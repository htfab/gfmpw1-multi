* NGSPICE file created from loopback9.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

.subckt loopback9 clk in[0] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17]
+ in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] out[0] out[10] out[11] out[1]
+ out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] rst_n vdd vss
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_172 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_15_139 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_11_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_120 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_31_215 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_16_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_13_109 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_16_Left_48 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA__12__A2 in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_79 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_23_173 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_14_259 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_19_Left_51 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_13_270 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_28_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_11_121 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_4_Left_36 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_31_216 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA__33__I clk vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_195 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_85 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_29_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_18_149 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_23_174 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_27_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_20_Left_52 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_10_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_24_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_30_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_12_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__24__A1 in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_119 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_7_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__15__A1 in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_16_97 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_1_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_175 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_131 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_239 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_70 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_29_ _09_ out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA__15__A2 rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_197 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_31_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_132 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_14_218 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_31_208 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_71 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_28_ in[14] in[15] out[7] _09_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor3_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_26_185 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_109 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_31_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_82 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_14_133 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_20_158 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_31_209 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_24_Left_56 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_72 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__27__A1 in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA__18__A1 in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
X_27_ in[14] out[7] out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_1
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_4_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_11_Left_43 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_26_186 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_3_83 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_134 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_20_159 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_30_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_26_ _08_ out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XTAP_TAPCELL_ROW_26_187 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_84 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_14_135 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_13_254 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_11_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_25_ in[12] in[13] out[5] _08_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor3_1
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_95 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_26_188 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_0_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_3_85 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_13_222 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_27_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_18_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_64 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_7_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_15_169 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_24_ in[12] out[5] out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_1
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_96 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_189 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_17_145 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_15_Left_47 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_16_253 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_22_170 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_11_118 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_13_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_18_Left_50 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_24_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_0_65 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_3_Left_35 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
X_23_ _07_ out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_4_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_6_97 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_25_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_146 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_22_171 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_119 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_203 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_0_66 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_20_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_22_ in[10] in[11] out[3] _07_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor3_1
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_29_199 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_6_98 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_3_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__11__A1 in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_17_147 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_299 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_8_104 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_204 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_67 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_21_ in[10] out[3] out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_1
XTAP_TAPCELL_ROW_6_99 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__11__A2 in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_25_181 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_17_148 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_16_267 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_8_105 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_205 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_68 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
X_20_ _06_ out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_7_Left_39 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_14_151 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_25_182 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_257 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_202 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_0_324 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_106 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_13_130 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_85 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_0_69 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_30_206 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_23_Left_55 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_20_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_11_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_183 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_31_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_16_214 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_107 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_10_Left_42 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_90 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_30_207 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_128 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_14_131 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_25_184 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_108 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_16_140 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_10_113 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_121 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_141 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_29_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_114 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_14_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_9_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_194 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_27_Left_59 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_3_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_25_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_142 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_0_328 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_22_167 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_14_Left_46 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_10_115 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_89 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_20_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_14_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_2_Left_34 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_28_195 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_16_143 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_218 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_22_168 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_7_100 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_31_Left_63 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_10_116 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_73 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_28_196 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_144 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_24_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_169 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_7_101 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_10_117 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_17_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_74 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_6_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_147 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_28_197 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_102 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_15_220 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_15_275 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_14_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_1_75 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_198 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_19_154 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_6_Left_38 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_7_103 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_13_127 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_9_Left_41 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_4_86 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_31_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_13_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_15_92 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_1_76 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_22_Left_54 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_19_155 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_180 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_13_128 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_87 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_31_70 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_9_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_31_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_156 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_267 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_13_129 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
X_19_ in[8] in[9] _05_ _06_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor3_1
XFILLER_0_26_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_4_88 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_6_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_190 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_19_157 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_21_163 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_18_ in[8] _05_ out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor2_1
XTAP_TAPCELL_ROW_4_89 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__31__A1 in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__22__A1 in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_5_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_10_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__13__A1 in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_27_191 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_26_Left_58 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_164 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_17_ _05_ out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_29_Left_61 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_13_Left_45 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__22__A2 in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__31__A2 in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__13__A2 in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_27_192 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_33_ clk out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_1_Left_33 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_21_165 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
X_16_ in[7] _03_ _04_ _05_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor3_1
XFILLER_0_31_324 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_30_Left_62 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_16_195 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_27_193 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_2_80 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_32_ _10_ out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_15_216 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_29_200 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_21_166 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_122 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_15_ in[0] rst_n _04_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor2_1
XFILLER_0_19_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_5_91 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__25__A1 in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__16__A1 in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_163 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_18_150 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_2_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_81 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_31_ in[16] in[17] out[9] _10_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor3_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_29_201 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_12_123 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_14_ _00_ _01_ _02_ _03_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor3_1
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_17_Left_49 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_5_92 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__25__A2 in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_88 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_18_151 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_176 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_30_ in[16] out[9] out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_202 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_5_Left_37 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_12_124 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_295 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_13_ in[1] in[2] _02_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_8_Left_40 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_5_93 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_16_143 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_113 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_18_152 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_24_177 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XPHY_EDGE_ROW_21_Left_53 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_125 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_263 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_28_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_12_ in[3] in[5] _01_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor2_1
XFILLER_0_29_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_25_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_31_328 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__28__A1 in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__19__A1 in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_5_94 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_5_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_27_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_153 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_24_178 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_110 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_126 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_11_ in[4] in[6] _00_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor2_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_31_210 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__28__A2 in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__19__A2 in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_16_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_123 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_16_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_13_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_137 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_2_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_179 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_9_111 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_160 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_31_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_211 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_36 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_21_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_138 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_1_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_9_112 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_15_136 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_222 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_20_161 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_28_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_25_Left_57 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_19_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_212 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_28_Left_60 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_12_Left_44 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_13_106 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_137 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_162 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_0_Left_32 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_31_213 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_13_129 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_93 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_77 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_138 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_14_235 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_31_214 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__21__A1 in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__30__A1 in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__12__A1 in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_78 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
.ends

