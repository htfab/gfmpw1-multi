magic
tech gf180mcuD
magscale 1 5
timestamp 1702357553
<< obsm1 >>
rect 672 1538 59304 58438
<< metal2 >>
rect 0 0 56 400
rect 26544 0 26600 400
rect 28560 0 28616 400
rect 28896 0 28952 400
rect 30576 0 30632 400
rect 30912 0 30968 400
rect 31920 0 31976 400
rect 32592 0 32648 400
rect 32928 0 32984 400
rect 33264 0 33320 400
rect 33600 0 33656 400
rect 33936 0 33992 400
rect 34272 0 34328 400
rect 34608 0 34664 400
rect 34944 0 35000 400
rect 37968 0 38024 400
rect 39984 0 40040 400
rect 40992 0 41048 400
<< obsm2 >>
rect 2238 430 59122 58427
rect 2238 400 26514 430
rect 26630 400 28530 430
rect 28646 400 28866 430
rect 28982 400 30546 430
rect 30662 400 30882 430
rect 30998 400 31890 430
rect 32006 400 32562 430
rect 32678 400 32898 430
rect 33014 400 33234 430
rect 33350 400 33570 430
rect 33686 400 33906 430
rect 34022 400 34242 430
rect 34358 400 34578 430
rect 34694 400 34914 430
rect 35030 400 37938 430
rect 38054 400 39954 430
rect 40070 400 40962 430
rect 41078 400 59122 430
<< metal3 >>
rect 59600 28896 60000 28952
rect 59600 28560 60000 28616
rect 59600 28224 60000 28280
rect 59600 27888 60000 27944
rect 59600 27552 60000 27608
rect 59600 27216 60000 27272
rect 59600 21840 60000 21896
rect 59600 20832 60000 20888
rect 59600 19152 60000 19208
rect 59600 18816 60000 18872
rect 59600 18480 60000 18536
rect 59600 18144 60000 18200
rect 59600 17808 60000 17864
rect 59600 17472 60000 17528
rect 59600 17136 60000 17192
<< obsm3 >>
rect 2233 28982 59600 58422
rect 2233 28866 59570 28982
rect 2233 28646 59600 28866
rect 2233 28530 59570 28646
rect 2233 28310 59600 28530
rect 2233 28194 59570 28310
rect 2233 27974 59600 28194
rect 2233 27858 59570 27974
rect 2233 27638 59600 27858
rect 2233 27522 59570 27638
rect 2233 27302 59600 27522
rect 2233 27186 59570 27302
rect 2233 21926 59600 27186
rect 2233 21810 59570 21926
rect 2233 20918 59600 21810
rect 2233 20802 59570 20918
rect 2233 19238 59600 20802
rect 2233 19122 59570 19238
rect 2233 18902 59600 19122
rect 2233 18786 59570 18902
rect 2233 18566 59600 18786
rect 2233 18450 59570 18566
rect 2233 18230 59600 18450
rect 2233 18114 59570 18230
rect 2233 17894 59600 18114
rect 2233 17778 59570 17894
rect 2233 17558 59600 17778
rect 2233 17442 59570 17558
rect 2233 17222 59600 17442
rect 2233 17106 59570 17222
rect 2233 1554 59600 17106
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
<< obsm4 >>
rect 17206 14177 17554 48767
rect 17774 14177 25234 48767
rect 25454 14177 32914 48767
rect 33134 14177 40594 48767
rect 40814 14177 41986 48767
<< labels >>
rlabel metal2 s 26544 0 26600 400 6 clk
port 1 nsew signal input
rlabel metal2 s 28896 0 28952 400 6 in[0]
port 2 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 in[10]
port 3 nsew signal input
rlabel metal2 s 34944 0 35000 400 6 in[11]
port 4 nsew signal input
rlabel metal2 s 40992 0 41048 400 6 in[12]
port 5 nsew signal input
rlabel metal3 s 59600 17136 60000 17192 6 in[13]
port 6 nsew signal input
rlabel metal2 s 39984 0 40040 400 6 in[14]
port 7 nsew signal input
rlabel metal3 s 59600 18816 60000 18872 6 in[15]
port 8 nsew signal input
rlabel metal3 s 59600 20832 60000 20888 6 in[16]
port 9 nsew signal input
rlabel metal3 s 59600 19152 60000 19208 6 in[17]
port 10 nsew signal input
rlabel metal3 s 59600 18480 60000 18536 6 in[18]
port 11 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 in[1]
port 12 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 in[2]
port 13 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 in[3]
port 14 nsew signal input
rlabel metal2 s 30912 0 30968 400 6 in[4]
port 15 nsew signal input
rlabel metal2 s 32592 0 32648 400 6 in[5]
port 16 nsew signal input
rlabel metal2 s 33936 0 33992 400 6 in[6]
port 17 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 in[7]
port 18 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 in[8]
port 19 nsew signal input
rlabel metal2 s 34608 0 34664 400 6 in[9]
port 20 nsew signal input
rlabel metal2 s 33600 0 33656 400 6 out[0]
port 21 nsew signal output
rlabel metal3 s 59600 28896 60000 28952 6 out[10]
port 22 nsew signal output
rlabel metal3 s 59600 28560 60000 28616 6 out[11]
port 23 nsew signal output
rlabel metal2 s 37968 0 38024 400 6 out[1]
port 24 nsew signal output
rlabel metal3 s 59600 21840 60000 21896 6 out[2]
port 25 nsew signal output
rlabel metal3 s 59600 17808 60000 17864 6 out[3]
port 26 nsew signal output
rlabel metal3 s 59600 17472 60000 17528 6 out[4]
port 27 nsew signal output
rlabel metal3 s 59600 18144 60000 18200 6 out[5]
port 28 nsew signal output
rlabel metal3 s 59600 27888 60000 27944 6 out[6]
port 29 nsew signal output
rlabel metal3 s 59600 28224 60000 28280 6 out[7]
port 30 nsew signal output
rlabel metal3 s 59600 27216 60000 27272 6 out[8]
port 31 nsew signal output
rlabel metal3 s 59600 27552 60000 27608 6 out[9]
port 32 nsew signal output
rlabel metal2 s 0 0 56 400 6 rst_n
port 33 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 35 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4221210
string GDS_FILE /home/htamas/test/caravel_user_project/openlane/unigate/runs/23_12_12_05_59/results/signoff/unigate.magic.gds
string GDS_START 403414
<< end >>

