magic
tech gf180mcuD
magscale 1 5
timestamp 1702354388
<< obsm1 >>
rect 672 1538 31304 30214
<< metal2 >>
rect 8064 31600 8120 32000
rect 13104 31600 13160 32000
rect 14784 31600 14840 32000
rect 19152 31600 19208 32000
rect 23856 31600 23912 32000
rect 24192 31600 24248 32000
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 3696 0 3752 400
rect 14784 0 14840 400
rect 15792 0 15848 400
rect 16128 0 16184 400
rect 16464 0 16520 400
rect 17136 0 17192 400
rect 19152 0 19208 400
<< obsm2 >>
rect 462 31570 8034 31600
rect 8150 31570 13074 31600
rect 13190 31570 14754 31600
rect 14870 31570 19122 31600
rect 19238 31570 23826 31600
rect 23942 31570 24162 31600
rect 24278 31570 31514 31600
rect 462 430 31514 31570
rect 462 350 642 430
rect 758 350 978 430
rect 1094 350 3666 430
rect 3782 350 14754 430
rect 14870 350 15762 430
rect 15878 350 16098 430
rect 16214 350 16434 430
rect 16550 350 17106 430
rect 17222 350 19122 430
rect 19238 350 31514 430
<< metal3 >>
rect 31600 29232 32000 29288
rect 0 27216 400 27272
rect 0 22176 400 22232
rect 31600 21504 32000 21560
rect 0 16800 400 16856
rect 31600 16464 32000 16520
rect 0 15456 400 15512
rect 31600 15456 32000 15512
rect 31600 15120 32000 15176
rect 31600 14784 32000 14840
rect 31600 14448 32000 14504
rect 31600 14112 32000 14168
rect 31600 13776 32000 13832
rect 0 12432 400 12488
rect 0 12096 400 12152
rect 0 5712 400 5768
<< obsm3 >>
rect 400 29318 31600 30282
rect 400 29202 31570 29318
rect 400 27302 31600 29202
rect 430 27186 31600 27302
rect 400 22262 31600 27186
rect 430 22146 31600 22262
rect 400 21590 31600 22146
rect 400 21474 31570 21590
rect 400 16886 31600 21474
rect 430 16770 31600 16886
rect 400 16550 31600 16770
rect 400 16434 31570 16550
rect 400 15542 31600 16434
rect 430 15426 31570 15542
rect 400 15206 31600 15426
rect 400 15090 31570 15206
rect 400 14870 31600 15090
rect 400 14754 31570 14870
rect 400 14534 31600 14754
rect 400 14418 31570 14534
rect 400 14198 31600 14418
rect 400 14082 31570 14198
rect 400 13862 31600 14082
rect 400 13746 31570 13862
rect 400 12518 31600 13746
rect 430 12402 31600 12518
rect 400 12182 31600 12402
rect 430 12066 31600 12182
rect 400 5798 31600 12066
rect 430 5682 31600 5798
rect 400 1470 31600 5682
<< metal4 >>
rect 2224 1538 2384 30214
rect 9904 1538 10064 30214
rect 17584 1538 17744 30214
rect 25264 1538 25424 30214
<< obsm4 >>
rect 854 1508 2194 29279
rect 2414 1508 9874 29279
rect 10094 1508 17554 29279
rect 17774 1508 25234 29279
rect 25454 1508 31122 29279
rect 854 1465 31122 1508
<< labels >>
rlabel metal2 s 0 0 56 400 6 clk
port 1 nsew signal input
rlabel metal3 s 0 27216 400 27272 6 in[0]
port 2 nsew signal input
rlabel metal3 s 31600 14784 32000 14840 6 in[10]
port 3 nsew signal input
rlabel metal3 s 31600 15120 32000 15176 6 in[11]
port 4 nsew signal input
rlabel metal2 s 16128 0 16184 400 6 in[12]
port 5 nsew signal input
rlabel metal2 s 16464 0 16520 400 6 in[13]
port 6 nsew signal input
rlabel metal3 s 31600 14448 32000 14504 6 in[14]
port 7 nsew signal input
rlabel metal3 s 31600 13776 32000 13832 6 in[15]
port 8 nsew signal input
rlabel metal3 s 31600 14112 32000 14168 6 in[16]
port 9 nsew signal input
rlabel metal2 s 336 0 392 400 6 in[17]
port 10 nsew signal input
rlabel metal2 s 672 0 728 400 6 in[18]
port 11 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 in[1]
port 12 nsew signal input
rlabel metal3 s 31600 16464 32000 16520 6 in[2]
port 13 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 in[3]
port 14 nsew signal input
rlabel metal2 s 14784 0 14840 400 6 in[4]
port 15 nsew signal input
rlabel metal3 s 0 5712 400 5768 6 in[5]
port 16 nsew signal input
rlabel metal3 s 0 12432 400 12488 6 in[6]
port 17 nsew signal input
rlabel metal3 s 0 15456 400 15512 6 in[7]
port 18 nsew signal input
rlabel metal3 s 0 22176 400 22232 6 in[8]
port 19 nsew signal input
rlabel metal2 s 14784 31600 14840 32000 6 in[9]
port 20 nsew signal input
rlabel metal3 s 31600 21504 32000 21560 6 out[0]
port 21 nsew signal output
rlabel metal3 s 31600 29232 32000 29288 6 out[10]
port 22 nsew signal output
rlabel metal2 s 19152 31600 19208 32000 6 out[11]
port 23 nsew signal output
rlabel metal3 s 31600 15456 32000 15512 6 out[1]
port 24 nsew signal output
rlabel metal2 s 19152 0 19208 400 6 out[2]
port 25 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 out[3]
port 26 nsew signal output
rlabel metal3 s 0 16800 400 16856 6 out[4]
port 27 nsew signal output
rlabel metal2 s 8064 31600 8120 32000 6 out[5]
port 28 nsew signal output
rlabel metal2 s 13104 31600 13160 32000 6 out[6]
port 29 nsew signal output
rlabel metal2 s 24192 31600 24248 32000 6 out[7]
port 30 nsew signal output
rlabel metal2 s 23856 31600 23912 32000 6 out[8]
port 31 nsew signal output
rlabel metal2 s 3696 0 3752 400 6 out[9]
port 32 nsew signal output
rlabel metal2 s 1008 0 1064 400 6 rst_n
port 33 nsew signal input
rlabel metal4 s 2224 1538 2384 30214 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 30214 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 30214 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 30214 6 vss
port 35 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32000 32000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3979300
string GDS_FILE /home/htamas/progs/gfmpw1-multi/openlane/rotfpga2a/runs/23_12_12_05_08/results/signoff/rotfpga2a.magic.gds
string GDS_START 228290
<< end >>

