module cells9 (clk,
    rst_n,
    vdd,
    vss,
    in,
    out);
 input clk;
 input rst_n;
 input vdd;
 input vss;
 input [17:0] in;
 output [11:0] out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire \cm_inst.cc_inst.in[0] ;
 wire \cm_inst.cc_inst.in[1] ;
 wire \cm_inst.cc_inst.in[2] ;
 wire \cm_inst.cc_inst.in[3] ;
 wire \cm_inst.cc_inst.in[4] ;
 wire \cm_inst.cc_inst.in[5] ;
 wire \cm_inst.cc_inst.out_notouch_[0] ;
 wire \cm_inst.cc_inst.out_notouch_[100] ;
 wire \cm_inst.cc_inst.out_notouch_[101] ;
 wire \cm_inst.cc_inst.out_notouch_[102] ;
 wire \cm_inst.cc_inst.out_notouch_[103] ;
 wire \cm_inst.cc_inst.out_notouch_[104] ;
 wire \cm_inst.cc_inst.out_notouch_[105] ;
 wire \cm_inst.cc_inst.out_notouch_[106] ;
 wire \cm_inst.cc_inst.out_notouch_[107] ;
 wire \cm_inst.cc_inst.out_notouch_[108] ;
 wire \cm_inst.cc_inst.out_notouch_[109] ;
 wire \cm_inst.cc_inst.out_notouch_[10] ;
 wire \cm_inst.cc_inst.out_notouch_[110] ;
 wire \cm_inst.cc_inst.out_notouch_[111] ;
 wire \cm_inst.cc_inst.out_notouch_[112] ;
 wire \cm_inst.cc_inst.out_notouch_[113] ;
 wire \cm_inst.cc_inst.out_notouch_[114] ;
 wire \cm_inst.cc_inst.out_notouch_[115] ;
 wire \cm_inst.cc_inst.out_notouch_[116] ;
 wire \cm_inst.cc_inst.out_notouch_[117] ;
 wire \cm_inst.cc_inst.out_notouch_[118] ;
 wire \cm_inst.cc_inst.out_notouch_[119] ;
 wire \cm_inst.cc_inst.out_notouch_[11] ;
 wire \cm_inst.cc_inst.out_notouch_[120] ;
 wire \cm_inst.cc_inst.out_notouch_[121] ;
 wire \cm_inst.cc_inst.out_notouch_[122] ;
 wire \cm_inst.cc_inst.out_notouch_[123] ;
 wire \cm_inst.cc_inst.out_notouch_[124] ;
 wire \cm_inst.cc_inst.out_notouch_[125] ;
 wire \cm_inst.cc_inst.out_notouch_[126] ;
 wire \cm_inst.cc_inst.out_notouch_[127] ;
 wire \cm_inst.cc_inst.out_notouch_[128] ;
 wire \cm_inst.cc_inst.out_notouch_[129] ;
 wire \cm_inst.cc_inst.out_notouch_[12] ;
 wire \cm_inst.cc_inst.out_notouch_[130] ;
 wire \cm_inst.cc_inst.out_notouch_[131] ;
 wire \cm_inst.cc_inst.out_notouch_[132] ;
 wire \cm_inst.cc_inst.out_notouch_[133] ;
 wire \cm_inst.cc_inst.out_notouch_[134] ;
 wire \cm_inst.cc_inst.out_notouch_[135] ;
 wire \cm_inst.cc_inst.out_notouch_[136] ;
 wire \cm_inst.cc_inst.out_notouch_[137] ;
 wire \cm_inst.cc_inst.out_notouch_[138] ;
 wire \cm_inst.cc_inst.out_notouch_[139] ;
 wire \cm_inst.cc_inst.out_notouch_[13] ;
 wire \cm_inst.cc_inst.out_notouch_[140] ;
 wire \cm_inst.cc_inst.out_notouch_[141] ;
 wire \cm_inst.cc_inst.out_notouch_[142] ;
 wire \cm_inst.cc_inst.out_notouch_[143] ;
 wire \cm_inst.cc_inst.out_notouch_[144] ;
 wire \cm_inst.cc_inst.out_notouch_[145] ;
 wire \cm_inst.cc_inst.out_notouch_[146] ;
 wire \cm_inst.cc_inst.out_notouch_[147] ;
 wire \cm_inst.cc_inst.out_notouch_[148] ;
 wire \cm_inst.cc_inst.out_notouch_[149] ;
 wire \cm_inst.cc_inst.out_notouch_[14] ;
 wire \cm_inst.cc_inst.out_notouch_[150] ;
 wire \cm_inst.cc_inst.out_notouch_[151] ;
 wire \cm_inst.cc_inst.out_notouch_[152] ;
 wire \cm_inst.cc_inst.out_notouch_[153] ;
 wire \cm_inst.cc_inst.out_notouch_[154] ;
 wire \cm_inst.cc_inst.out_notouch_[155] ;
 wire \cm_inst.cc_inst.out_notouch_[156] ;
 wire \cm_inst.cc_inst.out_notouch_[157] ;
 wire \cm_inst.cc_inst.out_notouch_[158] ;
 wire \cm_inst.cc_inst.out_notouch_[159] ;
 wire \cm_inst.cc_inst.out_notouch_[15] ;
 wire \cm_inst.cc_inst.out_notouch_[160] ;
 wire \cm_inst.cc_inst.out_notouch_[161] ;
 wire \cm_inst.cc_inst.out_notouch_[162] ;
 wire \cm_inst.cc_inst.out_notouch_[163] ;
 wire \cm_inst.cc_inst.out_notouch_[164] ;
 wire \cm_inst.cc_inst.out_notouch_[165] ;
 wire \cm_inst.cc_inst.out_notouch_[166] ;
 wire \cm_inst.cc_inst.out_notouch_[167] ;
 wire \cm_inst.cc_inst.out_notouch_[168] ;
 wire \cm_inst.cc_inst.out_notouch_[169] ;
 wire \cm_inst.cc_inst.out_notouch_[16] ;
 wire \cm_inst.cc_inst.out_notouch_[170] ;
 wire \cm_inst.cc_inst.out_notouch_[171] ;
 wire \cm_inst.cc_inst.out_notouch_[172] ;
 wire \cm_inst.cc_inst.out_notouch_[173] ;
 wire \cm_inst.cc_inst.out_notouch_[174] ;
 wire \cm_inst.cc_inst.out_notouch_[175] ;
 wire \cm_inst.cc_inst.out_notouch_[176] ;
 wire \cm_inst.cc_inst.out_notouch_[177] ;
 wire \cm_inst.cc_inst.out_notouch_[178] ;
 wire \cm_inst.cc_inst.out_notouch_[179] ;
 wire \cm_inst.cc_inst.out_notouch_[17] ;
 wire \cm_inst.cc_inst.out_notouch_[180] ;
 wire \cm_inst.cc_inst.out_notouch_[181] ;
 wire \cm_inst.cc_inst.out_notouch_[182] ;
 wire \cm_inst.cc_inst.out_notouch_[183] ;
 wire \cm_inst.cc_inst.out_notouch_[184] ;
 wire \cm_inst.cc_inst.out_notouch_[185] ;
 wire \cm_inst.cc_inst.out_notouch_[186] ;
 wire \cm_inst.cc_inst.out_notouch_[187] ;
 wire \cm_inst.cc_inst.out_notouch_[188] ;
 wire \cm_inst.cc_inst.out_notouch_[189] ;
 wire \cm_inst.cc_inst.out_notouch_[18] ;
 wire \cm_inst.cc_inst.out_notouch_[190] ;
 wire \cm_inst.cc_inst.out_notouch_[191] ;
 wire \cm_inst.cc_inst.out_notouch_[192] ;
 wire \cm_inst.cc_inst.out_notouch_[193] ;
 wire \cm_inst.cc_inst.out_notouch_[194] ;
 wire \cm_inst.cc_inst.out_notouch_[195] ;
 wire \cm_inst.cc_inst.out_notouch_[196] ;
 wire \cm_inst.cc_inst.out_notouch_[197] ;
 wire \cm_inst.cc_inst.out_notouch_[198] ;
 wire \cm_inst.cc_inst.out_notouch_[199] ;
 wire \cm_inst.cc_inst.out_notouch_[19] ;
 wire \cm_inst.cc_inst.out_notouch_[1] ;
 wire \cm_inst.cc_inst.out_notouch_[200] ;
 wire \cm_inst.cc_inst.out_notouch_[201] ;
 wire \cm_inst.cc_inst.out_notouch_[202] ;
 wire \cm_inst.cc_inst.out_notouch_[203] ;
 wire \cm_inst.cc_inst.out_notouch_[204] ;
 wire \cm_inst.cc_inst.out_notouch_[205] ;
 wire \cm_inst.cc_inst.out_notouch_[206] ;
 wire \cm_inst.cc_inst.out_notouch_[208] ;
 wire \cm_inst.cc_inst.out_notouch_[209] ;
 wire \cm_inst.cc_inst.out_notouch_[20] ;
 wire \cm_inst.cc_inst.out_notouch_[21] ;
 wire \cm_inst.cc_inst.out_notouch_[22] ;
 wire \cm_inst.cc_inst.out_notouch_[23] ;
 wire \cm_inst.cc_inst.out_notouch_[24] ;
 wire \cm_inst.cc_inst.out_notouch_[25] ;
 wire \cm_inst.cc_inst.out_notouch_[26] ;
 wire \cm_inst.cc_inst.out_notouch_[27] ;
 wire \cm_inst.cc_inst.out_notouch_[28] ;
 wire \cm_inst.cc_inst.out_notouch_[29] ;
 wire \cm_inst.cc_inst.out_notouch_[2] ;
 wire \cm_inst.cc_inst.out_notouch_[30] ;
 wire \cm_inst.cc_inst.out_notouch_[31] ;
 wire \cm_inst.cc_inst.out_notouch_[32] ;
 wire \cm_inst.cc_inst.out_notouch_[33] ;
 wire \cm_inst.cc_inst.out_notouch_[34] ;
 wire \cm_inst.cc_inst.out_notouch_[35] ;
 wire \cm_inst.cc_inst.out_notouch_[36] ;
 wire \cm_inst.cc_inst.out_notouch_[37] ;
 wire \cm_inst.cc_inst.out_notouch_[38] ;
 wire \cm_inst.cc_inst.out_notouch_[39] ;
 wire \cm_inst.cc_inst.out_notouch_[3] ;
 wire \cm_inst.cc_inst.out_notouch_[40] ;
 wire \cm_inst.cc_inst.out_notouch_[41] ;
 wire \cm_inst.cc_inst.out_notouch_[42] ;
 wire \cm_inst.cc_inst.out_notouch_[43] ;
 wire \cm_inst.cc_inst.out_notouch_[44] ;
 wire \cm_inst.cc_inst.out_notouch_[45] ;
 wire \cm_inst.cc_inst.out_notouch_[46] ;
 wire \cm_inst.cc_inst.out_notouch_[47] ;
 wire \cm_inst.cc_inst.out_notouch_[48] ;
 wire \cm_inst.cc_inst.out_notouch_[49] ;
 wire \cm_inst.cc_inst.out_notouch_[4] ;
 wire \cm_inst.cc_inst.out_notouch_[50] ;
 wire \cm_inst.cc_inst.out_notouch_[51] ;
 wire \cm_inst.cc_inst.out_notouch_[52] ;
 wire \cm_inst.cc_inst.out_notouch_[53] ;
 wire \cm_inst.cc_inst.out_notouch_[54] ;
 wire \cm_inst.cc_inst.out_notouch_[55] ;
 wire \cm_inst.cc_inst.out_notouch_[56] ;
 wire \cm_inst.cc_inst.out_notouch_[57] ;
 wire \cm_inst.cc_inst.out_notouch_[58] ;
 wire \cm_inst.cc_inst.out_notouch_[59] ;
 wire \cm_inst.cc_inst.out_notouch_[5] ;
 wire \cm_inst.cc_inst.out_notouch_[60] ;
 wire \cm_inst.cc_inst.out_notouch_[61] ;
 wire \cm_inst.cc_inst.out_notouch_[62] ;
 wire \cm_inst.cc_inst.out_notouch_[63] ;
 wire \cm_inst.cc_inst.out_notouch_[64] ;
 wire \cm_inst.cc_inst.out_notouch_[65] ;
 wire \cm_inst.cc_inst.out_notouch_[66] ;
 wire \cm_inst.cc_inst.out_notouch_[67] ;
 wire \cm_inst.cc_inst.out_notouch_[68] ;
 wire \cm_inst.cc_inst.out_notouch_[69] ;
 wire \cm_inst.cc_inst.out_notouch_[6] ;
 wire \cm_inst.cc_inst.out_notouch_[70] ;
 wire \cm_inst.cc_inst.out_notouch_[71] ;
 wire \cm_inst.cc_inst.out_notouch_[72] ;
 wire \cm_inst.cc_inst.out_notouch_[73] ;
 wire \cm_inst.cc_inst.out_notouch_[74] ;
 wire \cm_inst.cc_inst.out_notouch_[75] ;
 wire \cm_inst.cc_inst.out_notouch_[76] ;
 wire \cm_inst.cc_inst.out_notouch_[77] ;
 wire \cm_inst.cc_inst.out_notouch_[78] ;
 wire \cm_inst.cc_inst.out_notouch_[79] ;
 wire \cm_inst.cc_inst.out_notouch_[7] ;
 wire \cm_inst.cc_inst.out_notouch_[80] ;
 wire \cm_inst.cc_inst.out_notouch_[81] ;
 wire \cm_inst.cc_inst.out_notouch_[82] ;
 wire \cm_inst.cc_inst.out_notouch_[83] ;
 wire \cm_inst.cc_inst.out_notouch_[84] ;
 wire \cm_inst.cc_inst.out_notouch_[85] ;
 wire \cm_inst.cc_inst.out_notouch_[86] ;
 wire \cm_inst.cc_inst.out_notouch_[87] ;
 wire \cm_inst.cc_inst.out_notouch_[88] ;
 wire \cm_inst.cc_inst.out_notouch_[89] ;
 wire \cm_inst.cc_inst.out_notouch_[8] ;
 wire \cm_inst.cc_inst.out_notouch_[90] ;
 wire \cm_inst.cc_inst.out_notouch_[91] ;
 wire \cm_inst.cc_inst.out_notouch_[92] ;
 wire \cm_inst.cc_inst.out_notouch_[93] ;
 wire \cm_inst.cc_inst.out_notouch_[94] ;
 wire \cm_inst.cc_inst.out_notouch_[95] ;
 wire \cm_inst.cc_inst.out_notouch_[96] ;
 wire \cm_inst.cc_inst.out_notouch_[97] ;
 wire \cm_inst.cc_inst.out_notouch_[98] ;
 wire \cm_inst.cc_inst.out_notouch_[99] ;
 wire \cm_inst.cc_inst.out_notouch_[9] ;
 wire \cm_inst.page[0] ;
 wire \cm_inst.page[1] ;
 wire \cm_inst.page[2] ;
 wire \cm_inst.page[3] ;
 wire \cm_inst.page[4] ;
 wire \cm_inst.page[5] ;
 wire \ro_inst.counter[0] ;
 wire \ro_inst.counter[10] ;
 wire \ro_inst.counter[11] ;
 wire \ro_inst.counter[12] ;
 wire \ro_inst.counter[13] ;
 wire \ro_inst.counter[14] ;
 wire \ro_inst.counter[15] ;
 wire \ro_inst.counter[16] ;
 wire \ro_inst.counter[17] ;
 wire \ro_inst.counter[18] ;
 wire \ro_inst.counter[19] ;
 wire \ro_inst.counter[1] ;
 wire \ro_inst.counter[20] ;
 wire \ro_inst.counter[21] ;
 wire \ro_inst.counter[22] ;
 wire \ro_inst.counter[23] ;
 wire \ro_inst.counter[24] ;
 wire \ro_inst.counter[25] ;
 wire \ro_inst.counter[26] ;
 wire \ro_inst.counter[27] ;
 wire \ro_inst.counter[28] ;
 wire \ro_inst.counter[29] ;
 wire \ro_inst.counter[2] ;
 wire \ro_inst.counter[30] ;
 wire \ro_inst.counter[31] ;
 wire \ro_inst.counter[32] ;
 wire \ro_inst.counter[33] ;
 wire \ro_inst.counter[34] ;
 wire \ro_inst.counter[3] ;
 wire \ro_inst.counter[4] ;
 wire \ro_inst.counter[5] ;
 wire \ro_inst.counter[6] ;
 wire \ro_inst.counter[7] ;
 wire \ro_inst.counter[8] ;
 wire \ro_inst.counter[9] ;
 wire \ro_inst.counter_n[0] ;
 wire \ro_inst.counter_n[10] ;
 wire \ro_inst.counter_n[11] ;
 wire \ro_inst.counter_n[12] ;
 wire \ro_inst.counter_n[13] ;
 wire \ro_inst.counter_n[14] ;
 wire \ro_inst.counter_n[15] ;
 wire \ro_inst.counter_n[16] ;
 wire \ro_inst.counter_n[17] ;
 wire \ro_inst.counter_n[18] ;
 wire \ro_inst.counter_n[19] ;
 wire \ro_inst.counter_n[1] ;
 wire \ro_inst.counter_n[20] ;
 wire \ro_inst.counter_n[21] ;
 wire \ro_inst.counter_n[22] ;
 wire \ro_inst.counter_n[23] ;
 wire \ro_inst.counter_n[24] ;
 wire \ro_inst.counter_n[25] ;
 wire \ro_inst.counter_n[26] ;
 wire \ro_inst.counter_n[27] ;
 wire \ro_inst.counter_n[28] ;
 wire \ro_inst.counter_n[29] ;
 wire \ro_inst.counter_n[2] ;
 wire \ro_inst.counter_n[30] ;
 wire \ro_inst.counter_n[31] ;
 wire \ro_inst.counter_n[32] ;
 wire \ro_inst.counter_n[33] ;
 wire \ro_inst.counter_n[34] ;
 wire \ro_inst.counter_n[3] ;
 wire \ro_inst.counter_n[4] ;
 wire \ro_inst.counter_n[5] ;
 wire \ro_inst.counter_n[6] ;
 wire \ro_inst.counter_n[7] ;
 wire \ro_inst.counter_n[8] ;
 wire \ro_inst.counter_n[9] ;
 wire \ro_inst.enable ;
 wire \ro_inst.ring[0] ;
 wire \ro_inst.ring[1] ;
 wire \ro_inst.ring[2] ;
 wire \ro_inst.running ;
 wire \ro_inst.saved_signal ;
 wire \ro_inst.signal ;
 wire \ro_inst.slow_clk_n ;
 wire \ro_sel[0] ;
 wire \ro_sel[1] ;
 wire \ro_sel[2] ;

 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__249__I (.I(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__250__I (.I(\cm_inst.page[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__262__I (.I(_033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__263__S0 (.I(_031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__263__S1 (.I(_034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__264__I (.I(\cm_inst.page[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__269__I (.I(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__270__S (.I(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__280__S (.I(_051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__281__A1 (.I(_034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__284__A2 (.I(_035_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__290__I (.I(\cm_inst.page[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__291__S0 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__291__S1 (.I(_061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__292__I (.I(\cm_inst.page[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__294__S0 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__294__S1 (.I(_064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__297__S0 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__297__S1 (.I(_061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__300__S1 (.I(_064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__302__S (.I(_033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__303__A2 (.I(_073_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__305__I (.I(_075_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__308__S0 (.I(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__309__S (.I(_051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__319__A2 (.I(_080_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__322__S0 (.I(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__324__I (.I(_093_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__326__S1 (.I(_095_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__327__S (.I(_051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__328__I (.I(_061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__330__S (.I(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__333__I (.I(_093_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__338__I (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__339__S (.I(_108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__340__B (.I(_031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__349__I (.I(_093_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__357__B (.I(_075_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__363__S1 (.I(_095_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__365__S (.I(_133_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__366__S (.I(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__368__S1 (.I(_064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__372__S1 (.I(_064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__376__S (.I(_033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__377__A2 (.I(_145_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__381__S1 (.I(_095_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__382__I (.I(_093_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__383__I (.I(_061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__385__I1 (.I(_152_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__385__S (.I(_133_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__386__S (.I(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__391__S (.I(_108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__392__B (.I(_031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__402__B (.I(_034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__406__I (.I(_075_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__409__S (.I(_133_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__420__S (.I(_033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__421__A2 (.I(_187_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__424__S1 (.I(_095_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__426__S (.I(_133_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__432__B (.I(_031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__442__B (.I(_034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__451__S (.I(_051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__452__S (.I(_075_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__454__S0 (.I(_108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__455__S0 (.I(_108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__470__I (.I(in[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__471__I (.I(in[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__472__I (.I(in[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__473__B (.I(in[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__475__I0 (.I(in[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__476__I0 (.I(in[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__477__I0 (.I(in[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__478__I (.I(in[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__483__I0 (.I(in[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__483__I1 (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__485__I0 (.I(in[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__485__I1 (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__486__I0 (.I(in[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__486__I1 (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__487__I0 (.I(in[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__487__I1 (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__488__I0 (.I(in[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__488__I1 (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__489__I0 (.I(in[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__489__I1 (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__492__A1 (.I(in[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__492__A2 (.I(in[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__492__A3 (.I(in[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__492__A4 (.I(in[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__493__I0 (.I(in[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__494__I0 (.I(in[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__495__I0 (.I(in[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__496__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__497__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__498__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__499__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__500__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__501__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__502__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__503__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__504__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__505__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__506__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__507__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__508__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__509__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__510__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA__511__CLK (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addf_1_inst_A  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addf_1_inst_B  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addf_1_inst_CI  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addf_2_inst_A  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addf_2_inst_B  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addf_2_inst_CI  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addf_4_inst_A  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addf_4_inst_B  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addf_4_inst_CI  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addh_1_inst_A  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addh_1_inst_B  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addh_2_inst_A  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addh_2_inst_B  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addh_4_inst_A  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.addh_4_inst_B  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and2_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and2_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and2_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and2_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and2_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and2_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and3_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and3_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and3_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and3_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and3_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and3_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and3_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and3_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and3_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_1_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_2_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.and4_4_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_1_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_1_inst_C  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_2_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_2_inst_C  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_4_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi211_4_inst_C  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi21_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi21_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi21_1_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi21_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi21_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi21_2_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi21_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi21_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi21_4_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_1_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_1_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_1_inst_C  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_2_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_2_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_2_inst_C  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_4_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_4_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi221_4_inst_C  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_1_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_1_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_1_inst_C1  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_1_inst_C2  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_2_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_2_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_2_inst_C1  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_2_inst_C2  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_4_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_4_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_4_inst_C1  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi222_4_inst_C2  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_1_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_1_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_2_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_2_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_4_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.aoi22_4_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.buf_12_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.buf_16_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.buf_1_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.buf_20_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.buf_2_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.buf_3_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.buf_4_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.buf_8_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_12_inst_EN  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_12_inst_I  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_16_inst_EN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_16_inst_I  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_1_inst_EN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_1_inst_I  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_2_inst_EN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_2_inst_I  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_3_inst_EN  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_3_inst_I  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_4_inst_EN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_4_inst_I  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_8_inst_EN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.bufz_8_inst_I  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkbuf_12_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkbuf_16_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkbuf_1_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkbuf_20_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkbuf_2_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkbuf_3_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkbuf_4_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkbuf_8_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkinv_12_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkinv_16_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkinv_1_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkinv_20_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkinv_2_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkinv_3_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkinv_4_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.clkinv_8_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnq_1_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnq_2_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnq_4_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_SETN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_SETN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_SETN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffq_1_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffq_2_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffq_4_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrnq_1_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrnq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrnq_1_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrnq_2_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrnq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrnq_2_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrnq_4_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrnq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrnq_4_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffsnq_1_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffsnq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffsnq_1_inst_SETN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffsnq_2_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffsnq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffsnq_2_inst_SETN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffsnq_4_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffsnq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dffsnq_4_inst_SETN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlya_1_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlya_2_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlya_4_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlyb_1_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlyb_2_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlyb_4_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlyc_1_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlyc_2_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlyc_4_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlyd_1_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlyd_2_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.dlyd_4_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtn_1_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtn_1_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtn_1_inst_TE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtn_2_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtn_2_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtn_2_inst_TE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtn_4_inst_CLKN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtn_4_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtn_4_inst_TE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtp_2_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtp_2_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtp_2_inst_TE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtp_4_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtp_4_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.icgtp_4_inst_TE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.inv_12_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.inv_16_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.inv_1_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.inv_20_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.inv_2_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.inv_3_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.inv_4_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.inv_8_inst_I  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_12_inst_EN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_12_inst_I  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_1_inst_EN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_1_inst_I  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_2_inst_EN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_2_inst_I  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_3_inst_EN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_3_inst_I  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_4_inst_EN  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_4_inst_I  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_8_inst_EN  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.invz_8_inst_I  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latq_1_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latq_1_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latq_2_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latq_2_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latq_4_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latq_4_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrnq_1_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrnq_1_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrnq_1_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrnq_2_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrnq_2_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrnq_2_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrnq_4_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrnq_4_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrnq_4_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latsnq_1_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latsnq_1_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latsnq_1_inst_SETN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latsnq_2_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latsnq_2_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latsnq_2_inst_SETN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latsnq_4_inst_D  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latsnq_4_inst_E  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.latsnq_4_inst_SETN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux2_1_inst_I0  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux2_1_inst_I1  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux2_1_inst_S  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux2_2_inst_I0  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux2_2_inst_I1  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux2_2_inst_S  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux2_4_inst_I0  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux2_4_inst_I1  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux2_4_inst_S  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_1_inst_I0  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_1_inst_I1  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_1_inst_I2  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_1_inst_I3  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_1_inst_S0  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_1_inst_S1  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_2_inst_I0  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_2_inst_I1  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_2_inst_I2  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_2_inst_I3  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_2_inst_S0  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_2_inst_S1  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_4_inst_I0  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_4_inst_I1  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_4_inst_I2  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_4_inst_I3  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_4_inst_S0  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.mux4_4_inst_S1  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand2_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand2_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand2_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand2_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand2_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand2_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand3_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand3_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand3_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand3_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand3_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand3_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand3_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand3_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand3_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_1_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_2_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nand4_4_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor2_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor2_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor2_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor2_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor2_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor2_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor3_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor3_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor3_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor3_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor3_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor3_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor3_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor3_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor3_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_1_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_2_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.nor4_4_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_1_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_1_inst_C  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_2_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_2_inst_C  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_4_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai211_4_inst_C  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai21_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai21_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai21_1_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai21_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai21_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai21_2_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai21_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai21_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai21_4_inst_B  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_1_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_1_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_1_inst_C  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_2_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_2_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_2_inst_C  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_4_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_4_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai221_4_inst_C  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_1_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_1_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_1_inst_C1  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_1_inst_C2  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_2_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_2_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_2_inst_C1  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_2_inst_C2  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_4_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_4_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_4_inst_C1  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai222_4_inst_C2  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_1_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_1_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_2_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_2_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_4_inst_B1  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai22_4_inst_B2  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_1_inst_B  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_2_inst_B  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai31_4_inst_B  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_1_inst_B1  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_1_inst_B2  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_2_inst_B1  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_2_inst_B2  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_4_inst_B1  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai32_4_inst_B2  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_1_inst_B1  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_1_inst_B2  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_1_inst_B3  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_2_inst_B1  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_2_inst_B2  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_2_inst_B3  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_4_inst_B1  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_4_inst_B2  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.oai33_4_inst_B3  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or2_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or2_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or2_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or2_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or2_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or2_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or3_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or3_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or3_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or3_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or3_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or3_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or3_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or3_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or3_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_1_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_2_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.or4_4_inst_A4  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_1_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_1_inst_SE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_1_inst_SI  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_2_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_2_inst_SE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_2_inst_SI  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_4_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_4_inst_SE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffq_4_inst_SI  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_SE  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_SI  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SE  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SI  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_SE  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_SI  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SE  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SETN  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SI  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SE  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SETN  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SI  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_RN  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SE  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SETN  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SI  (.I(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SI  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SI  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_CLK  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_D  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SE  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SETN  (.I(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SI  (.I(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor2_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor2_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor2_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor2_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor2_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor2_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor3_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor3_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor3_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor3_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor3_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor3_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor3_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor3_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xnor3_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor2_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor2_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor2_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor2_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor2_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor2_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor3_1_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor3_1_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor3_1_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor3_2_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor3_2_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor3_2_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor3_4_inst_A1  (.I(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor3_4_inst_A2  (.I(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_cm_inst.cc_inst.xor3_4_inst_A3  (.I(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[10].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[11].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[12].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[13].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[14].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[15].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[16].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[17].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[18].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[19].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[1].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[20].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[21].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[22].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[23].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[24].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[25].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[26].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[27].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[28].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[29].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[2].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[30].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[31].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[32].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[33].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[34].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[3].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[4].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[5].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[6].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[7].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[8].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.gcount[9].div_flop_RN  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__antenna \ANTENNA_ro_inst.slow_clock_inv_I  (.I(in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_0_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_0_494 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_0_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_0_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_0_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_0_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_10_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_10_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_10_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_10_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_10_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_10_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_10_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_10_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_10_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_10_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_10_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_10_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_10_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_10_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_10_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_10_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_10_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_11_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_11_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_11_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_11_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_11_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_11_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_11_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_11_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_11_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_11_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_11_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_11_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_11_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_433 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_449 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_11_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_11_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_11_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_11_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_11_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_12_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_12_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_12_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_12_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_12_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_12_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_12_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_12_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_12_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_12_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_12_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_12_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_12_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_12_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_12_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_12_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_12_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_12_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_12_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_12_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_12_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_433 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_12_449 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_491 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_495 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_499 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_12_503 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_12_507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_13_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_13_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_13_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_13_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_13_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_13_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_13_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_13_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_13_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_13_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_13_436 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_13_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_13_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_13_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_13_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_13_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_13_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_13_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_14_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_14_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_14_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_14_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_14_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_14_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_14_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_14_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_14_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_14_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_14_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_14_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_14_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_14_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_14_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_14_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_14_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_14_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_449 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_14_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_14_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_15_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_15_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_15_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_15_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_15_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_15_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_15_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_15_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_15_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_15_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_15_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_15_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_15_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_16_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_16_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_16_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_16_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_16_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_16_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_16_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_16_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_16_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_16_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_16_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_16_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_16_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_449 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_493 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_16_497 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_16_501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_17_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_17_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_17_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_17_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_17_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_17_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_17_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_17_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_17_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_17_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_17_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_17_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_17_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_17_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_17_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_17_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_17_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_17_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_17_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_17_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_17_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_17_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_18_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_18_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_18_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_18_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_18_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_18_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_18_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_18_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_18_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_18_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_18_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_18_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_18_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_18_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_18_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_18_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_18_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_18_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_18_423 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_18_429 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_436 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_18_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_18_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_18_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_18_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_18_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_18_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_18_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_19_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_19_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_19_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_19_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_19_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_19_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_19_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_19_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_19_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_19_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_19_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_19_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_19_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_19_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_19_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_19_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_1_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_1_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_1_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_1_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_1_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_1_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_1_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_1_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_1_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_1_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_1_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_1_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_1_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_20_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_20_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_20_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_20_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_20_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_20_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_20_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_20_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_20_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_436 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_20_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_20_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_21_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_21_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_21_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_21_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_21_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_21_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_21_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_21_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_21_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_21_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_476 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_480 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_21_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_21_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_21_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_21_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_21_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_21_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_22_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_22_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_22_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_22_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_22_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_22_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_22_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_22_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_22_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_22_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_22_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_22_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_22_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_22_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_22_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_22_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_23_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_23_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_23_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_23_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_23_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_23_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_23_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_23_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_23_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_23_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_23_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_23_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_446 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_23_458 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_23_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_23_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_23_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_23_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_23_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_23_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_23_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_23_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_24_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_24_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_423 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_24_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_24_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_24_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_24_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_24_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_24_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_24_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_24_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_25_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_25_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_25_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_439 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_25_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_25_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_25_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_25_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_25_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_26_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_26_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_26_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_26_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_26_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_26_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_26_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_26_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_26_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_26_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_26_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_26_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_26_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_26_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_26_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_26_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_26_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_26_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_26_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_26_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_26_463 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_26_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_26_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_26_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_26_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_26_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_27_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_27_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_27_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_27_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_27_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_27_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_27_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_27_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_27_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_27_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_27_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_27_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_27_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_27_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_27_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_27_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_27_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_27_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_28_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_28_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_28_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_28_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_28_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_28_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_28_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_28_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_28_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_28_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_28_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_28_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_28_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_495 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_28_499 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_28_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_28_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_28_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_29_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_29_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_29_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_29_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_29_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_29_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_29_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_29_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_29_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_29_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_29_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_446 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_450 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_467 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_471 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_29_475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_29_481 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_485 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_29_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_29_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_29_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_29_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_29_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_29_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_29_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_2_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_2_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_2_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_2_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_2_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_2_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_2_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_2_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_2_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_2_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_2_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_2_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_2_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_2_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_2_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_30_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_30_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_30_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_30_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_30_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_30_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_30_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_30_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_30_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_30_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_30_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_30_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_30_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_30_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_30_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_30_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_30_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_30_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_30_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_30_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_439 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_30_474 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_483 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_491 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_30_495 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_30_503 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_30_507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_31_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_31_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_31_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_31_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_31_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_31_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_31_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_31_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_31_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_31_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_31_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_31_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_31_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_31_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_31_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_31_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_31_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_31_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_31_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_31_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_31_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_31_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_31_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_32_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_32_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_32_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_32_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_32_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_32_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_32_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_32_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_32_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_32_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_32_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_32_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_32_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_464 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_32_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_32_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_33_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_33_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_180 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_33_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_33_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_33_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_33_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_33_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_33_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_33_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_33_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_33_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_33_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_33_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_33_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_33_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_33_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_33_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_33_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_33_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_33_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_33_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_33_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_34_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_34_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_34_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_34_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_34_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_34_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_34_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_34_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_34_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_34_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_34_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_34_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_34_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_34_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_470 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_474 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_34_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_490 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_494 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_34_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_34_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_34_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_35_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_35_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_35_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_35_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_35_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_35_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_35_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_35_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_35_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_35_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_35_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_35_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_35_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_35_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_35_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_35_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_35_449 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_35_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_35_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_35_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_36_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_36_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_36_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_36_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_36_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_36_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_423 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_429 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_36_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_36_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_36_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_36_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_36_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_37_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_37_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_37_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_37_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_37_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_37_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_37_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_37_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_37_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_37_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_474 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_476 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_37_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_37_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_37_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_37_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_37_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_37_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_37_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_37_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_38_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_38_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_38_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_38_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_38_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_38_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_38_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_38_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_38_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_38_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_38_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_38_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_38_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_38_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_38_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_38_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_420 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_38_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_446 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_38_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_450 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_38_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_490 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_494 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_38_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_38_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_38_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_38_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_39_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_39_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_39_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_39_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_39_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_39_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_39_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_39_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_39_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_39_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_39_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_39_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_39_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_39_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_39_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_39_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_39_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_39_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_39_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_39_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_456 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_39_458 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_39_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_39_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_39_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_39_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_39_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_3_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_3_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_3_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_3_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_3_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_3_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_3_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_3_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_3_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_3_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_3_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_3_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_3_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_3_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_3_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_3_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_3_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_3_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_3_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_3_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_3_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_3_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_3_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_3_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_3_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_3_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_3_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_3_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_40_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_40_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_40_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_40_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_40_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_40_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_40_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_40_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_40_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_40_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_40_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_40_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_40_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_40_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_40_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_40_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_40_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_40_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_40_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_40_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_41_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_41_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_41_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_41_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_41_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_41_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_41_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_41_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_476 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_480 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_41_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_41_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_41_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_41_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_41_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_41_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_42_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_42_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_42_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_42_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_42_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_42_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_42_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_42_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_42_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_42_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_42_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_42_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_42_473 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_42_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_43_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_43_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_43_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_43_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_43_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_43_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_43_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_43_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_43_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_43_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_43_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_43_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_43_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_43_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_43_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_43_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_43_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_450 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_43_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_455 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_459 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_463 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_43_467 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_43_483 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_43_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_43_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_43_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_43_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_43_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_43_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_44_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_44_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_44_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_44_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_44_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_44_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_44_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_44_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_44_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_44_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_44_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_44_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_44_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_44_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_44_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_44_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_44_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_44_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_44_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_44_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_44_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_44_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_44_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_44_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_44_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_44_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_44_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_45_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_45_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_45_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_45_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_45_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_45_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_45_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_45_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_45_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_45_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_45_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_45_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_45_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_45_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_45_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_45_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_46_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_46_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_46_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_46_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_46_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_46_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_46_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_46_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_46_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_46_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_46_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_46_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_46_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_46_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_46_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_46_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_46_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_47_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_47_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_47_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_47_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_47_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_47_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_47_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_47_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_47_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_47_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_47_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_47_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_47_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_47_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_47_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_47_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_48_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_48_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_48_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_48_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_48_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_48_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_48_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_48_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_48_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_48_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_48_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_48_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_48_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_48_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_48_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_48_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_48_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_49_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_49_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_49_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_49_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_49_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_49_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_49_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_49_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_49_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_49_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_49_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_49_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_49_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_49_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_49_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_49_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_49_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_49_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_49_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_49_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_4_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_4_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_4_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_4_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_4_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_4_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_4_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_4_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_4_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_4_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_4_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_4_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_4_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_4_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_4_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_4_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_4_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_4_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_4_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_4_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_4_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_50_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_50_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_50_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_50_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_50_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_50_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_50_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_50_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_50_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_50_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_50_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_50_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_50_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_50_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_50_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_50_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_50_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_51_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_51_494 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_51_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_51_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_51_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_51_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_5_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_5_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_5_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_5_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_5_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_5_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_5_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_5_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_5_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_5_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_5_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_5_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_5_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_5_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_5_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_5_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_5_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_5_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_5_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_5_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_5_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_5_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_5_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_5_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_5_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_5_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_6_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_6_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_6_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_6_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_6_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_6_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_6_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_6_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_6_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_6_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_6_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_6_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_6_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_6_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_6_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_6_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_6_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_6_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_6_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_6_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_6_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_6_464 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_6_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_6_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_6_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_7_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_7_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_7_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_7_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_7_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_7_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_7_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_7_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_7_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_7_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_7_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_7_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_7_450 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_7_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_7_463 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_7_466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_7_470 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_7_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_7_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_7_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_7_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_7_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_8_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_8_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_8_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_8_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_8_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_8_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_8_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_8_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_8_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_8_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_8_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_8_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_8_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_8_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_8_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_8_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_8_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_8_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_8_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_8_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_449 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_8_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_8_463 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_8_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_8_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_9_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_9_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_9_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_9_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_9_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_9_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_9_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_9_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_9_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_9_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_9_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_9_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_9_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_9_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_9_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_9_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_0_9_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _244_ (.I(\ro_inst.enable ),
    .Z(_016_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _245_ (.I(\cm_inst.page[4] ),
    .Z(_017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _246_ (.I(_017_),
    .Z(_018_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _247_ (.I(\cm_inst.page[0] ),
    .Z(_019_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _248_ (.I(_019_),
    .Z(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _249_ (.I(_020_),
    .Z(_021_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _250_ (.I(\cm_inst.page[1] ),
    .Z(_022_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _251_ (.I(_022_),
    .Z(_023_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _252_ (.I(_023_),
    .Z(_024_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _253_ (.I0(\cm_inst.cc_inst.out_notouch_[96] ),
    .I1(\cm_inst.cc_inst.out_notouch_[104] ),
    .I2(\cm_inst.cc_inst.out_notouch_[112] ),
    .I3(\cm_inst.cc_inst.out_notouch_[120] ),
    .S0(_021_),
    .S1(_024_),
    .Z(_025_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _254_ (.I0(\cm_inst.cc_inst.out_notouch_[64] ),
    .I1(\cm_inst.cc_inst.out_notouch_[72] ),
    .I2(\cm_inst.cc_inst.out_notouch_[80] ),
    .I3(\cm_inst.cc_inst.out_notouch_[88] ),
    .S0(_021_),
    .S1(_024_),
    .Z(_026_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _255_ (.I0(\cm_inst.cc_inst.out_notouch_[32] ),
    .I1(\cm_inst.cc_inst.out_notouch_[40] ),
    .I2(\cm_inst.cc_inst.out_notouch_[48] ),
    .I3(\cm_inst.cc_inst.out_notouch_[56] ),
    .S0(_021_),
    .S1(_024_),
    .Z(_027_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _256_ (.I0(\cm_inst.cc_inst.out_notouch_[0] ),
    .I1(\cm_inst.cc_inst.out_notouch_[8] ),
    .I2(\cm_inst.cc_inst.out_notouch_[16] ),
    .I3(\cm_inst.cc_inst.out_notouch_[24] ),
    .S0(_021_),
    .S1(_024_),
    .Z(_028_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _257_ (.I(\cm_inst.page[2] ),
    .ZN(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _258_ (.I(_029_),
    .Z(_030_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _259_ (.I(_030_),
    .Z(_031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _260_ (.I(\cm_inst.page[3] ),
    .ZN(_032_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _261_ (.I(_032_),
    .Z(_033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _262_ (.I(_033_),
    .Z(_034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _263_ (.I0(_025_),
    .I1(_026_),
    .I2(_027_),
    .I3(_028_),
    .S0(_031_),
    .S1(_034_),
    .Z(_035_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _264_ (.I(\cm_inst.page[1] ),
    .ZN(_036_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _265_ (.I(_036_),
    .Z(_037_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _266_ (.I(_019_),
    .Z(_038_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _267_ (.I(_038_),
    .Z(_039_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _268_ (.A1(_037_),
    .A2(_039_),
    .ZN(_040_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _269_ (.I(_020_),
    .Z(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _270_ (.I0(\cm_inst.cc_inst.out_notouch_[192] ),
    .I1(\cm_inst.cc_inst.out_notouch_[200] ),
    .S(_041_),
    .Z(_042_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _271_ (.A1(\cm_inst.cc_inst.out_notouch_[208] ),
    .A2(_040_),
    .B1(_042_),
    .B2(_037_),
    .ZN(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _272_ (.I(_029_),
    .Z(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _273_ (.I(\cm_inst.page[3] ),
    .Z(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _274_ (.A1(_044_),
    .A2(_045_),
    .ZN(_046_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _275_ (.I(_017_),
    .Z(_047_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _276_ (.I(_019_),
    .Z(_048_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _277_ (.I0(\cm_inst.cc_inst.out_notouch_[160] ),
    .I1(\cm_inst.cc_inst.out_notouch_[168] ),
    .I2(\cm_inst.cc_inst.out_notouch_[176] ),
    .I3(\cm_inst.cc_inst.out_notouch_[184] ),
    .S0(_048_),
    .S1(_023_),
    .Z(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _278_ (.I0(\cm_inst.cc_inst.out_notouch_[128] ),
    .I1(\cm_inst.cc_inst.out_notouch_[136] ),
    .I2(\cm_inst.cc_inst.out_notouch_[144] ),
    .I3(\cm_inst.cc_inst.out_notouch_[152] ),
    .S0(_048_),
    .S1(_023_),
    .Z(_050_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _279_ (.I(_044_),
    .Z(_051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _280_ (.I0(_049_),
    .I1(_050_),
    .S(_051_),
    .Z(_052_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _281_ (.A1(_034_),
    .A2(_052_),
    .ZN(_053_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _282_ (.A1(_043_),
    .A2(_046_),
    .B(_047_),
    .C(_053_),
    .ZN(_054_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _283_ (.I(\cm_inst.page[5] ),
    .ZN(_055_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _284_ (.A1(_018_),
    .A2(_035_),
    .B(_054_),
    .C(_055_),
    .ZN(_056_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _285_ (.A1(\ro_inst.counter[0] ),
    .A2(\ro_inst.enable ),
    .ZN(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _286_ (.A1(_016_),
    .A2(_056_),
    .B(_057_),
    .ZN(out[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _287_ (.I(\cm_inst.page[5] ),
    .Z(_058_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _288_ (.I(\cm_inst.page[4] ),
    .Z(_059_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _289_ (.I(\cm_inst.page[0] ),
    .Z(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _290_ (.I(\cm_inst.page[1] ),
    .Z(_061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _291_ (.I0(\cm_inst.cc_inst.out_notouch_[97] ),
    .I1(\cm_inst.cc_inst.out_notouch_[105] ),
    .I2(\cm_inst.cc_inst.out_notouch_[113] ),
    .I3(\cm_inst.cc_inst.out_notouch_[121] ),
    .S0(_060_),
    .S1(_061_),
    .Z(_062_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _292_ (.I(\cm_inst.page[1] ),
    .Z(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _293_ (.I(_063_),
    .Z(_064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _294_ (.I0(\cm_inst.cc_inst.out_notouch_[65] ),
    .I1(\cm_inst.cc_inst.out_notouch_[73] ),
    .I2(\cm_inst.cc_inst.out_notouch_[81] ),
    .I3(\cm_inst.cc_inst.out_notouch_[89] ),
    .S0(_060_),
    .S1(_064_),
    .Z(_065_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _295_ (.I(_029_),
    .Z(_066_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _296_ (.I0(_062_),
    .I1(_065_),
    .S(_066_),
    .Z(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _297_ (.I0(\cm_inst.cc_inst.out_notouch_[33] ),
    .I1(\cm_inst.cc_inst.out_notouch_[41] ),
    .I2(\cm_inst.cc_inst.out_notouch_[49] ),
    .I3(\cm_inst.cc_inst.out_notouch_[57] ),
    .S0(_060_),
    .S1(_061_),
    .Z(_068_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _298_ (.I(\cm_inst.page[0] ),
    .Z(_069_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _299_ (.I(_069_),
    .Z(_070_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _300_ (.I0(\cm_inst.cc_inst.out_notouch_[1] ),
    .I1(\cm_inst.cc_inst.out_notouch_[9] ),
    .I2(\cm_inst.cc_inst.out_notouch_[17] ),
    .I3(\cm_inst.cc_inst.out_notouch_[25] ),
    .S0(_070_),
    .S1(_064_),
    .Z(_071_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _301_ (.I0(_068_),
    .I1(_071_),
    .S(_066_),
    .Z(_072_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _302_ (.I0(_067_),
    .I1(_072_),
    .S(_033_),
    .Z(_073_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _303_ (.A1(_059_),
    .A2(_073_),
    .ZN(_074_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _304_ (.I(_032_),
    .Z(_075_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _305_ (.I(_075_),
    .Z(_076_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _306_ (.I0(\cm_inst.cc_inst.out_notouch_[161] ),
    .I1(\cm_inst.cc_inst.out_notouch_[169] ),
    .I2(\cm_inst.cc_inst.out_notouch_[177] ),
    .I3(\cm_inst.cc_inst.out_notouch_[185] ),
    .S0(_048_),
    .S1(_023_),
    .Z(_077_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _307_ (.I(_022_),
    .Z(_078_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _308_ (.I0(\cm_inst.cc_inst.out_notouch_[129] ),
    .I1(\cm_inst.cc_inst.out_notouch_[137] ),
    .I2(\cm_inst.cc_inst.out_notouch_[145] ),
    .I3(\cm_inst.cc_inst.out_notouch_[153] ),
    .S0(_020_),
    .S1(_078_),
    .Z(_079_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _309_ (.I0(_077_),
    .I1(_079_),
    .S(_051_),
    .Z(_080_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _310_ (.I(_078_),
    .Z(_081_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _311_ (.I(_048_),
    .ZN(_082_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _312_ (.I(_082_),
    .Z(_083_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _313_ (.A1(_081_),
    .A2(_083_),
    .A3(\cm_inst.cc_inst.out_notouch_[209] ),
    .ZN(_084_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _314_ (.I(_019_),
    .Z(_085_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _315_ (.I0(\cm_inst.cc_inst.out_notouch_[193] ),
    .I1(\cm_inst.cc_inst.out_notouch_[201] ),
    .S(_085_),
    .Z(_086_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _316_ (.A1(_037_),
    .A2(_086_),
    .ZN(_087_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _317_ (.A1(_084_),
    .A2(_087_),
    .B(_046_),
    .ZN(_088_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _318_ (.I(\cm_inst.page[4] ),
    .ZN(_089_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _319_ (.A1(_076_),
    .A2(_080_),
    .B(_088_),
    .C(_089_),
    .ZN(_090_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _320_ (.A1(_058_),
    .A2(_074_),
    .A3(_090_),
    .ZN(_091_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _321_ (.I0(_091_),
    .I1(\ro_inst.counter[1] ),
    .S(_016_),
    .Z(out[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _322_ (.I0(\cm_inst.cc_inst.out_notouch_[162] ),
    .I1(\cm_inst.cc_inst.out_notouch_[170] ),
    .I2(\cm_inst.cc_inst.out_notouch_[178] ),
    .I3(\cm_inst.cc_inst.out_notouch_[186] ),
    .S0(_020_),
    .S1(_078_),
    .Z(_092_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _323_ (.I(\cm_inst.page[0] ),
    .Z(_093_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _324_ (.I(_093_),
    .Z(_094_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _325_ (.I(_022_),
    .Z(_095_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _326_ (.I0(\cm_inst.cc_inst.out_notouch_[130] ),
    .I1(\cm_inst.cc_inst.out_notouch_[138] ),
    .I2(\cm_inst.cc_inst.out_notouch_[146] ),
    .I3(\cm_inst.cc_inst.out_notouch_[154] ),
    .S0(_094_),
    .S1(_095_),
    .Z(_096_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _327_ (.I0(_092_),
    .I1(_096_),
    .S(_051_),
    .Z(_097_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _328_ (.I(_061_),
    .Z(_098_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _329_ (.A1(_098_),
    .A2(_046_),
    .ZN(_099_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _330_ (.I0(\cm_inst.cc_inst.out_notouch_[194] ),
    .I1(\cm_inst.cc_inst.out_notouch_[202] ),
    .S(_041_),
    .Z(_100_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _331_ (.A1(_076_),
    .A2(_097_),
    .B1(_099_),
    .B2(_100_),
    .ZN(_101_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _332_ (.I(_082_),
    .Z(_102_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _333_ (.I(_093_),
    .Z(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _334_ (.A1(_103_),
    .A2(\cm_inst.cc_inst.out_notouch_[90] ),
    .Z(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _335_ (.I(_036_),
    .Z(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _336_ (.A1(_102_),
    .A2(\cm_inst.cc_inst.out_notouch_[82] ),
    .B(_104_),
    .C(_105_),
    .ZN(_106_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _337_ (.I(_098_),
    .Z(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _338_ (.I(_060_),
    .Z(_108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _339_ (.I0(\cm_inst.cc_inst.out_notouch_[66] ),
    .I1(\cm_inst.cc_inst.out_notouch_[74] ),
    .S(_108_),
    .Z(_109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _340_ (.A1(_107_),
    .A2(_109_),
    .B(_031_),
    .ZN(_110_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _341_ (.I(\cm_inst.page[2] ),
    .Z(_111_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _342_ (.I(_111_),
    .Z(_112_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _343_ (.I(_022_),
    .Z(_113_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _344_ (.I0(\cm_inst.cc_inst.out_notouch_[98] ),
    .I1(\cm_inst.cc_inst.out_notouch_[106] ),
    .I2(\cm_inst.cc_inst.out_notouch_[114] ),
    .I3(\cm_inst.cc_inst.out_notouch_[122] ),
    .S0(_085_),
    .S1(_113_),
    .Z(_114_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _345_ (.A1(_112_),
    .A2(_114_),
    .ZN(_115_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _346_ (.A1(_106_),
    .A2(_110_),
    .B(_045_),
    .C(_115_),
    .ZN(_116_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _347_ (.A1(_038_),
    .A2(\cm_inst.cc_inst.out_notouch_[26] ),
    .Z(_117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _348_ (.A1(_083_),
    .A2(\cm_inst.cc_inst.out_notouch_[18] ),
    .B(_117_),
    .C(_036_),
    .ZN(_118_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _349_ (.I(_093_),
    .Z(_119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _350_ (.I0(\cm_inst.cc_inst.out_notouch_[2] ),
    .I1(\cm_inst.cc_inst.out_notouch_[10] ),
    .S(_119_),
    .Z(_120_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _351_ (.I(_044_),
    .Z(_121_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _352_ (.A1(_081_),
    .A2(_120_),
    .B(_121_),
    .ZN(_122_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _353_ (.I(_069_),
    .Z(_123_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _354_ (.I(_063_),
    .Z(_124_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _355_ (.I0(\cm_inst.cc_inst.out_notouch_[34] ),
    .I1(\cm_inst.cc_inst.out_notouch_[42] ),
    .I2(\cm_inst.cc_inst.out_notouch_[50] ),
    .I3(\cm_inst.cc_inst.out_notouch_[58] ),
    .S0(_123_),
    .S1(_124_),
    .Z(_125_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _356_ (.A1(_111_),
    .A2(_125_),
    .ZN(_126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _357_ (.A1(_118_),
    .A2(_122_),
    .B(_075_),
    .C(_126_),
    .ZN(_127_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _358_ (.A1(_116_),
    .A2(_127_),
    .B(_017_),
    .ZN(_128_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _359_ (.I(\cm_inst.page[5] ),
    .Z(_129_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _360_ (.A1(_047_),
    .A2(_101_),
    .B(_128_),
    .C(_129_),
    .ZN(_130_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _361_ (.I0(_130_),
    .I1(\ro_inst.counter[2] ),
    .S(_016_),
    .Z(out[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _362_ (.I0(\cm_inst.cc_inst.out_notouch_[163] ),
    .I1(\cm_inst.cc_inst.out_notouch_[171] ),
    .I2(\cm_inst.cc_inst.out_notouch_[179] ),
    .I3(\cm_inst.cc_inst.out_notouch_[187] ),
    .S0(_094_),
    .S1(_078_),
    .Z(_131_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _363_ (.I0(\cm_inst.cc_inst.out_notouch_[131] ),
    .I1(\cm_inst.cc_inst.out_notouch_[139] ),
    .I2(\cm_inst.cc_inst.out_notouch_[147] ),
    .I3(\cm_inst.cc_inst.out_notouch_[155] ),
    .S0(_094_),
    .S1(_095_),
    .Z(_132_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _364_ (.I(_044_),
    .Z(_133_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _365_ (.I0(_131_),
    .I1(_132_),
    .S(_133_),
    .Z(_134_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _366_ (.I0(\cm_inst.cc_inst.out_notouch_[195] ),
    .I1(\cm_inst.cc_inst.out_notouch_[203] ),
    .S(_041_),
    .Z(_135_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _367_ (.A1(_076_),
    .A2(_134_),
    .B1(_135_),
    .B2(_099_),
    .ZN(_136_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _368_ (.I0(\cm_inst.cc_inst.out_notouch_[99] ),
    .I1(\cm_inst.cc_inst.out_notouch_[107] ),
    .I2(\cm_inst.cc_inst.out_notouch_[115] ),
    .I3(\cm_inst.cc_inst.out_notouch_[123] ),
    .S0(_070_),
    .S1(_064_),
    .Z(_137_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _369_ (.I(_063_),
    .Z(_138_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _370_ (.I0(\cm_inst.cc_inst.out_notouch_[67] ),
    .I1(\cm_inst.cc_inst.out_notouch_[75] ),
    .I2(\cm_inst.cc_inst.out_notouch_[83] ),
    .I3(\cm_inst.cc_inst.out_notouch_[91] ),
    .S0(_070_),
    .S1(_138_),
    .Z(_139_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _371_ (.I0(_137_),
    .I1(_139_),
    .S(_066_),
    .Z(_140_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _372_ (.I0(\cm_inst.cc_inst.out_notouch_[35] ),
    .I1(\cm_inst.cc_inst.out_notouch_[43] ),
    .I2(\cm_inst.cc_inst.out_notouch_[51] ),
    .I3(\cm_inst.cc_inst.out_notouch_[59] ),
    .S0(_070_),
    .S1(_064_),
    .Z(_141_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _373_ (.I(_069_),
    .Z(_142_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _374_ (.I0(\cm_inst.cc_inst.out_notouch_[3] ),
    .I1(\cm_inst.cc_inst.out_notouch_[11] ),
    .I2(\cm_inst.cc_inst.out_notouch_[19] ),
    .I3(\cm_inst.cc_inst.out_notouch_[27] ),
    .S0(_142_),
    .S1(_138_),
    .Z(_143_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _375_ (.I0(_141_),
    .I1(_143_),
    .S(_066_),
    .Z(_144_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _376_ (.I0(_140_),
    .I1(_144_),
    .S(_033_),
    .Z(_145_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _377_ (.A1(_059_),
    .A2(_145_),
    .ZN(_146_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _378_ (.A1(_047_),
    .A2(_136_),
    .B(_146_),
    .C(_129_),
    .ZN(_147_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _379_ (.I(\ro_inst.enable ),
    .Z(_148_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _380_ (.I0(_147_),
    .I1(\ro_inst.counter[3] ),
    .S(_148_),
    .Z(out[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _381_ (.I0(\cm_inst.cc_inst.out_notouch_[164] ),
    .I1(\cm_inst.cc_inst.out_notouch_[172] ),
    .I2(\cm_inst.cc_inst.out_notouch_[180] ),
    .I3(\cm_inst.cc_inst.out_notouch_[188] ),
    .S0(_094_),
    .S1(_095_),
    .Z(_149_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _382_ (.I(_093_),
    .Z(_150_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _383_ (.I(_061_),
    .Z(_151_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _384_ (.I0(\cm_inst.cc_inst.out_notouch_[132] ),
    .I1(\cm_inst.cc_inst.out_notouch_[140] ),
    .I2(\cm_inst.cc_inst.out_notouch_[148] ),
    .I3(\cm_inst.cc_inst.out_notouch_[156] ),
    .S0(_150_),
    .S1(_151_),
    .Z(_152_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _385_ (.I0(_149_),
    .I1(_152_),
    .S(_133_),
    .Z(_153_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _386_ (.I0(\cm_inst.cc_inst.out_notouch_[196] ),
    .I1(\cm_inst.cc_inst.out_notouch_[204] ),
    .S(_041_),
    .Z(_154_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _387_ (.I(_099_),
    .Z(_155_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _388_ (.A1(_076_),
    .A2(_153_),
    .B1(_154_),
    .B2(_155_),
    .ZN(_156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _389_ (.A1(_103_),
    .A2(\cm_inst.cc_inst.out_notouch_[92] ),
    .Z(_157_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _390_ (.A1(_102_),
    .A2(\cm_inst.cc_inst.out_notouch_[84] ),
    .B(_157_),
    .C(_105_),
    .ZN(_158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _391_ (.I0(\cm_inst.cc_inst.out_notouch_[68] ),
    .I1(\cm_inst.cc_inst.out_notouch_[76] ),
    .S(_108_),
    .Z(_159_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _392_ (.A1(_107_),
    .A2(_159_),
    .B(_031_),
    .ZN(_160_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _393_ (.I0(\cm_inst.cc_inst.out_notouch_[100] ),
    .I1(\cm_inst.cc_inst.out_notouch_[108] ),
    .I2(\cm_inst.cc_inst.out_notouch_[116] ),
    .I3(\cm_inst.cc_inst.out_notouch_[124] ),
    .S0(_085_),
    .S1(_113_),
    .Z(_161_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _394_ (.A1(_112_),
    .A2(_161_),
    .ZN(_162_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _395_ (.A1(_158_),
    .A2(_160_),
    .B(_045_),
    .C(_162_),
    .ZN(_163_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _396_ (.A1(_038_),
    .A2(\cm_inst.cc_inst.out_notouch_[28] ),
    .Z(_164_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _397_ (.A1(_083_),
    .A2(\cm_inst.cc_inst.out_notouch_[20] ),
    .B(_164_),
    .C(_105_),
    .ZN(_165_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _398_ (.I0(\cm_inst.cc_inst.out_notouch_[4] ),
    .I1(\cm_inst.cc_inst.out_notouch_[12] ),
    .S(_119_),
    .Z(_166_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _399_ (.A1(_081_),
    .A2(_166_),
    .B(_121_),
    .ZN(_167_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _400_ (.I0(\cm_inst.cc_inst.out_notouch_[36] ),
    .I1(\cm_inst.cc_inst.out_notouch_[44] ),
    .I2(\cm_inst.cc_inst.out_notouch_[52] ),
    .I3(\cm_inst.cc_inst.out_notouch_[60] ),
    .S0(_123_),
    .S1(_124_),
    .Z(_168_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _401_ (.A1(_111_),
    .A2(_168_),
    .ZN(_169_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _402_ (.A1(_165_),
    .A2(_167_),
    .B(_034_),
    .C(_169_),
    .ZN(_170_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _403_ (.A1(_163_),
    .A2(_170_),
    .B(_017_),
    .ZN(_171_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _404_ (.A1(_018_),
    .A2(_156_),
    .B(_171_),
    .C(_129_),
    .ZN(_172_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _405_ (.I0(_172_),
    .I1(\ro_inst.counter[4] ),
    .S(_148_),
    .Z(out[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _406_ (.I(_075_),
    .Z(_173_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _407_ (.I0(\cm_inst.cc_inst.out_notouch_[165] ),
    .I1(\cm_inst.cc_inst.out_notouch_[173] ),
    .I2(\cm_inst.cc_inst.out_notouch_[181] ),
    .I3(\cm_inst.cc_inst.out_notouch_[189] ),
    .S0(_150_),
    .S1(_151_),
    .Z(_174_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _408_ (.I0(\cm_inst.cc_inst.out_notouch_[133] ),
    .I1(\cm_inst.cc_inst.out_notouch_[141] ),
    .I2(\cm_inst.cc_inst.out_notouch_[149] ),
    .I3(\cm_inst.cc_inst.out_notouch_[157] ),
    .S0(_119_),
    .S1(_151_),
    .Z(_175_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _409_ (.I0(_174_),
    .I1(_175_),
    .S(_133_),
    .Z(_176_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _410_ (.I0(\cm_inst.cc_inst.out_notouch_[197] ),
    .I1(\cm_inst.cc_inst.out_notouch_[205] ),
    .S(_039_),
    .Z(_177_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _411_ (.A1(_173_),
    .A2(_176_),
    .B1(_177_),
    .B2(_155_),
    .ZN(_178_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _412_ (.I0(\cm_inst.cc_inst.out_notouch_[101] ),
    .I1(\cm_inst.cc_inst.out_notouch_[109] ),
    .I2(\cm_inst.cc_inst.out_notouch_[117] ),
    .I3(\cm_inst.cc_inst.out_notouch_[125] ),
    .S0(_142_),
    .S1(_138_),
    .Z(_179_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _413_ (.I(_063_),
    .Z(_180_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _414_ (.I0(\cm_inst.cc_inst.out_notouch_[69] ),
    .I1(\cm_inst.cc_inst.out_notouch_[77] ),
    .I2(\cm_inst.cc_inst.out_notouch_[85] ),
    .I3(\cm_inst.cc_inst.out_notouch_[93] ),
    .S0(_142_),
    .S1(_180_),
    .Z(_181_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _415_ (.I0(_179_),
    .I1(_181_),
    .S(_030_),
    .Z(_182_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _416_ (.I0(\cm_inst.cc_inst.out_notouch_[37] ),
    .I1(\cm_inst.cc_inst.out_notouch_[45] ),
    .I2(\cm_inst.cc_inst.out_notouch_[53] ),
    .I3(\cm_inst.cc_inst.out_notouch_[61] ),
    .S0(_142_),
    .S1(_138_),
    .Z(_183_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _417_ (.I(_069_),
    .Z(_184_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _418_ (.I0(\cm_inst.cc_inst.out_notouch_[5] ),
    .I1(\cm_inst.cc_inst.out_notouch_[13] ),
    .I2(\cm_inst.cc_inst.out_notouch_[21] ),
    .I3(\cm_inst.cc_inst.out_notouch_[29] ),
    .S0(_184_),
    .S1(_180_),
    .Z(_185_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _419_ (.I0(_183_),
    .I1(_185_),
    .S(_030_),
    .Z(_186_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _420_ (.I0(_182_),
    .I1(_186_),
    .S(_033_),
    .Z(_187_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _421_ (.A1(_059_),
    .A2(_187_),
    .ZN(_188_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _422_ (.A1(_018_),
    .A2(_178_),
    .B(_188_),
    .C(_058_),
    .ZN(_189_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _423_ (.I0(_189_),
    .I1(\ro_inst.counter[5] ),
    .S(_148_),
    .Z(out[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _424_ (.I0(\cm_inst.cc_inst.out_notouch_[166] ),
    .I1(\cm_inst.cc_inst.out_notouch_[174] ),
    .I2(\cm_inst.cc_inst.out_notouch_[182] ),
    .I3(\cm_inst.cc_inst.out_notouch_[190] ),
    .S0(_150_),
    .S1(_095_),
    .Z(_190_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _425_ (.I0(\cm_inst.cc_inst.out_notouch_[134] ),
    .I1(\cm_inst.cc_inst.out_notouch_[142] ),
    .I2(\cm_inst.cc_inst.out_notouch_[150] ),
    .I3(\cm_inst.cc_inst.out_notouch_[158] ),
    .S0(_150_),
    .S1(_151_),
    .Z(_191_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _426_ (.I0(_190_),
    .I1(_191_),
    .S(_133_),
    .Z(_192_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _427_ (.I0(\cm_inst.cc_inst.out_notouch_[198] ),
    .I1(\cm_inst.cc_inst.out_notouch_[206] ),
    .S(_039_),
    .Z(_193_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _428_ (.A1(_173_),
    .A2(_192_),
    .B1(_193_),
    .B2(_155_),
    .ZN(_194_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _429_ (.A1(_103_),
    .A2(\cm_inst.cc_inst.out_notouch_[94] ),
    .Z(_195_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _430_ (.A1(_102_),
    .A2(\cm_inst.cc_inst.out_notouch_[86] ),
    .B(_195_),
    .C(_037_),
    .ZN(_196_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _431_ (.I0(\cm_inst.cc_inst.out_notouch_[70] ),
    .I1(\cm_inst.cc_inst.out_notouch_[78] ),
    .S(_038_),
    .Z(_197_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _432_ (.A1(_107_),
    .A2(_197_),
    .B(_031_),
    .ZN(_198_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _433_ (.I0(\cm_inst.cc_inst.out_notouch_[102] ),
    .I1(\cm_inst.cc_inst.out_notouch_[110] ),
    .I2(\cm_inst.cc_inst.out_notouch_[118] ),
    .I3(\cm_inst.cc_inst.out_notouch_[126] ),
    .S0(_085_),
    .S1(_113_),
    .Z(_199_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _434_ (.A1(_112_),
    .A2(_199_),
    .ZN(_200_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _435_ (.A1(_196_),
    .A2(_198_),
    .B(_045_),
    .C(_200_),
    .ZN(_201_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _436_ (.A1(_103_),
    .A2(\cm_inst.cc_inst.out_notouch_[30] ),
    .Z(_202_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _437_ (.A1(_083_),
    .A2(\cm_inst.cc_inst.out_notouch_[22] ),
    .B(_202_),
    .C(_105_),
    .ZN(_203_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _438_ (.I0(\cm_inst.cc_inst.out_notouch_[6] ),
    .I1(\cm_inst.cc_inst.out_notouch_[14] ),
    .S(_119_),
    .Z(_204_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _439_ (.A1(_081_),
    .A2(_204_),
    .B(_121_),
    .ZN(_205_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _440_ (.I0(\cm_inst.cc_inst.out_notouch_[38] ),
    .I1(\cm_inst.cc_inst.out_notouch_[46] ),
    .I2(\cm_inst.cc_inst.out_notouch_[54] ),
    .I3(\cm_inst.cc_inst.out_notouch_[62] ),
    .S0(_123_),
    .S1(_113_),
    .Z(_206_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _441_ (.A1(_111_),
    .A2(_206_),
    .ZN(_207_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _442_ (.A1(_203_),
    .A2(_205_),
    .B(_034_),
    .C(_207_),
    .ZN(_208_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _443_ (.A1(_201_),
    .A2(_208_),
    .B(_059_),
    .ZN(_209_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _444_ (.A1(_018_),
    .A2(_194_),
    .B(_209_),
    .C(_058_),
    .ZN(_210_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _445_ (.I0(_210_),
    .I1(\ro_inst.counter[34] ),
    .S(_148_),
    .Z(out[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _446_ (.I0(\cm_inst.cc_inst.out_notouch_[103] ),
    .I1(\cm_inst.cc_inst.out_notouch_[111] ),
    .I2(\cm_inst.cc_inst.out_notouch_[119] ),
    .I3(\cm_inst.cc_inst.out_notouch_[127] ),
    .S0(_184_),
    .S1(_180_),
    .Z(_211_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _447_ (.I0(\cm_inst.cc_inst.out_notouch_[71] ),
    .I1(\cm_inst.cc_inst.out_notouch_[79] ),
    .I2(\cm_inst.cc_inst.out_notouch_[87] ),
    .I3(\cm_inst.cc_inst.out_notouch_[95] ),
    .S0(_184_),
    .S1(_124_),
    .Z(_212_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _448_ (.I0(_211_),
    .I1(_212_),
    .S(_030_),
    .Z(_213_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _449_ (.I0(\cm_inst.cc_inst.out_notouch_[39] ),
    .I1(\cm_inst.cc_inst.out_notouch_[47] ),
    .I2(\cm_inst.cc_inst.out_notouch_[55] ),
    .I3(\cm_inst.cc_inst.out_notouch_[63] ),
    .S0(_184_),
    .S1(_180_),
    .Z(_214_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _450_ (.I0(\cm_inst.cc_inst.out_notouch_[7] ),
    .I1(\cm_inst.cc_inst.out_notouch_[15] ),
    .I2(\cm_inst.cc_inst.out_notouch_[23] ),
    .I3(\cm_inst.cc_inst.out_notouch_[31] ),
    .S0(_123_),
    .S1(_124_),
    .Z(_215_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _451_ (.I0(_214_),
    .I1(_215_),
    .S(_051_),
    .Z(_216_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _452_ (.I0(_213_),
    .I1(_216_),
    .S(_075_),
    .Z(_217_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _453_ (.A1(_047_),
    .A2(_217_),
    .ZN(_218_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _454_ (.I0(\cm_inst.cc_inst.out_notouch_[167] ),
    .I1(\cm_inst.cc_inst.out_notouch_[175] ),
    .I2(\cm_inst.cc_inst.out_notouch_[183] ),
    .I3(\cm_inst.cc_inst.out_notouch_[191] ),
    .S0(_108_),
    .S1(_098_),
    .Z(_219_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _455_ (.I0(\cm_inst.cc_inst.out_notouch_[135] ),
    .I1(\cm_inst.cc_inst.out_notouch_[143] ),
    .I2(\cm_inst.cc_inst.out_notouch_[151] ),
    .I3(\cm_inst.cc_inst.out_notouch_[159] ),
    .S0(_108_),
    .S1(_098_),
    .Z(_220_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _456_ (.I0(_219_),
    .I1(_220_),
    .S(_121_),
    .Z(_221_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _457_ (.A1(_102_),
    .A2(\cm_inst.cc_inst.out_notouch_[199] ),
    .Z(_222_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _458_ (.A1(_173_),
    .A2(_221_),
    .B1(_222_),
    .B2(_155_),
    .C(_089_),
    .ZN(_223_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _459_ (.A1(_058_),
    .A2(_218_),
    .A3(_223_),
    .ZN(_224_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _460_ (.I0(_224_),
    .I1(\ro_inst.saved_signal ),
    .S(\ro_inst.enable ),
    .Z(out[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _461_ (.I(\ro_sel[0] ),
    .Z(_225_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _462_ (.I(\ro_sel[0] ),
    .ZN(_226_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__or4_1 _463_ (.A1(_129_),
    .A2(_226_),
    .A3(_074_),
    .A4(_090_),
    .Z(_227_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _464_ (.A1(_225_),
    .A2(_056_),
    .B(_227_),
    .ZN(_228_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _465_ (.I0(_172_),
    .I1(_189_),
    .S(_225_),
    .Z(_229_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _466_ (.I0(_130_),
    .I1(_147_),
    .S(\ro_sel[0] ),
    .Z(_230_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _467_ (.I0(_210_),
    .I1(_224_),
    .S(_225_),
    .Z(_231_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 _468_ (.I0(_228_),
    .I1(_229_),
    .I2(_230_),
    .I3(_231_),
    .S0(\ro_sel[2] ),
    .S1(\ro_sel[1] ),
    .Z(_232_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _469_ (.I(_232_),
    .Z(\ro_inst.signal ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _470_ (.I(in[5]),
    .ZN(_233_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _471_ (.I(in[6]),
    .ZN(_234_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _472_ (.I(in[7]),
    .ZN(_235_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _473_ (.A1(_233_),
    .A2(_234_),
    .A3(_235_),
    .B(in[1]),
    .ZN(_236_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _474_ (.I(_236_),
    .Z(_237_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _475_ (.I0(in[2]),
    .I1(_039_),
    .S(_237_),
    .Z(_000_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _476_ (.I0(in[3]),
    .I1(_107_),
    .S(_236_),
    .Z(_001_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _477_ (.I0(in[4]),
    .I1(_112_),
    .S(_236_),
    .Z(_002_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _478_ (.I(in[1]),
    .Z(_238_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _479_ (.I(_238_),
    .Z(_239_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _480_ (.A1(_233_),
    .A2(_239_),
    .B1(_173_),
    .B2(_237_),
    .ZN(_003_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _481_ (.A1(_234_),
    .A2(_239_),
    .B1(_089_),
    .B2(_237_),
    .ZN(_004_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _482_ (.A1(_235_),
    .A2(_239_),
    .B1(_055_),
    .B2(_237_),
    .ZN(_005_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _483_ (.I0(in[2]),
    .I1(\cm_inst.cc_inst.in[0] ),
    .S(_239_),
    .Z(_006_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 _484_ (.I(_238_),
    .Z(_240_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _485_ (.I0(in[3]),
    .I1(\cm_inst.cc_inst.in[1] ),
    .S(_240_),
    .Z(_007_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _486_ (.I0(in[4]),
    .I1(\cm_inst.cc_inst.in[2] ),
    .S(_240_),
    .Z(_008_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _487_ (.I0(in[5]),
    .I1(\cm_inst.cc_inst.in[3] ),
    .S(_240_),
    .Z(_009_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _488_ (.I0(in[6]),
    .I1(\cm_inst.cc_inst.in[4] ),
    .S(_240_),
    .Z(_010_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _489_ (.I0(in[7]),
    .I1(\cm_inst.cc_inst.in[5] ),
    .S(_238_),
    .Z(_011_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _490_ (.A1(_238_),
    .A2(_016_),
    .B(_236_),
    .ZN(_241_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _491_ (.I(_241_),
    .ZN(_012_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _492_ (.A1(in[5]),
    .A2(in[6]),
    .A3(in[7]),
    .A4(in[1]),
    .ZN(_242_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _493_ (.I0(in[2]),
    .I1(_225_),
    .S(_242_),
    .Z(_013_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _494_ (.I0(in[3]),
    .I1(\ro_sel[1] ),
    .S(_242_),
    .Z(_014_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _495_ (.I0(in[4]),
    .I1(\ro_sel[2] ),
    .S(_242_),
    .Z(_015_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _496_ (.D(_000_),
    .CLK(in[0]),
    .Q(\cm_inst.page[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _497_ (.D(_001_),
    .CLK(in[0]),
    .Q(\cm_inst.page[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _498_ (.D(_002_),
    .CLK(in[0]),
    .Q(\cm_inst.page[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _499_ (.D(_003_),
    .CLK(in[0]),
    .Q(\cm_inst.page[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _500_ (.D(_004_),
    .CLK(in[0]),
    .Q(\cm_inst.page[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _501_ (.D(_005_),
    .CLK(in[0]),
    .Q(\cm_inst.page[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _502_ (.D(_006_),
    .CLK(in[0]),
    .Q(\cm_inst.cc_inst.in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _503_ (.D(_007_),
    .CLK(in[0]),
    .Q(\cm_inst.cc_inst.in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _504_ (.D(_008_),
    .CLK(in[0]),
    .Q(\cm_inst.cc_inst.in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _505_ (.D(_009_),
    .CLK(in[0]),
    .Q(\cm_inst.cc_inst.in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _506_ (.D(_010_),
    .CLK(in[0]),
    .Q(\cm_inst.cc_inst.in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _507_ (.D(_011_),
    .CLK(in[0]),
    .Q(\cm_inst.cc_inst.in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _508_ (.D(_012_),
    .CLK(in[0]),
    .Q(\ro_inst.enable ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _509_ (.D(_013_),
    .CLK(in[0]),
    .Q(\ro_sel[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _510_ (.D(_014_),
    .CLK(in[0]),
    .Q(\ro_sel[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _511_ (.D(_015_),
    .CLK(in[0]),
    .Q(\ro_sel[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _512_ (.ZN(_243_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _513_ (.ZN(out[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _514_ (.ZN(out[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _515_ (.ZN(out[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _516_ (.ZN(out[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 \cm_inst.cc_inst.addf_1_inst  (.A(\cm_inst.cc_inst.in[0] ),
    .B(\cm_inst.cc_inst.in[1] ),
    .CI(\cm_inst.cc_inst.in[2] ),
    .CO(\cm_inst.cc_inst.out_notouch_[105] ),
    .S(\cm_inst.cc_inst.out_notouch_[106] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 \cm_inst.cc_inst.addf_2_inst  (.A(\cm_inst.cc_inst.in[0] ),
    .B(\cm_inst.cc_inst.in[1] ),
    .CI(\cm_inst.cc_inst.in[2] ),
    .CO(\cm_inst.cc_inst.out_notouch_[107] ),
    .S(\cm_inst.cc_inst.out_notouch_[108] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__addf_4 \cm_inst.cc_inst.addf_4_inst  (.A(\cm_inst.cc_inst.in[0] ),
    .B(\cm_inst.cc_inst.in[1] ),
    .CI(\cm_inst.cc_inst.in[2] ),
    .CO(\cm_inst.cc_inst.out_notouch_[109] ),
    .S(\cm_inst.cc_inst.out_notouch_[110] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 \cm_inst.cc_inst.addh_1_inst  (.A(\cm_inst.cc_inst.in[0] ),
    .B(\cm_inst.cc_inst.in[1] ),
    .CO(\cm_inst.cc_inst.out_notouch_[111] ),
    .S(\cm_inst.cc_inst.out_notouch_[112] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 \cm_inst.cc_inst.addh_2_inst  (.A(\cm_inst.cc_inst.in[0] ),
    .B(\cm_inst.cc_inst.in[1] ),
    .CO(\cm_inst.cc_inst.out_notouch_[113] ),
    .S(\cm_inst.cc_inst.out_notouch_[114] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 \cm_inst.cc_inst.addh_4_inst  (.A(\cm_inst.cc_inst.in[0] ),
    .B(\cm_inst.cc_inst.in[1] ),
    .CO(\cm_inst.cc_inst.out_notouch_[115] ),
    .S(\cm_inst.cc_inst.out_notouch_[116] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 \cm_inst.cc_inst.and2_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[18] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 \cm_inst.cc_inst.and2_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[19] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 \cm_inst.cc_inst.and2_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[20] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 \cm_inst.cc_inst.and3_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[21] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 \cm_inst.cc_inst.and3_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[22] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 \cm_inst.cc_inst.and3_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[23] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and4_1 \cm_inst.cc_inst.and4_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .Z(\cm_inst.cc_inst.out_notouch_[24] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 \cm_inst.cc_inst.and4_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .Z(\cm_inst.cc_inst.out_notouch_[25] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 \cm_inst.cc_inst.and4_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .Z(\cm_inst.cc_inst.out_notouch_[26] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 \cm_inst.cc_inst.aoi211_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .C(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[72] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 \cm_inst.cc_inst.aoi211_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .C(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[73] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 \cm_inst.cc_inst.aoi211_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .C(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[74] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 \cm_inst.cc_inst.aoi21_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[66] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 \cm_inst.cc_inst.aoi21_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[67] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 \cm_inst.cc_inst.aoi21_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[68] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 \cm_inst.cc_inst.aoi221_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C(\cm_inst.cc_inst.in[4] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[75] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 \cm_inst.cc_inst.aoi221_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C(\cm_inst.cc_inst.in[4] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[76] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 \cm_inst.cc_inst.aoi221_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C(\cm_inst.cc_inst.in[4] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[77] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_1 \cm_inst.cc_inst.aoi222_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C1(\cm_inst.cc_inst.in[4] ),
    .C2(\cm_inst.cc_inst.in[5] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[78] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 \cm_inst.cc_inst.aoi222_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C1(\cm_inst.cc_inst.in[4] ),
    .C2(\cm_inst.cc_inst.in[5] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[79] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 \cm_inst.cc_inst.aoi222_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C1(\cm_inst.cc_inst.in[4] ),
    .C2(\cm_inst.cc_inst.in[5] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[80] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 \cm_inst.cc_inst.aoi22_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[69] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 \cm_inst.cc_inst.aoi22_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[70] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 \cm_inst.cc_inst.aoi22_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[71] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 \cm_inst.cc_inst.buf_12_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 \cm_inst.cc_inst.buf_16_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[8] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 \cm_inst.cc_inst.buf_1_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 \cm_inst.cc_inst.buf_20_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 \cm_inst.cc_inst.buf_2_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 \cm_inst.cc_inst.buf_3_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 \cm_inst.cc_inst.buf_4_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 \cm_inst.cc_inst.buf_8_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__bufz_12 \cm_inst.cc_inst.bufz_12_inst  (.EN(\cm_inst.cc_inst.in[4] ),
    .I(\cm_inst.cc_inst.in[5] ),
    .Z(\cm_inst.cc_inst.out_notouch_[172] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__bufz_16 \cm_inst.cc_inst.bufz_16_inst  (.EN(\cm_inst.cc_inst.in[0] ),
    .I(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[173] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__bufz_1 \cm_inst.cc_inst.bufz_1_inst  (.EN(\cm_inst.cc_inst.in[0] ),
    .I(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[171] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__bufz_2 \cm_inst.cc_inst.bufz_2_inst  (.EN(\cm_inst.cc_inst.in[2] ),
    .I(\cm_inst.cc_inst.in[3] ),
    .Z(\cm_inst.cc_inst.out_notouch_[171] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__bufz_3 \cm_inst.cc_inst.bufz_3_inst  (.EN(\cm_inst.cc_inst.in[4] ),
    .I(\cm_inst.cc_inst.in[5] ),
    .Z(\cm_inst.cc_inst.out_notouch_[171] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__bufz_4 \cm_inst.cc_inst.bufz_4_inst  (.EN(\cm_inst.cc_inst.in[0] ),
    .I(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[172] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__bufz_8 \cm_inst.cc_inst.bufz_8_inst  (.EN(\cm_inst.cc_inst.in[2] ),
    .I(\cm_inst.cc_inst.in[3] ),
    .Z(\cm_inst.cc_inst.out_notouch_[172] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 \cm_inst.cc_inst.clkbuf_12_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[193] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 \cm_inst.cc_inst.clkbuf_16_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[194] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 \cm_inst.cc_inst.clkbuf_1_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[188] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 \cm_inst.cc_inst.clkbuf_20_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[195] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 \cm_inst.cc_inst.clkbuf_2_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[189] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 \cm_inst.cc_inst.clkbuf_3_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[190] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 \cm_inst.cc_inst.clkbuf_4_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[191] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 \cm_inst.cc_inst.clkbuf_8_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[192] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 \cm_inst.cc_inst.clkinv_12_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[201] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 \cm_inst.cc_inst.clkinv_16_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[202] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 \cm_inst.cc_inst.clkinv_1_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[196] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 \cm_inst.cc_inst.clkinv_20_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[203] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 \cm_inst.cc_inst.clkinv_2_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[197] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 \cm_inst.cc_inst.clkinv_3_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[198] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 \cm_inst.cc_inst.clkinv_4_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[199] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 \cm_inst.cc_inst.clkinv_8_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[200] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnq_1 \cm_inst.cc_inst.dffnq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[135] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnq_2 \cm_inst.cc_inst.dffnq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[136] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnq_4 \cm_inst.cc_inst.dffnq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[137] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1 \cm_inst.cc_inst.dffnrnq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[138] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \cm_inst.cc_inst.dffnrnq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[139] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 \cm_inst.cc_inst.dffnrnq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[140] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 \cm_inst.cc_inst.dffnrsnq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[141] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2 \cm_inst.cc_inst.dffnrsnq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[142] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4 \cm_inst.cc_inst.dffnrsnq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[143] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1 \cm_inst.cc_inst.dffnsnq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SETN(\cm_inst.cc_inst.in[2] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[144] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 \cm_inst.cc_inst.dffnsnq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SETN(\cm_inst.cc_inst.in[2] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[145] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4 \cm_inst.cc_inst.dffnsnq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SETN(\cm_inst.cc_inst.in[2] ),
    .CLKN(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[146] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 \cm_inst.cc_inst.dffq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[147] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \cm_inst.cc_inst.dffq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[148] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \cm_inst.cc_inst.dffq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[149] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \cm_inst.cc_inst.dffrnq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[150] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cm_inst.cc_inst.dffrnq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[151] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \cm_inst.cc_inst.dffrnq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[152] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1 \cm_inst.cc_inst.dffrsnq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[153] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2 \cm_inst.cc_inst.dffrsnq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[154] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4 \cm_inst.cc_inst.dffrsnq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[155] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 \cm_inst.cc_inst.dffsnq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SETN(\cm_inst.cc_inst.in[2] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[156] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \cm_inst.cc_inst.dffsnq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SETN(\cm_inst.cc_inst.in[2] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[157] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \cm_inst.cc_inst.dffsnq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SETN(\cm_inst.cc_inst.in[2] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[158] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlya_1 \cm_inst.cc_inst.dlya_1_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[176] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 \cm_inst.cc_inst.dlya_2_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[177] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 \cm_inst.cc_inst.dlya_4_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[178] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_1 \cm_inst.cc_inst.dlyb_1_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[179] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 \cm_inst.cc_inst.dlyb_2_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[180] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_4 \cm_inst.cc_inst.dlyb_4_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[181] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_1 \cm_inst.cc_inst.dlyc_1_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[182] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 \cm_inst.cc_inst.dlyc_2_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[183] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_4 \cm_inst.cc_inst.dlyc_4_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[184] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlyd_1 \cm_inst.cc_inst.dlyd_1_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[185] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlyd_2 \cm_inst.cc_inst.dlyd_2_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[186] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dlyd_4 \cm_inst.cc_inst.dlyd_4_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .Z(\cm_inst.cc_inst.out_notouch_[187] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__hold \cm_inst.cc_inst.hold_inst  (.Z(\cm_inst.cc_inst.out_notouch_[173] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__icgtn_1 \cm_inst.cc_inst.icgtn_1_inst  (.CLKN(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .TE(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[204] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__icgtn_2 \cm_inst.cc_inst.icgtn_2_inst  (.CLKN(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .TE(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[205] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__icgtn_4 \cm_inst.cc_inst.icgtn_4_inst  (.CLKN(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .TE(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[206] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__icgtp_2 \cm_inst.cc_inst.icgtp_2_inst  (.CLK(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .TE(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[208] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__icgtp_4 \cm_inst.cc_inst.icgtp_4_inst  (.CLK(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .TE(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[209] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 \cm_inst.cc_inst.inv_12_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[15] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 \cm_inst.cc_inst.inv_16_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[16] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \cm_inst.cc_inst.inv_1_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[10] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 \cm_inst.cc_inst.inv_20_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[17] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 \cm_inst.cc_inst.inv_2_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[11] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 \cm_inst.cc_inst.inv_3_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[12] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 \cm_inst.cc_inst.inv_4_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[13] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 \cm_inst.cc_inst.inv_8_inst  (.I(\cm_inst.cc_inst.in[0] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[14] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__invz_12 \cm_inst.cc_inst.invz_12_inst  (.EN(\cm_inst.cc_inst.in[2] ),
    .I(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[175] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__invz_1 \cm_inst.cc_inst.invz_1_inst  (.EN(\cm_inst.cc_inst.in[2] ),
    .I(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[173] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__invz_2 \cm_inst.cc_inst.invz_2_inst  (.EN(\cm_inst.cc_inst.in[0] ),
    .I(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[174] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__invz_3 \cm_inst.cc_inst.invz_3_inst  (.EN(\cm_inst.cc_inst.in[2] ),
    .I(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[174] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__invz_4 \cm_inst.cc_inst.invz_4_inst  (.EN(\cm_inst.cc_inst.in[4] ),
    .I(\cm_inst.cc_inst.in[5] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[174] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__invz_8 \cm_inst.cc_inst.invz_8_inst  (.EN(\cm_inst.cc_inst.in[0] ),
    .I(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[175] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latq_1 \cm_inst.cc_inst.latq_1_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .Q(\cm_inst.cc_inst.out_notouch_[123] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latq_2 \cm_inst.cc_inst.latq_2_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .Q(\cm_inst.cc_inst.out_notouch_[124] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latq_4 \cm_inst.cc_inst.latq_4_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .Q(\cm_inst.cc_inst.out_notouch_[125] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latrnq_1 \cm_inst.cc_inst.latrnq_1_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[126] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latrnq_2 \cm_inst.cc_inst.latrnq_2_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[127] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latrnq_4 \cm_inst.cc_inst.latrnq_4_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[128] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 \cm_inst.cc_inst.latrsnq_1_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .Q(\cm_inst.cc_inst.out_notouch_[129] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latrsnq_2 \cm_inst.cc_inst.latrsnq_2_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .Q(\cm_inst.cc_inst.out_notouch_[130] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latrsnq_4 \cm_inst.cc_inst.latrsnq_4_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .Q(\cm_inst.cc_inst.out_notouch_[131] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latsnq_1 \cm_inst.cc_inst.latsnq_1_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .SETN(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[132] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latsnq_2 \cm_inst.cc_inst.latsnq_2_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .SETN(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[133] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latsnq_4 \cm_inst.cc_inst.latsnq_4_inst  (.D(\cm_inst.cc_inst.in[0] ),
    .E(\cm_inst.cc_inst.in[1] ),
    .SETN(\cm_inst.cc_inst.in[2] ),
    .Q(\cm_inst.cc_inst.out_notouch_[134] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 \cm_inst.cc_inst.mux2_1_inst  (.I0(\cm_inst.cc_inst.in[0] ),
    .I1(\cm_inst.cc_inst.in[1] ),
    .S(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[117] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 \cm_inst.cc_inst.mux2_2_inst  (.I0(\cm_inst.cc_inst.in[0] ),
    .I1(\cm_inst.cc_inst.in[1] ),
    .S(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[118] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 \cm_inst.cc_inst.mux2_4_inst  (.I0(\cm_inst.cc_inst.in[0] ),
    .I1(\cm_inst.cc_inst.in[1] ),
    .S(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[119] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_1 \cm_inst.cc_inst.mux4_1_inst  (.I0(\cm_inst.cc_inst.in[0] ),
    .I1(\cm_inst.cc_inst.in[1] ),
    .I2(\cm_inst.cc_inst.in[2] ),
    .I3(\cm_inst.cc_inst.in[3] ),
    .S0(\cm_inst.cc_inst.in[4] ),
    .S1(\cm_inst.cc_inst.in[5] ),
    .Z(\cm_inst.cc_inst.out_notouch_[120] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 \cm_inst.cc_inst.mux4_2_inst  (.I0(\cm_inst.cc_inst.in[0] ),
    .I1(\cm_inst.cc_inst.in[1] ),
    .I2(\cm_inst.cc_inst.in[2] ),
    .I3(\cm_inst.cc_inst.in[3] ),
    .S0(\cm_inst.cc_inst.in[4] ),
    .S1(\cm_inst.cc_inst.in[5] ),
    .Z(\cm_inst.cc_inst.out_notouch_[121] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 \cm_inst.cc_inst.mux4_4_inst  (.I0(\cm_inst.cc_inst.in[0] ),
    .I1(\cm_inst.cc_inst.in[1] ),
    .I2(\cm_inst.cc_inst.in[2] ),
    .I3(\cm_inst.cc_inst.in[3] ),
    .S0(\cm_inst.cc_inst.in[4] ),
    .S1(\cm_inst.cc_inst.in[5] ),
    .Z(\cm_inst.cc_inst.out_notouch_[122] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 \cm_inst.cc_inst.nand2_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[27] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 \cm_inst.cc_inst.nand2_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[28] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 \cm_inst.cc_inst.nand2_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[29] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 \cm_inst.cc_inst.nand3_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[30] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 \cm_inst.cc_inst.nand3_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[31] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 \cm_inst.cc_inst.nand3_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[32] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 \cm_inst.cc_inst.nand4_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[33] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 \cm_inst.cc_inst.nand4_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[34] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 \cm_inst.cc_inst.nand4_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[35] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 \cm_inst.cc_inst.nor2_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[36] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 \cm_inst.cc_inst.nor2_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[37] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 \cm_inst.cc_inst.nor2_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[38] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 \cm_inst.cc_inst.nor3_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[39] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 \cm_inst.cc_inst.nor3_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[40] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 \cm_inst.cc_inst.nor3_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[41] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor4_1 \cm_inst.cc_inst.nor4_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[42] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 \cm_inst.cc_inst.nor4_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[43] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 \cm_inst.cc_inst.nor4_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[44] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 \cm_inst.cc_inst.oai211_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .C(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[96] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 \cm_inst.cc_inst.oai211_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .C(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[97] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 \cm_inst.cc_inst.oai211_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .C(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[98] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 \cm_inst.cc_inst.oai21_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[81] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 \cm_inst.cc_inst.oai21_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[82] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 \cm_inst.cc_inst.oai21_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[83] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 \cm_inst.cc_inst.oai221_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C(\cm_inst.cc_inst.in[4] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[99] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 \cm_inst.cc_inst.oai221_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C(\cm_inst.cc_inst.in[4] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[100] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 \cm_inst.cc_inst.oai221_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C(\cm_inst.cc_inst.in[4] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[101] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai222_1 \cm_inst.cc_inst.oai222_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C1(\cm_inst.cc_inst.in[4] ),
    .C2(\cm_inst.cc_inst.in[5] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[102] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 \cm_inst.cc_inst.oai222_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C1(\cm_inst.cc_inst.in[4] ),
    .C2(\cm_inst.cc_inst.in[5] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[103] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai222_4 \cm_inst.cc_inst.oai222_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .C1(\cm_inst.cc_inst.in[4] ),
    .C2(\cm_inst.cc_inst.in[5] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[104] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 \cm_inst.cc_inst.oai22_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[84] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 \cm_inst.cc_inst.oai22_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[85] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 \cm_inst.cc_inst.oai22_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .B1(\cm_inst.cc_inst.in[2] ),
    .B2(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[86] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 \cm_inst.cc_inst.oai31_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .B(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[87] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 \cm_inst.cc_inst.oai31_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .B(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[88] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 \cm_inst.cc_inst.oai31_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .B(\cm_inst.cc_inst.in[3] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[89] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 \cm_inst.cc_inst.oai32_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .B1(\cm_inst.cc_inst.in[3] ),
    .B2(\cm_inst.cc_inst.in[4] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[90] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 \cm_inst.cc_inst.oai32_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .B1(\cm_inst.cc_inst.in[3] ),
    .B2(\cm_inst.cc_inst.in[4] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[91] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 \cm_inst.cc_inst.oai32_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .B1(\cm_inst.cc_inst.in[3] ),
    .B2(\cm_inst.cc_inst.in[4] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[92] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai33_1 \cm_inst.cc_inst.oai33_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .B1(\cm_inst.cc_inst.in[3] ),
    .B2(\cm_inst.cc_inst.in[4] ),
    .B3(\cm_inst.cc_inst.in[5] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[93] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 \cm_inst.cc_inst.oai33_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .B1(\cm_inst.cc_inst.in[3] ),
    .B2(\cm_inst.cc_inst.in[4] ),
    .B3(\cm_inst.cc_inst.in[5] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[94] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__oai33_4 \cm_inst.cc_inst.oai33_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .B1(\cm_inst.cc_inst.in[3] ),
    .B2(\cm_inst.cc_inst.in[4] ),
    .B3(\cm_inst.cc_inst.in[5] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[95] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 \cm_inst.cc_inst.or2_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[45] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 \cm_inst.cc_inst.or2_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[46] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 \cm_inst.cc_inst.or2_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[47] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__or3_1 \cm_inst.cc_inst.or3_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[48] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 \cm_inst.cc_inst.or3_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[49] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 \cm_inst.cc_inst.or3_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[50] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__or4_1 \cm_inst.cc_inst.or4_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .Z(\cm_inst.cc_inst.out_notouch_[51] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 \cm_inst.cc_inst.or4_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .Z(\cm_inst.cc_inst.out_notouch_[52] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 \cm_inst.cc_inst.or4_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .A4(\cm_inst.cc_inst.in[3] ),
    .Z(\cm_inst.cc_inst.out_notouch_[53] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffq_1 \cm_inst.cc_inst.sdffq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SE(\cm_inst.cc_inst.in[2] ),
    .SI(\cm_inst.cc_inst.in[3] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[159] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffq_2 \cm_inst.cc_inst.sdffq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SE(\cm_inst.cc_inst.in[2] ),
    .SI(\cm_inst.cc_inst.in[3] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[160] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffq_4 \cm_inst.cc_inst.sdffq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SE(\cm_inst.cc_inst.in[2] ),
    .SI(\cm_inst.cc_inst.in[3] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[161] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1 \cm_inst.cc_inst.sdffrnq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SE(\cm_inst.cc_inst.in[3] ),
    .SI(\cm_inst.cc_inst.in[4] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[162] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 \cm_inst.cc_inst.sdffrnq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SE(\cm_inst.cc_inst.in[3] ),
    .SI(\cm_inst.cc_inst.in[4] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[163] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4 \cm_inst.cc_inst.sdffrnq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SE(\cm_inst.cc_inst.in[3] ),
    .SI(\cm_inst.cc_inst.in[4] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[164] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1 \cm_inst.cc_inst.sdffrsnq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SE(\cm_inst.cc_inst.in[3] ),
    .SETN(\cm_inst.cc_inst.in[4] ),
    .SI(\cm_inst.cc_inst.in[5] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[165] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2 \cm_inst.cc_inst.sdffrsnq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SE(\cm_inst.cc_inst.in[3] ),
    .SETN(\cm_inst.cc_inst.in[4] ),
    .SI(\cm_inst.cc_inst.in[5] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[166] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4 \cm_inst.cc_inst.sdffrsnq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .RN(\cm_inst.cc_inst.in[2] ),
    .SE(\cm_inst.cc_inst.in[3] ),
    .SETN(\cm_inst.cc_inst.in[4] ),
    .SI(\cm_inst.cc_inst.in[5] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[167] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1 \cm_inst.cc_inst.sdffsnq_1_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SE(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .SI(\cm_inst.cc_inst.in[4] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[168] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2 \cm_inst.cc_inst.sdffsnq_2_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SE(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .SI(\cm_inst.cc_inst.in[4] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[169] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4 \cm_inst.cc_inst.sdffsnq_4_inst  (.D(\cm_inst.cc_inst.in[1] ),
    .SE(\cm_inst.cc_inst.in[2] ),
    .SETN(\cm_inst.cc_inst.in[3] ),
    .SI(\cm_inst.cc_inst.in[4] ),
    .CLK(\cm_inst.cc_inst.in[0] ),
    .Q(\cm_inst.cc_inst.out_notouch_[170] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tieh \cm_inst.cc_inst.tieh_inst  (.Z(\cm_inst.cc_inst.out_notouch_[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel \cm_inst.cc_inst.tiel_inst  (.ZN(\cm_inst.cc_inst.out_notouch_[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 \cm_inst.cc_inst.xnor2_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[54] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 \cm_inst.cc_inst.xnor2_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[55] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 \cm_inst.cc_inst.xnor2_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[56] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 \cm_inst.cc_inst.xnor3_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[57] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 \cm_inst.cc_inst.xnor3_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[58] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_4 \cm_inst.cc_inst.xnor3_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .ZN(\cm_inst.cc_inst.out_notouch_[59] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 \cm_inst.cc_inst.xor2_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[60] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 \cm_inst.cc_inst.xor2_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[61] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 \cm_inst.cc_inst.xor2_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .Z(\cm_inst.cc_inst.out_notouch_[62] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 \cm_inst.cc_inst.xor3_1_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[63] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 \cm_inst.cc_inst.xor3_2_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[64] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xor3_4 \cm_inst.cc_inst.xor3_4_inst  (.A1(\cm_inst.cc_inst.in[0] ),
    .A2(\cm_inst.cc_inst.in[1] ),
    .A3(\cm_inst.cc_inst.in[2] ),
    .Z(\cm_inst.cc_inst.out_notouch_[65] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__icgtp_2 \ro_inst.clock_gate  (.CLK(\ro_inst.ring[0] ),
    .E(\ro_inst.running ),
    .TE(_243_),
    .Q(\ro_inst.counter[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.clock_gate_inv  (.I(\ro_inst.counter[0] ),
    .ZN(\ro_inst.counter_n[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[10].div_flop  (.D(\ro_inst.counter_n[10] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[9] ),
    .Q(\ro_inst.counter[10] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[10].div_flop_inv  (.I(\ro_inst.counter[10] ),
    .ZN(\ro_inst.counter_n[10] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[11].div_flop  (.D(\ro_inst.counter_n[11] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[10] ),
    .Q(\ro_inst.counter[11] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[11].div_flop_inv  (.I(\ro_inst.counter[11] ),
    .ZN(\ro_inst.counter_n[11] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[12].div_flop  (.D(\ro_inst.counter_n[12] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[11] ),
    .Q(\ro_inst.counter[12] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[12].div_flop_inv  (.I(\ro_inst.counter[12] ),
    .ZN(\ro_inst.counter_n[12] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[13].div_flop  (.D(\ro_inst.counter_n[13] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[12] ),
    .Q(\ro_inst.counter[13] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[13].div_flop_inv  (.I(\ro_inst.counter[13] ),
    .ZN(\ro_inst.counter_n[13] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[14].div_flop  (.D(\ro_inst.counter_n[14] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[13] ),
    .Q(\ro_inst.counter[14] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[14].div_flop_inv  (.I(\ro_inst.counter[14] ),
    .ZN(\ro_inst.counter_n[14] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[15].div_flop  (.D(\ro_inst.counter_n[15] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[14] ),
    .Q(\ro_inst.counter[15] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[15].div_flop_inv  (.I(\ro_inst.counter[15] ),
    .ZN(\ro_inst.counter_n[15] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[16].div_flop  (.D(\ro_inst.counter_n[16] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[15] ),
    .Q(\ro_inst.counter[16] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[16].div_flop_inv  (.I(\ro_inst.counter[16] ),
    .ZN(\ro_inst.counter_n[16] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[17].div_flop  (.D(\ro_inst.counter_n[17] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[16] ),
    .Q(\ro_inst.counter[17] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[17].div_flop_inv  (.I(\ro_inst.counter[17] ),
    .ZN(\ro_inst.counter_n[17] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[18].div_flop  (.D(\ro_inst.counter_n[18] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[17] ),
    .Q(\ro_inst.counter[18] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[18].div_flop_inv  (.I(\ro_inst.counter[18] ),
    .ZN(\ro_inst.counter_n[18] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[19].div_flop  (.D(\ro_inst.counter_n[19] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[18] ),
    .Q(\ro_inst.counter[19] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[19].div_flop_inv  (.I(\ro_inst.counter[19] ),
    .ZN(\ro_inst.counter_n[19] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[1].div_flop  (.D(\ro_inst.counter_n[1] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[0] ),
    .Q(\ro_inst.counter[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[1].div_flop_inv  (.I(\ro_inst.counter[1] ),
    .ZN(\ro_inst.counter_n[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[20].div_flop  (.D(\ro_inst.counter_n[20] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[19] ),
    .Q(\ro_inst.counter[20] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[20].div_flop_inv  (.I(\ro_inst.counter[20] ),
    .ZN(\ro_inst.counter_n[20] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[21].div_flop  (.D(\ro_inst.counter_n[21] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[20] ),
    .Q(\ro_inst.counter[21] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[21].div_flop_inv  (.I(\ro_inst.counter[21] ),
    .ZN(\ro_inst.counter_n[21] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[22].div_flop  (.D(\ro_inst.counter_n[22] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[21] ),
    .Q(\ro_inst.counter[22] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[22].div_flop_inv  (.I(\ro_inst.counter[22] ),
    .ZN(\ro_inst.counter_n[22] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[23].div_flop  (.D(\ro_inst.counter_n[23] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[22] ),
    .Q(\ro_inst.counter[23] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[23].div_flop_inv  (.I(\ro_inst.counter[23] ),
    .ZN(\ro_inst.counter_n[23] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[24].div_flop  (.D(\ro_inst.counter_n[24] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[23] ),
    .Q(\ro_inst.counter[24] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[24].div_flop_inv  (.I(\ro_inst.counter[24] ),
    .ZN(\ro_inst.counter_n[24] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[25].div_flop  (.D(\ro_inst.counter_n[25] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[24] ),
    .Q(\ro_inst.counter[25] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[25].div_flop_inv  (.I(\ro_inst.counter[25] ),
    .ZN(\ro_inst.counter_n[25] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[26].div_flop  (.D(\ro_inst.counter_n[26] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[25] ),
    .Q(\ro_inst.counter[26] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[26].div_flop_inv  (.I(\ro_inst.counter[26] ),
    .ZN(\ro_inst.counter_n[26] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[27].div_flop  (.D(\ro_inst.counter_n[27] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[26] ),
    .Q(\ro_inst.counter[27] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[27].div_flop_inv  (.I(\ro_inst.counter[27] ),
    .ZN(\ro_inst.counter_n[27] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[28].div_flop  (.D(\ro_inst.counter_n[28] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[27] ),
    .Q(\ro_inst.counter[28] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[28].div_flop_inv  (.I(\ro_inst.counter[28] ),
    .ZN(\ro_inst.counter_n[28] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[29].div_flop  (.D(\ro_inst.counter_n[29] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[28] ),
    .Q(\ro_inst.counter[29] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[29].div_flop_inv  (.I(\ro_inst.counter[29] ),
    .ZN(\ro_inst.counter_n[29] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[2].div_flop  (.D(\ro_inst.counter_n[2] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[1] ),
    .Q(\ro_inst.counter[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[2].div_flop_inv  (.I(\ro_inst.counter[2] ),
    .ZN(\ro_inst.counter_n[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[30].div_flop  (.D(\ro_inst.counter_n[30] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[29] ),
    .Q(\ro_inst.counter[30] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[30].div_flop_inv  (.I(\ro_inst.counter[30] ),
    .ZN(\ro_inst.counter_n[30] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[31].div_flop  (.D(\ro_inst.counter_n[31] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[30] ),
    .Q(\ro_inst.counter[31] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[31].div_flop_inv  (.I(\ro_inst.counter[31] ),
    .ZN(\ro_inst.counter_n[31] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[32].div_flop  (.D(\ro_inst.counter_n[32] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[31] ),
    .Q(\ro_inst.counter[32] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[32].div_flop_inv  (.I(\ro_inst.counter[32] ),
    .ZN(\ro_inst.counter_n[32] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[33].div_flop  (.D(\ro_inst.counter_n[33] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[32] ),
    .Q(\ro_inst.counter[33] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[33].div_flop_inv  (.I(\ro_inst.counter[33] ),
    .ZN(\ro_inst.counter_n[33] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[34].div_flop  (.D(\ro_inst.counter_n[34] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[33] ),
    .Q(\ro_inst.counter[34] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[34].div_flop_inv  (.I(\ro_inst.counter[34] ),
    .ZN(\ro_inst.counter_n[34] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[3].div_flop  (.D(\ro_inst.counter_n[3] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[2] ),
    .Q(\ro_inst.counter[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[3].div_flop_inv  (.I(\ro_inst.counter[3] ),
    .ZN(\ro_inst.counter_n[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[4].div_flop  (.D(\ro_inst.counter_n[4] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[3] ),
    .Q(\ro_inst.counter[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[4].div_flop_inv  (.I(\ro_inst.counter[4] ),
    .ZN(\ro_inst.counter_n[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[5].div_flop  (.D(\ro_inst.counter_n[5] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[4] ),
    .Q(\ro_inst.counter[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[5].div_flop_inv  (.I(\ro_inst.counter[5] ),
    .ZN(\ro_inst.counter_n[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[6].div_flop  (.D(\ro_inst.counter_n[6] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[5] ),
    .Q(\ro_inst.counter[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[6].div_flop_inv  (.I(\ro_inst.counter[6] ),
    .ZN(\ro_inst.counter_n[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[7].div_flop  (.D(\ro_inst.counter_n[7] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[6] ),
    .Q(\ro_inst.counter[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[7].div_flop_inv  (.I(\ro_inst.counter[7] ),
    .ZN(\ro_inst.counter_n[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[8].div_flop  (.D(\ro_inst.counter_n[8] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[7] ),
    .Q(\ro_inst.counter[8] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[8].div_flop_inv  (.I(\ro_inst.counter[8] ),
    .ZN(\ro_inst.counter_n[8] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 \ro_inst.gcount[9].div_flop  (.D(\ro_inst.counter_n[9] ),
    .RN(in[0]),
    .CLK(\ro_inst.counter_n[8] ),
    .Q(\ro_inst.counter[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.gcount[9].div_flop_inv  (.I(\ro_inst.counter[9] ),
    .ZN(\ro_inst.counter_n[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 \ro_inst.ring_osc_0  (.A1(\ro_inst.ring[0] ),
    .A2(\ro_inst.enable ),
    .ZN(\ro_inst.ring[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.ring_osc_1  (.I(\ro_inst.ring[1] ),
    .ZN(\ro_inst.ring[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.ring_osc_2  (.I(\ro_inst.ring[2] ),
    .ZN(\ro_inst.ring[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 \ro_inst.sig_cmp  (.A1(\ro_inst.signal ),
    .A2(\ro_inst.saved_signal ),
    .ZN(\ro_inst.running ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__latq_1 \ro_inst.sig_latch  (.D(\ro_inst.signal ),
    .E(\ro_inst.slow_clk_n ),
    .Q(\ro_inst.saved_signal ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 \ro_inst.slow_clock_inv  (.I(in[0]),
    .ZN(\ro_inst.slow_clk_n ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
endmodule
