VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO loopback9
  CLASS BLOCK ;
  FOREIGN loopback9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.853500 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 196.000 74.480 200.000 ;
    END
  END clk
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.640 4.000 81.200 ;
    END
  END in[0]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.877500 ;
    ANTENNADIFFAREA 0.813600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 73.920 200.000 74.480 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.317000 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 127.680 200.000 128.240 ;
    END
  END in[11]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.877500 ;
    ANTENNADIFFAREA 0.813600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 84.000 200.000 84.560 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.317000 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 87.360 200.000 87.920 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.877500 ;
    ANTENNADIFFAREA 0.813600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 94.080 200.000 94.640 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.317000 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 80.640 200.000 81.200 ;
    END
  END in[15]
  PIN in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.877500 ;
    ANTENNADIFFAREA 0.813600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 97.440 200.000 98.000 ;
    END
  END in[16]
  PIN in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.317000 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 100.800 200.000 101.360 ;
    END
  END in[17]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 4.000 98.000 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.317000 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.877500 ;
    ANTENNADIFFAREA 0.813600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.317000 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END in[9]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 196.000 77.840 200.000 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 90.720 200.000 91.280 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 117.600 200.000 118.160 ;
    END
  END out[11]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.121000 ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 120.960 200.000 121.520 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 110.880 200.000 111.440 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.121000 ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 114.240 200.000 114.800 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 77.280 200.000 77.840 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.121000 ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 124.320 200.000 124.880 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 107.520 200.000 108.080 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.121000 ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 104.160 200.000 104.720 ;
    END
  END out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 29.230 19.860 30.830 181.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 75.850 19.860 77.450 181.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.470 19.860 124.070 181.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.090 19.860 170.690 181.740 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 52.540 19.860 54.140 181.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.160 19.860 100.760 181.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 145.780 19.860 147.380 181.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 192.400 19.860 194.000 181.740 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 19.710 194.000 181.890 ;
      LAYER Metal2 ;
        RECT 20.300 195.700 73.620 196.000 ;
        RECT 74.780 195.700 76.980 196.000 ;
        RECT 78.140 195.700 193.860 196.000 ;
        RECT 20.300 19.970 193.860 195.700 ;
      LAYER Metal3 ;
        RECT 4.000 128.540 196.000 181.580 ;
        RECT 4.000 127.380 195.700 128.540 ;
        RECT 4.000 125.180 196.000 127.380 ;
        RECT 4.000 124.020 195.700 125.180 ;
        RECT 4.000 121.820 196.000 124.020 ;
        RECT 4.300 120.660 195.700 121.820 ;
        RECT 4.000 118.460 196.000 120.660 ;
        RECT 4.300 117.300 195.700 118.460 ;
        RECT 4.000 115.100 196.000 117.300 ;
        RECT 4.300 113.940 195.700 115.100 ;
        RECT 4.000 111.740 196.000 113.940 ;
        RECT 4.300 110.580 195.700 111.740 ;
        RECT 4.000 108.380 196.000 110.580 ;
        RECT 4.300 107.220 195.700 108.380 ;
        RECT 4.000 105.020 196.000 107.220 ;
        RECT 4.300 103.860 195.700 105.020 ;
        RECT 4.000 101.660 196.000 103.860 ;
        RECT 4.300 100.500 195.700 101.660 ;
        RECT 4.000 98.300 196.000 100.500 ;
        RECT 4.300 97.140 195.700 98.300 ;
        RECT 4.000 94.940 196.000 97.140 ;
        RECT 4.300 93.780 195.700 94.940 ;
        RECT 4.000 91.580 196.000 93.780 ;
        RECT 4.300 90.420 195.700 91.580 ;
        RECT 4.000 88.220 196.000 90.420 ;
        RECT 4.300 87.060 195.700 88.220 ;
        RECT 4.000 84.860 196.000 87.060 ;
        RECT 4.300 83.700 195.700 84.860 ;
        RECT 4.000 81.500 196.000 83.700 ;
        RECT 4.300 80.340 195.700 81.500 ;
        RECT 4.000 78.140 196.000 80.340 ;
        RECT 4.000 76.980 195.700 78.140 ;
        RECT 4.000 74.780 196.000 76.980 ;
        RECT 4.000 73.620 195.700 74.780 ;
        RECT 4.000 20.020 196.000 73.620 ;
  END
END loopback9
END LIBRARY

