* NGSPICE file created from cells7.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2 D RN SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2 D SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_1 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_16 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_1 D SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2 D RN SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__addf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__addf_2 A B CI CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_4 D SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_2 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1 D RN SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__icgtp_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__icgtp_1 CLK E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__bufz_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_1 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_2 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4 D RN SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__icgtp_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__icgtp_4 CLK E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_2 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__bufz_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_4 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latsnq_1 D E SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__bufz_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_16 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_12 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2 D RN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_8 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latsnq_4 D E SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 D RN SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2 D RN SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1 D SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1 D RN SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4 D SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4 D RN SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4 D SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__addf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__addf_1 A B CI CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4 D RN SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_1 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__bufz_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_12 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__addh_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__addh_2 A B CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrsnq_2 D E RN SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__icgtn_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__icgtn_2 CLKN E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__addf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__addf_4 A B CI CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_4 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_1 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__bufz_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_3 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_20 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_2 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_4 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_4 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1 D RN SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4 D RN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4 D RN SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__hold abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__hold Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_16 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_2 D SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_12 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__addh_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__addh_1 A B CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrsnq_1 D E RN SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__icgtn_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__icgtn_1 CLKN E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_3 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2 D RN SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__icgtp_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__icgtp_2 CLK E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__bufz_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_2 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__addh_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__addh_4 A B CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrsnq_4 D E RN SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_20 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__icgtn_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__icgtn_4 CLKN E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latsnq_2 D E SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_2 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_4 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_12 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2 D SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__bufz_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_8 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

.subckt cells7 clk in[0] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[1]
+ in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] out[0] out[10] out[11] out[1] out[2]
+ out[3] out[4] out[5] out[6] out[7] out[8] out[9] rst_n vdd vss
XTAP_TAPCELL_ROW_52_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_432_ cm_inst.cc_inst.out_notouch_\[39\] cm_inst.cc_inst.out_notouch_\[47\] cm_inst.cc_inst.out_notouch_\[55\]
+ cm_inst.cc_inst.out_notouch_\[63\] _071_ _072_ _198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_501_ _007_ net297 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_363_ cm_inst.cc_inst.out_notouch_\[99\] cm_inst.cc_inst.out_notouch_\[107\] cm_inst.cc_inst.out_notouch_\[115\]
+ cm_inst.cc_inst.out_notouch_\[123\] _025_ _021_ _133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_294_ cm_inst.page\[3\] _066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout105 net108 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout127 net128 net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout138 net139 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout149 net150 net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout116 net118 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.dffrsnq_2_inst net191 net120 net62 net284 cm_inst.cc_inst.out_notouch_\[154\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2
XTAP_TAPCELL_ROW_5_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_346_ cm_inst.cc_inst.out_notouch_\[34\] cm_inst.cc_inst.out_notouch_\[42\] cm_inst.cc_inst.out_notouch_\[50\]
+ cm_inst.cc_inst.out_notouch_\[58\] _115_ _116_ _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_415_ cm_inst.cc_inst.out_notouch_\[102\] cm_inst.cc_inst.out_notouch_\[110\] cm_inst.cc_inst.out_notouch_\[118\]
+ cm_inst.cc_inst.out_notouch_\[126\] _105_ _106_ _182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_277_ _049_ _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_11_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout19_I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_4_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xro_inst.gcount\[20\].div_flop ro_inst.counter_n\[20\] net299 ro_inst.counter_n\[19\]
+ ro_inst.counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_fanout223_I net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_329_ _088_ _095_ _099_ _047_ _100_ _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_51_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__373__S _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xcm_inst.cc_inst.and3_2_inst net252 net168 net102 cm_inst.cc_inst.out_notouch_\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.sdffsnq_2_inst net179 net106 net62 net25 net283 cm_inst.cc_inst.out_notouch_\[169\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_50_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.mux2_1_inst net276 net185 net116 cm_inst.cc_inst.out_notouch_\[117\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_1
XFILLER_0_7_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.clkbuf_4_inst net256 cm_inst.cc_inst.out_notouch_\[191\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XPHY_EDGE_ROW_7_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xfanout309 net310 net309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.dlya_1_inst net229 cm_inst.cc_inst.out_notouch_\[176\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlya_1
Xcm_inst.cc_inst.xnor3_2_inst net262 net174 net105 cm_inst.cc_inst.out_notouch_\[58\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_500_ _006_ net296 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_431_ _197_ net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_362_ _130_ _131_ _074_ _132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_293_ _059_ _065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout106 net108 net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout117 net118 net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout139 net140 net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout128 cm_inst.cc_inst.in\[2\] net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_345_ _026_ _116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_276_ cm_inst.page\[0\] _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xro_inst.gcount\[10\].div_flop ro_inst.counter_n\[10\] net296 ro_inst.counter_n\[9\]
+ ro_inst.counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_414_ _181_ net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_11_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_259_ _031_ _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_328_ _059_ _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.clkinv_16_inst net220 cm_inst.cc_inst.out_notouch_\[202\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_16
XTAP_TAPCELL_ROW_47_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout31_I net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xcm_inst.cc_inst.dffsnq_2_inst net177 net107 net263 cm_inst.cc_inst.out_notouch_\[157\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_0_21_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.sdffq_1_inst net164 net100 net58 net248 cm_inst.cc_inst.out_notouch_\[159\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA_fanout79_I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.dffnrsnq_2_inst net184 net114 net61 net272 cm_inst.cc_inst.out_notouch_\[142\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2
XFILLER_0_21_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout283_I net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.oai32_1_inst net286 net194 net122 net65 net34 cm_inst.cc_inst.out_notouch_\[90\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput10 net10 out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.inv_2_inst net213 cm_inst.cc_inst.out_notouch_\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_1_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input3_I in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_430_ _196_ ro_inst.counter\[34\] _148_ _197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_361_ cm_inst.cc_inst.out_notouch_\[3\] cm_inst.cc_inst.out_notouch_\[11\] cm_inst.cc_inst.out_notouch_\[19\]
+ cm_inst.cc_inst.out_notouch_\[27\] _081_ _082_ _131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_292_ _064_ net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xro_inst.gcount\[7\].div_flop ro_inst.counter_n\[7\] net299 ro_inst.counter_n\[6\]
+ ro_inst.counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_23_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand3_1_inst_A2 net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout246_I net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout107 net108 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout129 net130 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout118 net126 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__281__I _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_413_ _180_ ro_inst.counter\[5\] _148_ _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_28_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_344_ _049_ _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__392__S _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_275_ _040_ _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.clock_gate_315 net315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xro_inst.gcount\[8\].div_flop_inv ro_inst.counter\[8\] ro_inst.counter_n\[8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_16_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_327_ _048_ _096_ _097_ _098_ _099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_258_ _030_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xcm_inst.cc_inst.mux4_2_inst net276 net159 net94 net48 net31 net19 cm_inst.cc_inst.out_notouch_\[121\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_24_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout24_I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xro_inst.gcount\[33\].div_flop_inv ro_inst.counter\[33\] ro_inst.counter_n\[33\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout290 net291 net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_36_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.aoi21_4_inst net227 net147 net86 cm_inst.cc_inst.out_notouch_\[68\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_46_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.dlyc_2_inst net257 cm_inst.cc_inst.out_notouch_\[183\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_0_21_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__374__I _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput9 net9 out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 net11 out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xcm_inst.cc_inst.oai222_2_inst net235 net154 net90 net46 net29 net18 cm_inst.cc_inst.out_notouch_\[103\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__279__I _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_360_ cm_inst.cc_inst.out_notouch_\[35\] cm_inst.cc_inst.out_notouch_\[43\] cm_inst.cc_inst.out_notouch_\[51\]
+ cm_inst.cc_inst.out_notouch_\[59\] _071_ _072_ _130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_291_ _062_ ro_inst.counter\[0\] _063_ _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xro_inst.gcount\[26\].div_flop_inv ro_inst.counter\[26\] ro_inst.counter_n\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_cm_inst.cc_inst.nand3_1_inst_A3 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_489_ _239_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout119 net120 net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout108 net109 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__336__S0 _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_412_ _065_ _174_ _179_ _102_ _180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_28_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_343_ _112_ _113_ _114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_274_ _046_ _047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_24_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.mux2_4_inst net234 net153 net89 cm_inst.cc_inst.out_notouch_\[119\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_4
XANTENNA_cm_inst.cc_inst.bufz_3_inst_I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_326_ _069_ _054_ cm_inst.cc_inst.out_notouch_\[209\] _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_16_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_257_ cm_inst.page\[2\] _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xfanout90 net91 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout17_I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xro_inst.gcount\[19\].div_flop_inv ro_inst.counter\[19\] ro_inst.counter_n\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout291 net292 net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout280 net291 net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_44_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_309_ _037_ _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_21_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.dlya_4_inst net240 cm_inst.cc_inst.out_notouch_\[178\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlya_4
Xcm_inst.cc_inst.or2_2_inst net253 net169 cm_inst.cc_inst.out_notouch_\[46\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_21_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_SETN net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__390__S1 _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.nor2_1_inst net260 net176 cm_inst.cc_inst.out_notouch_\[36\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__381__S1 _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.addf_2_inst net232 net152 net91 cm_inst.cc_inst.out_notouch_\[107\]
+ cm_inst.cc_inst.out_notouch_\[108\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__addf_2
Xoutput12 net12 out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xcm_inst.cc_inst.nand2_1_inst net212 net136 cm_inst.cc_inst.out_notouch_\[27\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_290_ ro_inst.enable _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_48_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_488_ net3 ro_sel\[0\] _238_ _239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout109 net110 net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_342_ cm_inst.cc_inst.out_notouch_\[2\] cm_inst.cc_inst.out_notouch_\[10\] cm_inst.cc_inst.out_notouch_\[18\]
+ cm_inst.cc_inst.out_notouch_\[26\] _089_ _027_ _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_411_ _088_ _177_ _178_ _125_ _100_ _179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_28_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_273_ _030_ cm_inst.page\[3\] _046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.sdffq_4_inst net192 net106 net56 net283 cm_inst.cc_inst.out_notouch_\[161\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffq_4
XFILLER_0_10_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcm_inst.cc_inst.aoi222_2_inst net237 net156 net92 net47 net30 net19 cm_inst.cc_inst.out_notouch_\[79\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_325_ _055_ cm_inst.cc_inst.out_notouch_\[201\] _097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout91 net97 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout80 net81 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_24_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_256_ cm_inst.cc_inst.out_notouch_\[0\] cm_inst.cc_inst.out_notouch_\[8\] cm_inst.cc_inst.out_notouch_\[16\]
+ cm_inst.cc_inst.out_notouch_\[24\] _025_ _021_ _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_19_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.oai32_4_inst net226 net147 net83 net43 net27 cm_inst.cc_inst.out_notouch_\[92\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_51_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout281 net282 net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout292 net293 net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcm_inst.cc_inst.oai21_1_inst net212 net138 net77 cm_inst.cc_inst.out_notouch_\[81\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout270 net274 net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_44_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_308_ _079_ _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xro_inst.gcount\[4\].div_flop_inv ro_inst.counter\[4\] ro_inst.counter_n\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.invz_2_inst net285 net195 cm_inst.cc_inst.out_notouch_\[174\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_12_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.sdffrsnq_1_inst net190 net119 net57 net35 net17 net281 cm_inst.cc_inst.out_notouch_\[165\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1
XPHY_EDGE_ROW_11_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput13 net13 out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.icgtp_1_inst net249 net166 net101 cm_inst.cc_inst.out_notouch_\[207\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XFILLER_0_7_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_487_ net6 net7 net8 net2 _238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xcm_inst.cc_inst.bufz_1_inst net256 net173 cm_inst.cc_inst.out_notouch_\[171\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__bufz_1
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_410_ cm_inst.cc_inst.out_notouch_\[197\] cm_inst.cc_inst.out_notouch_\[205\] _144_
+ _178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_272_ _041_ _043_ _044_ _045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_341_ _031_ _112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_28_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.and2_1_inst net250 net167 cm_inst.cc_inst.out_notouch_\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xro_inst.gcount\[22\].div_flop_inv ro_inst.counter\[22\] ro_inst.counter_n\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xro_inst.gcount\[6\].div_flop ro_inst.counter_n\[6\] net299 ro_inst.counter_n\[5\]
+ ro_inst.counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_18_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_255_ cm_inst.cc_inst.out_notouch_\[32\] cm_inst.cc_inst.out_notouch_\[40\] cm_inst.cc_inst.out_notouch_\[48\]
+ cm_inst.cc_inst.out_notouch_\[56\] _025_ _027_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_324_ _052_ cm_inst.cc_inst.out_notouch_\[193\] _096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout92 net96 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout81 net99 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout70 cm_inst.cc_inst.in\[3\] net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_38_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_41_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout282 net284 net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout260 net261 net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout271 net272 net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xcm_inst.cc_inst.nor4_2_inst net207 net135 net74 net38 cm_inst.cc_inst.out_notouch_\[43\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xfanout293 cm_inst.cc_inst.in\[0\] net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_44_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_307_ cm_inst.page\[2\] _079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.nand4_2_inst net260 net176 net106 net55 cm_inst.cc_inst.out_notouch_\[34\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_46_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout22_I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.oai211_2_inst net276 net186 net95 net59 cm_inst.cc_inst.out_notouch_\[97\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xcm_inst.cc_inst.xnor2_1_inst net253 net169 cm_inst.cc_inst.out_notouch_\[54\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_41_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xro_inst.gcount\[15\].div_flop_inv ro_inst.counter\[15\] ro_inst.counter_n\[15\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput14 net14 out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_34_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_486_ _237_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_271_ _031_ _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_340_ _107_ _110_ _044_ _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_469_ _218_ _228_ _065_ _221_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcm_inst.cc_inst.aoi22_1_inst net232 net151 net79 net40 cm_inst.cc_inst.out_notouch_\[69\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_323_ _091_ _093_ _094_ _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout60 net61 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_254_ _026_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout71 net72 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout82 net83 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout93 net96 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout187_I net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.nor2_4_inst net252 net168 cm_inst.cc_inst.out_notouch_\[38\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout261 net262 net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout283 net290 net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout272 net274 net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout250 net252 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xcm_inst.cc_inst.nand2_4_inst net210 net134 cm_inst.cc_inst.out_notouch_\[29\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xfanout294 net295 net294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_44_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_306_ _076_ _077_ _078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.clkinv_2_inst net254 cm_inst.cc_inst.out_notouch_\[197\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput15 net15 out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xro_inst.gcount\[29\].div_flop ro_inst.counter_n\[29\] net309 ro_inst.counter_n\[28\]
+ ro_inst.counter\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_43_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout267_I net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.buf_3_inst net271 cm_inst.cc_inst.out_notouch_\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_3
Xcm_inst.cc_inst.and4_2_inst net204 net132 net72 net39 cm_inst.cc_inst.out_notouch_\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_485_ _228_ _063_ _222_ _237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xcm_inst.cc_inst.aoi211_2_inst net213 net138 net77 net38 cm_inst.cc_inst.out_notouch_\[73\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__497__CLK net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.latq_2_inst net232 net151 cm_inst.cc_inst.out_notouch_\[124\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_48_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_270_ cm_inst.cc_inst.out_notouch_\[128\] cm_inst.cc_inst.out_notouch_\[136\] cm_inst.cc_inst.out_notouch_\[144\]
+ cm_inst.cc_inst.out_notouch_\[152\] _038_ _042_ _043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__420__S0 _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xcm_inst.cc_inst.oai21_4_inst net227 net146 net82 cm_inst.cc_inst.out_notouch_\[83\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_19_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.oai33_1_inst_B1 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_468_ _226_ _228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_27_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.inv_8_inst net271 cm_inst.cc_inst.out_notouch_\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_8
X_399_ cm_inst.cc_inst.out_notouch_\[5\] cm_inst.cc_inst.out_notouch_\[13\] cm_inst.cc_inst.out_notouch_\[21\]
+ cm_inst.cc_inst.out_notouch_\[29\] _071_ _072_ _167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_10_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SETN net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_322_ _030_ _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xcm_inst.cc_inst.dlyb_1_inst net257 cm_inst.cc_inst.out_notouch_\[179\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_253_ cm_inst.page\[1\] _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout83 net84 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout72 net78 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout50 net51 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout61 net68 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout94 net96 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.sdffrsnq_4_inst net173 net104 net54 net25 net23 net256 cm_inst.cc_inst.out_notouch_\[167\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4
XTAP_TAPCELL_ROW_38_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout240 net242 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout284 net290 net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout262 net265 net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout251 net252 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout273 net274 net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout295 net298 net295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.oai221_1_inst net235 net154 net89 net46 net28 cm_inst.cc_inst.out_notouch_\[99\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_305_ cm_inst.cc_inst.out_notouch_\[97\] cm_inst.cc_inst.out_notouch_\[105\] cm_inst.cc_inst.out_notouch_\[113\]
+ cm_inst.cc_inst.out_notouch_\[121\] _019_ _023_ _077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_12_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.icgtp_4_inst net218 net141 net80 cm_inst.cc_inst.out_notouch_\[209\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__icgtp_4
XFILLER_0_11_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.latrnq_2_inst net234 net153 net89 cm_inst.cc_inst.out_notouch_\[127\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latrnq_2
Xro_inst.gcount\[19\].div_flop ro_inst.counter_n\[19\] net295 ro_inst.counter_n\[18\]
+ ro_inst.counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_16_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.bufz_4_inst net239 net157 cm_inst.cc_inst.out_notouch_\[172\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__bufz_4
XFILLER_0_25_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput16 net16 out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.and2_4_inst net250 net167 cm_inst.cc_inst.out_notouch_\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_4_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xro_inst.gcount\[11\].div_flop_inv ro_inst.counter\[11\] ro_inst.counter_n\[11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_15_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcm_inst.cc_inst.latsnq_1_inst net228 net145 net85 cm_inst.cc_inst.out_notouch_\[132\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latsnq_1
XTAP_TAPCELL_ROW_8_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_484_ _219_ _227_ _236_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.bufz_16_inst net281 net190 cm_inst.cc_inst.out_notouch_\[173\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__bufz_16
XFILLER_0_13_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.oai33_1_inst net221 net142 net79 net41 net24 net17 cm_inst.cc_inst.out_notouch_\[93\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_0_48_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai33_1_inst_B2 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.dffq_2_inst net144 net224 cm_inst.cc_inst.out_notouch_\[148\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_398_ cm_inst.cc_inst.out_notouch_\[37\] cm_inst.cc_inst.out_notouch_\[45\] cm_inst.cc_inst.out_notouch_\[53\]
+ cm_inst.cc_inst.out_notouch_\[61\] _051_ _069_ _166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_467_ _217_ _227_ _036_ _221_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_27_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_18_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.xnor2_4_inst net269 net183 cm_inst.cc_inst.out_notouch_\[56\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
X_321_ cm_inst.cc_inst.out_notouch_\[129\] cm_inst.cc_inst.out_notouch_\[137\] cm_inst.cc_inst.out_notouch_\[145\]
+ cm_inst.cc_inst.out_notouch_\[153\] _092_ _090_ _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xfanout62 net67 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout73 net75 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout51 net52 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout40 net41 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_252_ _018_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout84 net85 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout95 net96 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.buf_20_inst net204 cm_inst.cc_inst.out_notouch_\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_0_27_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout263 net265 net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout252 net254 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout274 net280 net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_3_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xfanout230 net231 net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout241 net243 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout285 net288 net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout296 net298 net296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_304_ _030_ _076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xro_inst.gcount\[5\].div_flop ro_inst.counter_n\[5\] net300 ro_inst.counter_n\[4\]
+ ro_inst.counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_20_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_45_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_C net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcells7_316 out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout68_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xcm_inst.cc_inst.aoi221_1_inst net226 net146 net82 net42 net26 cm_inst.cc_inst.out_notouch_\[75\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_8_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.aoi22_4_inst net238 net156 net92 net45 cm_inst.cc_inst.out_notouch_\[71\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XPHY_EDGE_ROW_32_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_483_ _230_ net17 _236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.dlyd_2_inst net238 cm_inst.cc_inst.out_notouch_\[186\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlyd_2
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai33_1_inst_B3 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_466_ _226_ _227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_397_ _165_ net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_27_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout63 net67 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_320_ _049_ _092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_36_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_251_ cm_inst.cc_inst.out_notouch_\[64\] cm_inst.cc_inst.out_notouch_\[72\] cm_inst.cc_inst.out_notouch_\[80\]
+ cm_inst.cc_inst.out_notouch_\[88\] _019_ _023_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xfanout74 net75 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout85 net88 net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout30 net32 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout96 net97 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout41 net52 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout52 net70 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_449_ _062_ _103_ _128_ _147_ ro_sel\[0\] ro_sel\[1\] _214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_50_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout264 net265 net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout286 net288 net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout253 net254 net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout275 net279 net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout231 net245 net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout297 net298 net297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout220 net221 net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout242 net243 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_303_ _070_ _073_ _074_ _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_B2 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout98_I net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcells7_317 out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_29_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.clkinv_12_inst net218 cm_inst.cc_inst.out_notouch_\[201\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_12
Xcm_inst.cc_inst.dffnrnq_2_inst net172 net103 net258 cm_inst.cc_inst.out_notouch_\[139\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_482_ _218_ _227_ _235_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xcm_inst.cc_inst.dlyb_4_inst net281 cm_inst.cc_inst.out_notouch_\[181\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xcm_inst.cc_inst.invz_8_inst net259 net173 cm_inst.cc_inst.out_notouch_\[175\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_8
XFILLER_0_45_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.or3_2_inst net201 net131 net71 cm_inst.cc_inst.out_notouch_\[49\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout80_I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xro_inst.gcount\[28\].div_flop ro_inst.counter_n\[28\] net309 ro_inst.counter_n\[27\]
+ ro_inst.counter\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_36_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xcm_inst.cc_inst.oai221_4_inst net277 net186 net116 net60 net33 cm_inst.cc_inst.out_notouch_\[101\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
Xcm_inst.cc_inst.nor3_1_inst net207 net135 net74 cm_inst.cc_inst.out_notouch_\[39\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_465_ net2 _226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_19_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.dffnsnq_1_inst net144 net86 net225 cm_inst.cc_inst.out_notouch_\[144\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
X_396_ _164_ ro_inst.counter\[4\] _148_ _165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcm_inst.cc_inst.nand3_1_inst net272 net189 net102 cm_inst.cc_inst.out_notouch_\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.gcount\[29\].div_flop_inv ro_inst.counter\[29\] ro_inst.counter_n\[29\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_1_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout53 net57 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout64 net66 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_250_ _020_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout20 net21 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout75 net76 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout86 net88 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout42 net43 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout31 net32 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_24_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout97 net98 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_448_ _213_ net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_379_ _147_ ro_inst.counter\[3\] _148_ _149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout265 net266 net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout287 net289 net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout254 net255 net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout210 net211 net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout298 net302 net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout232 net233 net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout243 net244 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout221 net222 net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout276 net279 net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_302_ _031_ _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.latsnq_4_inst net278 net187 net114 cm_inst.cc_inst.out_notouch_\[134\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latsnq_4
Xcells7_318 out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__428__A2 _193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xcm_inst.cc_inst.oai33_4_inst net238 net156 net92 net45 net27 net18 cm_inst.cc_inst.out_notouch_\[95\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_4
XFILLER_0_7_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.oai22_1_inst net226 net147 net84 net42 cm_inst.cc_inst.out_notouch_\[84\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xro_inst.gcount\[18\].div_flop ro_inst.counter_n\[18\] net295 ro_inst.counter_n\[17\]
+ ro_inst.counter\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_31_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai22_2_inst_B2 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_481_ _230_ net24 _235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__350__S0 _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_464_ _076_ _222_ _225_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_27_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_395_ _016_ _158_ _163_ _164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_50_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.dffrsnq_1_inst net178 net107 net56 net264 cm_inst.cc_inst.out_notouch_\[153\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XFILLER_0_10_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout21 net22 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_1_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout54 net57 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout65 net66 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout43 net44 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout32 net36 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout76 net77 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout87 net88 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout98 net99 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.sdffrnq_2_inst net173 net104 net54 net25 net256 cm_inst.cc_inst.out_notouch_\[163\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2
XFILLER_0_35_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_378_ ro_inst.enable _148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_27_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_447_ _212_ ro_inst.saved_signal ro_inst.enable _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout36_I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout200 cm_inst.cc_inst.in\[1\] net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout211 net215 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout222 net223 net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__252__I _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout288 net289 net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout266 net267 net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout255 net267 net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout277 net278 net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout233 net236 net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout244 net245 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout299 net301 net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_301_ cm_inst.cc_inst.out_notouch_\[1\] cm_inst.cc_inst.out_notouch_\[9\] cm_inst.cc_inst.out_notouch_\[17\]
+ cm_inst.cc_inst.out_notouch_\[25\] _071_ _072_ _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__337__I _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.and3_1_inst net201 net132 net72 cm_inst.cc_inst.out_notouch_\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_46_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__247__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.aoi221_4_inst net232 net151 net79 net40 net24 cm_inst.cc_inst.out_notouch_\[77\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xcells7_319 out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_40_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.sdffsnq_1_inst net150 net87 net44 net30 net229 cm_inst.cc_inst.out_notouch_\[168\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1
Xcm_inst.cc_inst.clkbuf_3_inst net278 cm_inst.cc_inst.out_notouch_\[190\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_43_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.gcount\[4\].div_flop ro_inst.counter_n\[4\] net305 ro_inst.counter_n\[3\]
+ ro_inst.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_47_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xro_inst.gcount\[7\].div_flop_inv ro_inst.counter\[7\] ro_inst.counter_n\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_480_ _217_ _227_ _234_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xcm_inst.cc_inst.clkinv_8_inst net219 cm_inst.cc_inst.out_notouch_\[200\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_8
Xro_inst.gcount\[32\].div_flop_inv ro_inst.counter\[32\] ro_inst.counter_n\[32\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xcm_inst.cc_inst.xnor3_1_inst net203 net131 net71 cm_inst.cc_inst.out_notouch_\[57\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_13_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_36_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.dffrnq_2_inst net164 net100 net247 cm_inst.cc_inst.out_notouch_\[151\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_463_ net5 _222_ _225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_394_ _036_ _161_ _162_ _125_ _060_ _163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout55 net56 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout33 net35 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout44 net51 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout22 net23 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_24_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout66 net67 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_32_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout77 net78 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout88 net98 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout99 net128 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_446_ _060_ _206_ _211_ cm_inst.page\[5\] _212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_377_ _065_ _140_ _146_ _102_ _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_23_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout116_I net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout29_I net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout256 net257 net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout201 net202 net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xcm_inst.cc_inst.tiel_inst cm_inst.cc_inst.out_notouch_\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xfanout212 net214 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout223 net246 net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout245 net246 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout234 net236 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout289 net290 net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout278 net279 net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout267 net292 net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_300_ _039_ _072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xro_inst.gcount\[25\].div_flop_inv ro_inst.counter\[25\] ro_inst.counter_n\[25\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.dffsnq_1_inst net144 net85 net225 cm_inst.cc_inst.out_notouch_\[156\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_EDGE_ROW_39_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_43_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_429_ _102_ _190_ _195_ _196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_23_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput1 in[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.dffnrsnq_1_inst net177 net107 net56 net263 cm_inst.cc_inst.out_notouch_\[141\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1
XFILLER_0_7_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.nor3_4_inst net201 net129 net71 cm_inst.cc_inst.out_notouch_\[41\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xcm_inst.cc_inst.dffnsnq_4_inst net191 net119 net282 cm_inst.cc_inst.out_notouch_\[146\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4
XFILLER_0_40_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.nand3_4_inst net273 net182 net111 cm_inst.cc_inst.out_notouch_\[32\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xcm_inst.cc_inst.inv_1_inst net250 cm_inst.cc_inst.out_notouch_\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_10_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xro_inst.gcount\[18\].div_flop_inv ro_inst.counter\[18\] ro_inst.counter_n\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout313_I net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout59_I net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__271__I _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.xor2_2_inst net201 net129 cm_inst.cc_inst.out_notouch_\[61\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_39_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_462_ _224_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_393_ cm_inst.cc_inst.out_notouch_\[196\] cm_inst.cc_inst.out_notouch_\[204\] _052_
+ _162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout56 net57 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout67 net68 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout34 net35 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout78 net81 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__266__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout23 cm_inst.cc_inst.in\[5\] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout89 net97 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout45 net50 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_32_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_445_ _033_ _209_ _210_ _124_ _059_ _211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_376_ _088_ _143_ _145_ _124_ _100_ _146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_23_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xro_inst.gcount\[27\].div_flop ro_inst.counter_n\[27\] net308 ro_inst.counter_n\[26\]
+ ro_inst.counter\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.mux4_1_inst net241 net158 net89 net46 net28 net18 cm_inst.cc_inst.out_notouch_\[120\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xfanout257 net259 net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout279 net280 net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout268 net270 net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout224 net225 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout202 net203 net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout213 net214 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout246 net293 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout235 net236 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_428_ _088_ _193_ _194_ _125_ _100_ _195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_15_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_359_ _129_ net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcm_inst.cc_inst.oai22_4_inst net283 net192 net120 net62 cm_inst.cc_inst.out_notouch_\[86\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
Xinput2 in[1] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_fanout41_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.dlyc_1_inst net287 cm_inst.cc_inst.out_notouch_\[182\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_11_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.dffrsnq_4_inst net172 net103 net53 net258 cm_inst.cc_inst.out_notouch_\[155\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcm_inst.cc_inst.oai222_1_inst net275 net185 net116 net59 net33 net20 cm_inst.cc_inst.out_notouch_\[102\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA_cm_inst.cc_inst.bufz_3_inst_EN net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xro_inst.gcount\[3\].div_flop_inv ro_inst.counter\[3\] ro_inst.counter_n\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.and3_2_inst_A3 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_461_ net4 _048_ _220_ _224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_392_ _159_ _160_ _044_ _161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_10_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xro_inst.gcount\[17\].div_flop ro_inst.counter_n\[17\] net294 ro_inst.counter_n\[16\]
+ ro_inst.counter\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_14_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.and3_4_inst net207 net135 net76 cm_inst.cc_inst.out_notouch_\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout57 net58 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout35 net36 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_32_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout79 net80 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout24 net37 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout46 net50 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_24_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout68 net69 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_444_ cm_inst.cc_inst.out_notouch_\[199\] cm_inst.cc_inst.out_notouch_\[207\] _144_
+ _210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcm_inst.cc_inst.sdffsnq_4_inst net157 net92 net48 net31 net239 cm_inst.cc_inst.out_notouch_\[170\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4
XFILLER_0_35_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_375_ cm_inst.cc_inst.out_notouch_\[195\] cm_inst.cc_inst.out_notouch_\[203\] _144_
+ _145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout258 net266 net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout247 net248 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout269 net270 net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout225 net228 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout214 net215 net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout203 net204 net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout236 net244 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_427_ cm_inst.cc_inst.out_notouch_\[198\] cm_inst.cc_inst.out_notouch_\[206\] _144_
+ _194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_358_ _128_ ro_inst.counter\[2\] _063_ _129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_289_ _016_ _035_ _061_ _062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout34_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 in[2] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_40_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.xnor3_4_inst net205 net133 net73 cm_inst.cc_inst.out_notouch_\[59\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_4
Xro_inst.gcount\[21\].div_flop_inv ro_inst.counter\[21\] ro_inst.counter_n\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcm_inst.cc_inst.or2_1_inst net202 net130 cm_inst.cc_inst.out_notouch_\[45\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_11_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.addf_1_inst net240 net159 net94 cm_inst.cc_inst.out_notouch_\[105\]
+ cm_inst.cc_inst.out_notouch_\[106\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__addf_1
XFILLER_0_3_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.buf_16_inst net268 cm_inst.cc_inst.out_notouch_\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_0_38_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xro_inst.gcount\[3\].div_flop ro_inst.counter_n\[3\] net305 ro_inst.counter_n\[2\]
+ ro_inst.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_0_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_391_ cm_inst.cc_inst.out_notouch_\[132\] cm_inst.cc_inst.out_notouch_\[140\] cm_inst.cc_inst.out_notouch_\[148\]
+ cm_inst.cc_inst.out_notouch_\[156\] _135_ _042_ _160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_460_ _055_ _221_ _223_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_50_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.dffsnq_4_inst net184 net113 net273 cm_inst.cc_inst.out_notouch_\[158\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XANTENNA_cm_inst.cc_inst.icgtp_4_inst_TE net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xro_inst.gcount\[14\].div_flop_inv ro_inst.counter\[14\] ro_inst.counter_n\[14\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_18_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout25 net37 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout69 net70 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout58 net69 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout36 net37 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout47 net48 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_443_ _207_ _208_ _094_ _209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_374_ _051_ _144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xcm_inst.cc_inst.aoi222_1_inst net287 net193 net121 net64 net33 net20 cm_inst.cc_inst.out_notouch_\[78\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA_fanout199_I net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xcm_inst.cc_inst.dffnrsnq_4_inst net164 net101 net58 net247 cm_inst.cc_inst.out_notouch_\[143\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4
XFILLER_0_25_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout204 net217 net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_14_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout259 net266 net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout248 net249 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout226 net227 net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout215 net216 net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout237 net239 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_426_ _191_ _192_ _032_ _193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_357_ _016_ _120_ _127_ _128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_11_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_288_ _036_ _045_ _047_ _058_ _060_ _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xinput4 in[3] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_34_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_cm_inst.cc_inst.and4_1_inst_A4 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.inv_4_inst net211 cm_inst.cc_inst.out_notouch_\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_4
XTAP_TAPCELL_ROW_40_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_409_ _175_ _176_ _094_ _177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.invz_1_inst net119 net63 cm_inst.cc_inst.out_notouch_\[173\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_0_6_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout181_I net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.mux4_4_inst net240 net159 net94 net48 net31 net19 cm_inst.cc_inst.out_notouch_\[122\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__479__A2 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_390_ cm_inst.cc_inst.out_notouch_\[164\] cm_inst.cc_inst.out_notouch_\[172\] cm_inst.cc_inst.out_notouch_\[180\]
+ cm_inst.cc_inst.out_notouch_\[188\] _038_ _040_ _159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_10_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout26 net28 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout37 cm_inst.cc_inst.in\[4\] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout48 net50 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout59 net61 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_373_ _141_ _142_ _094_ _143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_442_ cm_inst.cc_inst.out_notouch_\[135\] cm_inst.cc_inst.out_notouch_\[143\] cm_inst.cc_inst.out_notouch_\[151\]
+ cm_inst.cc_inst.out_notouch_\[159\] _050_ _068_ _208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.dlyc_4_inst net229 cm_inst.cc_inst.out_notouch_\[184\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlyc_4
XFILLER_0_14_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout227 net228 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout205 net206 net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout216 net217 net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout238 net239 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout249 net255 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_17_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.or4_2_inst net262 net174 net105 net55 cm_inst.cc_inst.out_notouch_\[52\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_32_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.bufz_12_inst net30 net19 cm_inst.cc_inst.out_notouch_\[172\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__bufz_12
X_425_ cm_inst.cc_inst.out_notouch_\[134\] cm_inst.cc_inst.out_notouch_\[142\] cm_inst.cc_inst.out_notouch_\[150\]
+ cm_inst.cc_inst.out_notouch_\[158\] _108_ _023_ _192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_287_ _059_ _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_356_ _036_ _123_ _125_ _126_ _060_ _127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xcm_inst.cc_inst.nor4_1_inst net260 net174 net105 net55 cm_inst.cc_inst.out_notouch_\[42\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_36_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 in[4] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xcm_inst.cc_inst.oai222_4_inst net241 net158 net90 net46 net29 net18 cm_inst.cc_inst.out_notouch_\[104\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
Xcm_inst.cc_inst.addh_2_inst net241 net158 cm_inst.cc_inst.out_notouch_\[113\] cm_inst.cc_inst.out_notouch_\[114\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__addh_2
XTAP_TAPCELL_ROW_34_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.nand4_1_inst net210 net129 net72 net39 cm_inst.cc_inst.out_notouch_\[33\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_52_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xro_inst.gcount\[26\].div_flop ro_inst.counter_n\[26\] net308 ro_inst.counter_n\[25\]
+ ro_inst.counter\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_2_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.oai211_1_inst net241 net158 net94 net49 cm_inst.cc_inst.out_notouch_\[96\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_408_ cm_inst.cc_inst.out_notouch_\[133\] cm_inst.cc_inst.out_notouch_\[141\] cm_inst.cc_inst.out_notouch_\[149\]
+ cm_inst.cc_inst.out_notouch_\[157\] _092_ _090_ _176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_339_ cm_inst.cc_inst.out_notouch_\[66\] cm_inst.cc_inst.out_notouch_\[74\] cm_inst.cc_inst.out_notouch_\[82\]
+ cm_inst.cc_inst.out_notouch_\[90\] _108_ _109_ _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XPHY_EDGE_ROW_44_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__299__I _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.latrsnq_2_inst net289 net196 net124 net66 cm_inst.cc_inst.out_notouch_\[130\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latrsnq_2
XFILLER_0_33_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.icgtn_2_inst net248 net164 net100 cm_inst.cc_inst.out_notouch_\[205\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__icgtn_2
XFILLER_0_12_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout291_I net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout304_I net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout38 net39 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout27 net28 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout49 net50 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_441_ cm_inst.cc_inst.out_notouch_\[167\] cm_inst.cc_inst.out_notouch_\[175\] cm_inst.cc_inst.out_notouch_\[183\]
+ cm_inst.cc_inst.out_notouch_\[191\] _115_ _116_ _207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_372_ cm_inst.cc_inst.out_notouch_\[131\] cm_inst.cc_inst.out_notouch_\[139\] cm_inst.cc_inst.out_notouch_\[147\]
+ cm_inst.cc_inst.out_notouch_\[155\] _115_ _068_ _142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xro_inst.gcount\[10\].div_flop_inv ro_inst.counter\[10\] ro_inst.counter_n\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout228 net231 net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout206 net209 net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcm_inst.cc_inst.or2_4_inst net206 net134 cm_inst.cc_inst.out_notouch_\[47\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
Xfanout217 net223 net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout239 net243 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xro_inst.gcount\[16\].div_flop ro_inst.counter_n\[16\] net294 ro_inst.counter_n\[15\]
+ ro_inst.counter\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_424_ cm_inst.cc_inst.out_notouch_\[166\] cm_inst.cc_inst.out_notouch_\[174\] cm_inst.cc_inst.out_notouch_\[182\]
+ cm_inst.cc_inst.out_notouch_\[190\] _105_ _109_ _191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xcm_inst.cc_inst.addf_4_inst net275 net185 net116 cm_inst.cc_inst.out_notouch_\[109\]
+ cm_inst.cc_inst.out_notouch_\[110\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__addf_4
X_355_ cm_inst.cc_inst.out_notouch_\[194\] cm_inst.cc_inst.out_notouch_\[202\] _052_
+ _126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_286_ cm_inst.page\[4\] _059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 in[5] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_34_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_407_ cm_inst.cc_inst.out_notouch_\[165\] cm_inst.cc_inst.out_notouch_\[173\] cm_inst.cc_inst.out_notouch_\[181\]
+ cm_inst.cc_inst.out_notouch_\[189\] _092_ _090_ _175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_338_ _020_ _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_269_ _039_ _042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.clkinv_1_inst net221 cm_inst.cc_inst.out_notouch_\[196\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout32_I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.buf_2_inst net213 cm_inst.cc_inst.out_notouch_\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_2
Xcm_inst.cc_inst.and4_1_inst net268 net182 net111 net61 cm_inst.cc_inst.out_notouch_\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcm_inst.cc_inst.aoi222_4_inst net277 net187 net114 net59 net33 net20 cm_inst.cc_inst.out_notouch_\[80\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout284_I net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.aoi211_1_inst net276 net186 net114 net59 cm_inst.cc_inst.out_notouch_\[72\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_4_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__496__CLK net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.latq_1_inst net234 net153 cm_inst.cc_inst.out_notouch_\[123\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_38_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout28 net32 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout39 net41 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout17 net23 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xro_inst.gcount\[2\].div_flop ro_inst.counter_n\[2\] net305 ro_inst.counter_n\[1\]
+ ro_inst.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_371_ cm_inst.cc_inst.out_notouch_\[163\] cm_inst.cc_inst.out_notouch_\[171\] cm_inst.cc_inst.out_notouch_\[179\]
+ cm_inst.cc_inst.out_notouch_\[187\] _115_ _116_ _141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_440_ _067_ _200_ _205_ _206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_23_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout207 net208 net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout229 net230 net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout218 net219 net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xcm_inst.cc_inst.invz_4_inst net34 net21 cm_inst.cc_inst.out_notouch_\[174\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__invz_4
XTAP_TAPCELL_ROW_20_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_354_ _124_ _125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_423_ _085_ _184_ _189_ _017_ _190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_51_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_285_ _048_ _053_ _056_ _057_ _058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_23_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 in[6] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__288__A2 _045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_337_ _018_ _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xcm_inst.cc_inst.latrnq_1_inst net270 net183 net112 cm_inst.cc_inst.out_notouch_\[126\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_406_ _067_ _168_ _173_ _174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_268_ cm_inst.cc_inst.out_notouch_\[160\] cm_inst.cc_inst.out_notouch_\[168\] cm_inst.cc_inst.out_notouch_\[176\]
+ cm_inst.cc_inst.out_notouch_\[184\] _038_ _040_ _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout25_I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xcm_inst.cc_inst.bufz_3_inst net24 net17 cm_inst.cc_inst.out_notouch_\[171\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__bufz_3
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcm_inst.cc_inst.inv_20_inst net204 cm_inst.cc_inst.out_notouch_\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_20
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.nor4_4_inst net261 net176 net106 net55 cm_inst.cc_inst.out_notouch_\[44\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_1_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.dffq_1_inst net172 net258 cm_inst.cc_inst.out_notouch_\[147\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout18 net22 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout29 net32 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.nand4_4_inst net208 net136 net73 net38 cm_inst.cc_inst.out_notouch_\[35\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_370_ _067_ _132_ _139_ _140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.oai211_4_inst net242 net159 net95 net49 cm_inst.cc_inst.out_notouch_\[98\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_46_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_499_ _005_ net314 cm_inst.page\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout208 net209 net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout219 net220 net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_20_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xro_inst.sig_cmp ro_inst.signal ro_inst.saved_signal ro_inst.running vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_43_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_422_ _186_ _188_ _066_ _189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_284_ _048_ _055_ cm_inst.cc_inst.out_notouch_\[208\] _057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_353_ _069_ _046_ _124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_51_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.xor3_2_inst net277 net188 net115 cm_inst.cc_inst.out_notouch_\[64\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__302__I _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 in[7] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__323__S _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_267_ _039_ _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_405_ _170_ _172_ _138_ _173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_336_ cm_inst.cc_inst.out_notouch_\[98\] cm_inst.cc_inst.out_notouch_\[106\] cm_inst.cc_inst.out_notouch_\[114\]
+ cm_inst.cc_inst.out_notouch_\[122\] _105_ _106_ _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout18_I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.gcount\[28\].div_flop_inv ro_inst.counter\[28\] ro_inst.counter_n\[28\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xro_inst.slow_clock_inv net306 ro_inst.slow_clk_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_6_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_319_ cm_inst.cc_inst.out_notouch_\[161\] cm_inst.cc_inst.out_notouch_\[169\] cm_inst.cc_inst.out_notouch_\[177\]
+ cm_inst.cc_inst.out_notouch_\[185\] _089_ _090_ _091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xcm_inst.cc_inst.clkbuf_20_inst net247 cm_inst.cc_inst.out_notouch_\[195\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
Xro_inst.gcount\[25\].div_flop ro_inst.counter_n\[25\] net308 ro_inst.counter_n\[24\]
+ ro_inst.counter\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_47_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.oai31_2_inst net277 net188 net115 net60 cm_inst.cc_inst.out_notouch_\[88\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_47_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.dlyd_1_inst net261 cm_inst.cc_inst.out_notouch_\[185\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_0_7_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout19 net22 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.dffnq_2_inst net149 net230 cm_inst.cc_inst.out_notouch_\[136\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XFILLER_0_23_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_498_ _004_ net313 cm_inst.page\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.clkinv_4_inst net249 cm_inst.cc_inst.out_notouch_\[199\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
Xfanout209 net216 net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_421_ _079_ _187_ _188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_283_ _055_ cm_inst.cc_inst.out_notouch_\[200\] _056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_352_ _121_ _122_ _032_ _123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.and4_4_inst net250 net167 net102 net58 cm_inst.cc_inst.out_notouch_\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_4
X_404_ _080_ _171_ _172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xro_inst.ring_osc_0 ro_inst.ring\[0\] ro_inst.enable ro_inst.ring\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_38_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_266_ cm_inst.page\[1\] _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_335_ _020_ _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xro_inst.gcount\[15\].div_flop ro_inst.counter_n\[15\] net294 ro_inst.counter_n\[14\]
+ ro_inst.counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_22_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.aoi211_4_inst net285 net195 net123 net64 cm_inst.cc_inst.out_notouch_\[74\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__499__CLK net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xcm_inst.cc_inst.latq_4_inst net275 net185 cm_inst.cc_inst.out_notouch_\[125\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
Xcm_inst.cc_inst.tieh_inst cm_inst.cc_inst.out_notouch_\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_33_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_318_ _026_ _090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_249_ cm_inst.cc_inst.out_notouch_\[96\] cm_inst.cc_inst.out_notouch_\[104\] cm_inst.cc_inst.out_notouch_\[112\]
+ cm_inst.cc_inst.out_notouch_\[120\] _019_ _021_ _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xcm_inst.cc_inst.dffnrnq_1_inst net190 net124 net282 cm_inst.cc_inst.out_notouch_\[138\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XANTENNA_fanout30_I net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi22_1_inst_B2 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout78_I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.or3_1_inst net269 net182 net111 cm_inst.cc_inst.out_notouch_\[48\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_14_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__481__A2 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.latrnq_4_inst net230 net149 net86 cm_inst.cc_inst.out_notouch_\[128\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latrnq_4
Xro_inst.gcount\[6\].div_flop_inv ro_inst.counter\[6\] ro_inst.counter_n\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_497_ _003_ net313 cm_inst.page\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_351_ cm_inst.cc_inst.out_notouch_\[130\] cm_inst.cc_inst.out_notouch_\[138\] cm_inst.cc_inst.out_notouch_\[146\]
+ cm_inst.cc_inst.out_notouch_\[154\] _108_ _109_ _122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_420_ cm_inst.cc_inst.out_notouch_\[38\] cm_inst.cc_inst.out_notouch_\[46\] cm_inst.cc_inst.out_notouch_\[54\]
+ cm_inst.cc_inst.out_notouch_\[62\] _050_ _068_ _187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_51_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_282_ _054_ _055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xro_inst.gcount\[31\].div_flop_inv ro_inst.counter\[31\] ro_inst.counter_n\[31\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout245_I net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xro_inst.gcount\[1\].div_flop ro_inst.counter_n\[1\] net305 ro_inst.counter_n\[0\]
+ ro_inst.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_10_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout60_I net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_403_ cm_inst.cc_inst.out_notouch_\[69\] cm_inst.cc_inst.out_notouch_\[77\] cm_inst.cc_inst.out_notouch_\[85\]
+ cm_inst.cc_inst.out_notouch_\[93\] _081_ _082_ _171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_334_ _037_ _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xro_inst.ring_osc_1 ro_inst.ring\[1\] ro_inst.ring\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_265_ _037_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__268__S1 _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_317_ _049_ _089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_33_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout110_I net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_248_ _020_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xcm_inst.cc_inst.dffq_4_inst net177 net263 cm_inst.cc_inst.out_notouch_\[149\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_38_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout190 net192 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xro_inst.gcount\[24\].div_flop_inv ro_inst.counter\[24\] ro_inst.counter_n\[24\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_29_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SI net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__398__S0 _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_496_ _002_ net313 cm_inst.page\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xro_inst.gcount\[34\].div_flop ro_inst.counter_n\[34\] net311 ro_inst.counter_n\[33\]
+ ro_inst.counter\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_37_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.sdffrnq_1_inst net157 net93 net47 net31 net240 cm_inst.cc_inst.out_notouch_\[162\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1
XANTENNA__443__S _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_350_ cm_inst.cc_inst.out_notouch_\[162\] cm_inst.cc_inst.out_notouch_\[170\] cm_inst.cc_inst.out_notouch_\[178\]
+ cm_inst.cc_inst.out_notouch_\[186\] _105_ _106_ _121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_51_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xro_inst.gcount\[17\].div_flop_inv ro_inst.counter\[17\] ro_inst.counter_n\[17\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_281_ _018_ _054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_479_ _228_ net40 _234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xro_inst.ring_osc_2 ro_inst.ring\[2\] ro_inst.ring\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_264_ cm_inst.page\[0\] _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_333_ _104_ net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_402_ _076_ _169_ _170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout188_I net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.clkbuf_2_inst net281 cm_inst.cc_inst.out_notouch_\[189\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xcm_inst.cc_inst.dlyd_4_inst net257 cm_inst.cc_inst.out_notouch_\[187\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_33_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_247_ cm_inst.page\[1\] _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_316_ _033_ _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_cm_inst.cc_inst.and4_4_inst_A3 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout191 net192 net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout180 net181 net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_29_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xro_inst.gcount\[24\].div_flop ro_inst.counter_n\[24\] net308 ro_inst.counter_n\[23\]
+ ro_inst.counter\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_14_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.dffrnq_1_inst net184 net113 net272 cm_inst.cc_inst.out_notouch_\[150\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_17_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__398__S1 _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.buf_8_inst net271 cm_inst.cc_inst.out_notouch_\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_35_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_495_ _001_ net303 cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_45_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.buf_12_inst net224 cm_inst.cc_inst.out_notouch_\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_280_ _052_ cm_inst.cc_inst.out_notouch_\[192\] _053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_51_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__298__S0 _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_478_ _233_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcm_inst.cc_inst.dffnrnq_4_inst net144 net85 net224 cm_inst.cc_inst.out_notouch_\[140\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4
Xro_inst.gcount\[2\].div_flop_inv ro_inst.counter\[2\] ro_inst.counter_n\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__253__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_401_ cm_inst.cc_inst.out_notouch_\[101\] cm_inst.cc_inst.out_notouch_\[109\] cm_inst.cc_inst.out_notouch_\[117\]
+ cm_inst.cc_inst.out_notouch_\[125\] _019_ _023_ _169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_332_ _103_ ro_inst.counter\[1\] _063_ _104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_263_ _033_ _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SI net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xcm_inst.cc_inst.or3_4_inst net262 net174 net105 cm_inst.cc_inst.out_notouch_\[50\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_0_41_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_315_ _067_ _075_ _086_ _087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_26_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_246_ _018_ _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xro_inst.gcount\[14\].div_flop ro_inst.counter_n\[14\] net294 ro_inst.counter_n\[13\]
+ ro_inst.counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_46_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout192 net197 net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout170 net171 net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout181 net199 net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_29_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.xor2_1_inst net260 net175 cm_inst.cc_inst.out_notouch_\[60\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout163_I net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xro_inst.gcount\[20\].div_flop_inv ro_inst.counter\[20\] ro_inst.counter_n\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_cm_inst.cc_inst.icgtn_1_inst_TE net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_29_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_13_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_494_ _000_ net303 cm_inst.page\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__298__S1 _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout126_I net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_477_ net5 net80 _226_ _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SI net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout39_I net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_400_ _166_ _167_ _074_ _168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_331_ _065_ _087_ _101_ _102_ _103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_36_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_262_ _017_ _034_ _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xcm_inst.cc_inst.aoi21_2_inst net226 net146 net82 cm_inst.cc_inst.out_notouch_\[67\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xro_inst.gcount\[13\].div_flop_inv ro_inst.counter\[13\] ro_inst.counter_n\[13\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_314_ _078_ _084_ _085_ _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_245_ cm_inst.page\[0\] _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_15_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_43_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__259__I _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout193 net194 net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout182 net183 net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout171 net181 net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout160 net161 net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_29_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.sdffrnq_4_inst net156 net93 net47 net30 net237 cm_inst.cc_inst.out_notouch_\[164\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4
XFILLER_0_47_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout21_I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_493_ _241_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcm_inst.cc_inst.hold_inst cm_inst.cc_inst.out_notouch_\[173\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__hold
XFILLER_0_41_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__383__S _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_37_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.mux2_2_inst net275 net183 net112 cm_inst.cc_inst.out_notouch_\[118\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_476_ _232_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.gcount\[33\].div_flop ro_inst.counter_n\[33\] net311 ro_inst.counter_n\[32\]
+ ro_inst.counter\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_330_ cm_inst.page\[5\] _102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_261_ _022_ _024_ _028_ _029_ _032_ _033_ _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_8_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_459_ net3 _222_ _223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.dlya_2_inst net283 cm_inst.cc_inst.out_notouch_\[177\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.inv_16_inst net268 cm_inst.cc_inst.out_notouch_\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_16
XANTENNA_fanout51_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_313_ _066_ _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_244_ cm_inst.page\[4\] _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xcm_inst.cc_inst.dffrnq_4_inst net145 net86 net225 cm_inst.cc_inst.out_notouch_\[152\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XTAP_TAPCELL_ROW_15_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__275__I _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout172 net180 net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout150 net162 net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout161 net162 net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout183 net184 net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout194 net195 net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout101_I net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xro_inst.clock_gate ro_inst.ring\[0\] ro_inst.running net315 ro_inst.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XFILLER_0_18_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_492_ net5 ro_sel\[2\] _238_ _241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.sdffq_2_inst net149 net87 net44 net230 cm_inst.cc_inst.out_notouch_\[160\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffq_2
XTAP_TAPCELL_ROW_37_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.invz_12_inst net104 net53 cm_inst.cc_inst.out_notouch_\[175\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_12
XFILLER_0_40_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xro_inst.gcount\[23\].div_flop ro_inst.counter_n\[23\] net306 ro_inst.counter_n\[22\]
+ ro_inst.counter\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout81_I net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.clkbuf_16_inst net220 cm_inst.cc_inst.out_notouch_\[194\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_42_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.oai32_2_inst net227 net146 net82 net42 net26 cm_inst.cc_inst.out_notouch_\[91\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_475_ net4 net141 _230_ _232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__278__I _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_260_ cm_inst.page\[3\] _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xcm_inst.cc_inst.inv_3_inst net251 cm_inst.cc_inst.out_notouch_\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_8_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_458_ _220_ _222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_389_ _085_ _152_ _157_ _017_ _158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_27_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout310 net312 net310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_312_ _080_ _083_ _084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_243_ cm_inst.page\[5\] _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xcm_inst.cc_inst.xor2_4_inst net253 net169 cm_inst.cc_inst.out_notouch_\[62\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XTAP_TAPCELL_ROW_9_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout173 net180 net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout195 net196 net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout140 net143 net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout162 net163 net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout151 net155 net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout184 net189 net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.gcount\[13\].div_flop ro_inst.counter_n\[13\] net295 ro_inst.counter_n\[12\]
+ ro_inst.counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_29_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.sig_latch ro_inst.signal ro_inst.slow_clk_n ro_inst.saved_signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_491_ _240_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_474_ _231_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcm_inst.cc_inst.or4_1_inst net205 net133 net73 net38 cm_inst.cc_inst.out_notouch_\[51\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_22_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.addh_1_inst net234 net153 cm_inst.cc_inst.out_notouch_\[111\] cm_inst.cc_inst.out_notouch_\[112\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__addh_1
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_457_ _220_ _221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_388_ _154_ _156_ _138_ _157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xfanout311 net312 net311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout300 net301 net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_311_ cm_inst.cc_inst.out_notouch_\[65\] cm_inst.cc_inst.out_notouch_\[73\] cm_inst.cc_inst.out_notouch_\[81\]
+ cm_inst.cc_inst.out_notouch_\[89\] _081_ _082_ _083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_9_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_509_ _015_ net302 ro_sel\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_15_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.latrsnq_1_inst net282 net190 net119 net63 cm_inst.cc_inst.out_notouch_\[129\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latrsnq_1
XFILLER_0_46_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_5_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.icgtn_1_inst net221 net141 net81 cm_inst.cc_inst.out_notouch_\[204\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__icgtn_1
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout196 net197 net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout174 net175 net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout185 net187 net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout163 net200 net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout130 net131 net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout141 net143 net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout152 net155 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout289_I net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.clkbuf_8_inst net218 cm_inst.cc_inst.out_notouch_\[192\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_490_ net4 ro_sel\[1\] _238_ _240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xro_inst.clock_gate_inv ro_inst.counter\[0\] ro_inst.counter_n\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_8_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_34_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_473_ net3 net222 _230_ _231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_50_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.nor2_2_inst net210 net129 cm_inst.cc_inst.out_notouch_\[37\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_42_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.nand2_2_inst net251 net167 cm_inst.cc_inst.out_notouch_\[28\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xro_inst.gcount\[9\].div_flop_inv ro_inst.counter\[9\] ro_inst.counter_n\[9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_456_ _217_ _218_ _219_ net2 _220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA_fanout117_I net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_387_ _079_ _155_ _156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout312 net313 net312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout301 net302 net301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_310_ _039_ _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xro_inst.gcount\[34\].div_flop_inv ro_inst.counter\[34\] ro_inst.counter_n\[34\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_9_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_37_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xro_inst.gcount\[32\].div_flop ro_inst.counter_n\[32\] net310 ro_inst.counter_n\[31\]
+ ro_inst.counter\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_15_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_508_ _014_ net301 ro_sel\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_439_ _202_ _204_ _138_ _205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_21_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout120 net125 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout131 net132 net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout175 net176 net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout197 net198 net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout164 net166 net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_6_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout142 net143 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout153 net155 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout186 net187 net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.buf_1_inst net271 cm_inst.cc_inst.out_notouch_\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout184_I net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__477__I1 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.oai21_2_inst net286 net193 net121 cm_inst.cc_inst.out_notouch_\[82\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_39_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xro_inst.gcount\[27\].div_flop_inv ro_inst.counter\[27\] ro_inst.counter_n\[27\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_472_ _226_ _230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_50_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.invz_3_inst net123 net65 cm_inst.cc_inst.out_notouch_\[174\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
Xcm_inst.cc_inst.sdffrsnq_2_inst net194 net124 net64 net34 net20 net285 cm_inst.cc_inst.out_notouch_\[166\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2
XFILLER_0_45_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_386_ cm_inst.cc_inst.out_notouch_\[36\] cm_inst.cc_inst.out_notouch_\[44\] cm_inst.cc_inst.out_notouch_\[52\]
+ cm_inst.cc_inst.out_notouch_\[60\] _092_ _116_ _155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xro_inst.gcount\[22\].div_flop ro_inst.counter_n\[22\] net300 ro_inst.counter_n\[21\]
+ ro_inst.counter\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_455_ net8 _219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcm_inst.cc_inst.icgtp_2_inst net218 net141 net80 cm_inst.cc_inst.out_notouch_\[208\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__icgtp_2
XFILLER_0_18_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout313 net314 net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout302 net304 net302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xcm_inst.cc_inst.bufz_2_inst net103 net53 cm_inst.cc_inst.out_notouch_\[171\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__bufz_2
XFILLER_0_24_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_507_ _013_ net300 ro_sel\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_369_ _134_ _137_ _138_ _139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_438_ _080_ _203_ _204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout121 net122 net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout165 net166 net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout110 net127 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout132 net140 net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_6_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout143 net163 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout154 net155 net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout176 net179 net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout187 net189 net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xcm_inst.cc_inst.and2_2_inst net212 net138 cm_inst.cc_inst.out_notouch_\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xfanout198 net199 net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_49_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.or4_4_inst net203 net131 net71 net39 cm_inst.cc_inst.out_notouch_\[53\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_20_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.addh_4_inst net233 net151 cm_inst.cc_inst.out_notouch_\[115\] cm_inst.cc_inst.out_notouch_\[116\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__addh_4
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.xnor2_2_inst net205 net133 cm_inst.cc_inst.out_notouch_\[55\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_8_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.gcount\[12\].div_flop ro_inst.counter_n\[12\] net296 ro_inst.counter_n\[11\]
+ ro_inst.counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_471_ _219_ _228_ _229_ _221_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SI net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.latrsnq_4_inst net258 net172 net103 net53 cm_inst.cc_inst.out_notouch_\[131\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latrsnq_4
Xcm_inst.cc_inst.xor3_1_inst net205 net133 net73 cm_inst.cc_inst.out_notouch_\[63\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.clkinv_20_inst net247 cm_inst.cc_inst.out_notouch_\[203\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_20
XFILLER_0_32_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.icgtn_4_inst net249 net165 net100 cm_inst.cc_inst.out_notouch_\[206\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__icgtn_4
XFILLER_0_8_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_454_ net7 _218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_385_ _076_ _153_ _154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout314 net1 net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout303 net304 net303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_506_ _012_ net307 ro_inst.enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_299_ _050_ _071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xro_inst.gcount\[5\].div_flop_inv ro_inst.counter\[5\] ro_inst.counter_n\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_437_ cm_inst.cc_inst.out_notouch_\[71\] cm_inst.cc_inst.out_notouch_\[79\] cm_inst.cc_inst.out_notouch_\[87\]
+ cm_inst.cc_inst.out_notouch_\[95\] _135_ _106_ _203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_23_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_368_ cm_inst.page\[3\] _138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout35_I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout177 net179 net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout122 net123 net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout100 net101 net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout199 net200 net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout188 net189 net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout166 net171 net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout144 net148 net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_6_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout133 net134 net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout155 net161 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout111 net113 net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xro_inst.gcount\[30\].div_flop_inv ro_inst.counter\[30\] ro_inst.counter_n\[30\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.aoi22_2_inst net287 net193 net121 net64 cm_inst.cc_inst.out_notouch_\[70\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_17_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcm_inst.cc_inst.oai31_1_inst net233 net152 net91 net45 cm_inst.cc_inst.out_notouch_\[87\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_25_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xro_inst.gcount\[9\].div_flop ro_inst.counter_n\[9\] net297 ro_inst.counter_n\[8\]
+ ro_inst.counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_22_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.dffnq_1_inst net165 net248 cm_inst.cc_inst.out_notouch_\[135\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA_input7_I in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.clkinv_3_inst net253 cm_inst.cc_inst.out_notouch_\[198\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_12_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_470_ _016_ _229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xro_inst.gcount\[23\].div_flop_inv ro_inst.counter\[23\] ro_inst.counter_n\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_453_ net6 _217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_384_ cm_inst.cc_inst.out_notouch_\[4\] cm_inst.cc_inst.out_notouch_\[12\] cm_inst.cc_inst.out_notouch_\[20\]
+ cm_inst.cc_inst.out_notouch_\[28\] _089_ _027_ _153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.buf_4_inst net210 cm_inst.cc_inst.out_notouch_\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout304 net314 net304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_505_ _011_ net304 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_436_ _112_ _201_ _202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_298_ cm_inst.cc_inst.out_notouch_\[33\] cm_inst.cc_inst.out_notouch_\[41\] cm_inst.cc_inst.out_notouch_\[49\]
+ cm_inst.cc_inst.out_notouch_\[57\] _051_ _069_ _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_367_ _080_ _136_ _137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__498__CLK net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__409__S _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout28_I net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout178 net179 net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout123 net124 net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout112 net113 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout167 net170 net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout101 net102 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout189 net198 net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout134 net137 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout145 net148 net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_6_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout156 net157 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xro_inst.gcount\[16\].div_flop_inv ro_inst.counter\[16\] ro_inst.counter_n\[16\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_25_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_419_ _112_ _185_ _186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.gcount\[31\].div_flop ro_inst.counter_n\[31\] net310 ro_inst.counter_n\[30\]
+ ro_inst.counter\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xcm_inst.cc_inst.dlyb_2_inst net237 cm_inst.cc_inst.out_notouch_\[180\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlyb_2
XTAP_TAPCELL_ROW_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.oai221_2_inst net233 net152 net91 net45 net26 cm_inst.cc_inst.out_notouch_\[100\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_TAPCELL_ROW_22_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout312_I net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout58_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai31_4_inst_B net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_383_ _150_ _151_ _044_ _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_452_ _216_ ro_inst.signal vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.latsnq_2_inst net264 net178 net108 cm_inst.cc_inst.out_notouch_\[133\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latsnq_2
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout305 net307 net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_52_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__353__A1 _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__340__S _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_366_ cm_inst.cc_inst.out_notouch_\[67\] cm_inst.cc_inst.out_notouch_\[75\] cm_inst.cc_inst.out_notouch_\[83\]
+ cm_inst.cc_inst.out_notouch_\[91\] _135_ _042_ _136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_504_ _010_ net303 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_435_ cm_inst.cc_inst.out_notouch_\[103\] cm_inst.cc_inst.out_notouch_\[111\] cm_inst.cc_inst.out_notouch_\[119\]
+ cm_inst.cc_inst.out_notouch_\[127\] _025_ _021_ _201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_297_ _068_ _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.oai33_2_inst net287 net193 net121 net62 net35 net21 cm_inst.cc_inst.out_notouch_\[94\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_2
XFILLER_0_3_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout102 net110 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xro_inst.gcount\[21\].div_flop ro_inst.counter_n\[21\] net299 ro_inst.counter_n\[20\]
+ ro_inst.counter\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout113 net118 net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout179 net180 net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout124 net125 net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout168 net169 net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout135 net136 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout146 net148 net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout157 net160 net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__326__A1 _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_418_ cm_inst.cc_inst.out_notouch_\[6\] cm_inst.cc_inst.out_notouch_\[14\] cm_inst.cc_inst.out_notouch_\[22\]
+ cm_inst.cc_inst.out_notouch_\[30\] _089_ _027_ _185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_349_ _085_ _111_ _119_ _017_ _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_36_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xro_inst.gcount\[1\].div_flop_inv ro_inst.counter\[1\] ro_inst.counter_n\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout40_I net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcm_inst.cc_inst.xor3_4_inst net213 net139 net78 cm_inst.cc_inst.out_notouch_\[65\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_4
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout292_I net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SETN net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_cm_inst.cc_inst.icgtp_2_inst_TE net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_382_ cm_inst.cc_inst.out_notouch_\[68\] cm_inst.cc_inst.out_notouch_\[76\] cm_inst.cc_inst.out_notouch_\[84\]
+ cm_inst.cc_inst.out_notouch_\[92\] _135_ _042_ _151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_451_ _214_ _215_ ro_sel\[2\] _216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcm_inst.cc_inst.aoi221_2_inst net229 net149 net84 net42 net26 cm_inst.cc_inst.out_notouch_\[76\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_26_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.gcount\[11\].div_flop ro_inst.counter_n\[11\] net296 ro_inst.counter_n\[10\]
+ ro_inst.counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout306 net307 net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.clkbuf_1_inst net237 cm_inst.cc_inst.out_notouch_\[188\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_503_ _009_ net303 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_296_ _026_ _068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_434_ _198_ _199_ _074_ _200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcm_inst.cc_inst.oai31_4_inst net212 net138 net77 net41 cm_inst.cc_inst.out_notouch_\[89\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_365_ _037_ _135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout125 net126 net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout103 net109 net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout114 net117 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout136 net137 net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_6_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout147 net148 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout169 net170 net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout158 net160 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.dffnq_4_inst net178 net263 cm_inst.cc_inst.out_notouch_\[137\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_4
XFILLER_0_36_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_417_ _182_ _183_ _032_ _184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_348_ _114_ _118_ _066_ _119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_11_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_279_ _051_ _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout33_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xcm_inst.cc_inst.inv_12_inst net224 cm_inst.cc_inst.out_notouch_\[15\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_12
XFILLER_0_52_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xro_inst.gcount\[12\].div_flop_inv ro_inst.counter\[12\] ro_inst.counter_n\[12\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xro_inst.gcount\[8\].div_flop ro_inst.counter_n\[8\] net297 ro_inst.counter_n\[7\]
+ ro_inst.counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input5_I in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_381_ cm_inst.cc_inst.out_notouch_\[100\] cm_inst.cc_inst.out_notouch_\[108\] cm_inst.cc_inst.out_notouch_\[116\]
+ cm_inst.cc_inst.out_notouch_\[124\] _038_ _040_ _150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_450_ _164_ _180_ _196_ _212_ ro_sel\[0\] ro_sel\[1\] _215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__442__S0 _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout307 net312 net307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_433_ cm_inst.cc_inst.out_notouch_\[7\] cm_inst.cc_inst.out_notouch_\[15\] cm_inst.cc_inst.out_notouch_\[23\]
+ cm_inst.cc_inst.out_notouch_\[31\] _081_ _082_ _199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_502_ _008_ net301 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_cm_inst.cc_inst.oai33_2_inst_B2 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__424__S0 _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_295_ _066_ _067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_364_ _112_ _133_ _134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcm_inst.cc_inst.clkbuf_12_inst net211 cm_inst.cc_inst.out_notouch_\[193\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XANTENNA_fanout198_I net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__415__S0 _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout104 net109 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout115 net117 net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout126 net127 net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout148 net150 net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout137 net139 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout159 net160 net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xcm_inst.cc_inst.nor3_2_inst net268 net182 net111 cm_inst.cc_inst.out_notouch_\[40\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_52_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xcm_inst.cc_inst.dffnsnq_2_inst net177 net107 net264 cm_inst.cc_inst.out_notouch_\[145\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2
XFILLER_0_49_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.nand3_2_inst net207 net135 net76 cm_inst.cc_inst.out_notouch_\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_416_ cm_inst.cc_inst.out_notouch_\[70\] cm_inst.cc_inst.out_notouch_\[78\] cm_inst.cc_inst.out_notouch_\[86\]
+ cm_inst.cc_inst.out_notouch_\[94\] _108_ _109_ _183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_278_ _050_ _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_11_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout113_I net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_347_ _079_ _117_ _118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__341__I _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xcm_inst.cc_inst.bufz_8_inst net93 net47 cm_inst.cc_inst.out_notouch_\[172\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_0_18_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__483__A2 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_16_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__272__S _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__246__I _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xro_inst.gcount\[30\].div_flop ro_inst.counter_n\[30\] net309 ro_inst.counter_n\[29\]
+ ro_inst.counter\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_12_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_380_ _149_ net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcm_inst.cc_inst.oai22_2_inst net220 net142 net79 net40 cm_inst.cc_inst.out_notouch_\[85\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcm_inst.cc_inst.aoi21_1_inst net285 net195 net123 cm_inst.cc_inst.out_notouch_\[66\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout308 net310 net308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
.ends

