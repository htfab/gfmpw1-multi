VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cells9
  CLASS BLOCK ;
  FOREIGN cells9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END clk
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 82.550995 ;
    ANTENNADIFFAREA 20.746799 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END in[0]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 0.000 7.280 4.000 ;
    END
  END in[11]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 4.000 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 0.000 20.720 4.000 ;
    END
  END in[15]
  PIN in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END in[16]
  PIN in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END in[17]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.900000 ;
    ANTENNADIFFAREA 1.220400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 1.220400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 4.000 182.000 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 1.220400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 296.000 138.320 300.000 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.560500 ;
    ANTENNADIFFAREA 1.220400 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 296.000 148.400 300.000 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.638500 ;
    ANTENNADIFFAREA 1.220400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.240 4.000 198.800 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.638500 ;
    ANTENNADIFFAREA 1.220400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.638500 ;
    ANTENNADIFFAREA 1.220400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END in[9]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.911900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.290400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.720 4.000 259.280 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.290400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 4.000 34.160 ;
    END
  END out[11]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.840 4.000 148.400 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.360 4.000 171.920 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.290400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 4.000 30.800 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.290400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 268.800 300.000 269.360 ;
    END
  END out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 19.860 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 19.860 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 19.860 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 19.860 254.240 282.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 19.710 292.880 282.690 ;
      LAYER Metal2 ;
        RECT 8.540 295.700 137.460 296.660 ;
        RECT 138.620 295.700 147.540 296.660 ;
        RECT 148.700 295.700 291.060 296.660 ;
        RECT 8.540 19.970 291.060 295.700 ;
      LAYER Metal3 ;
        RECT 4.000 269.660 296.000 282.380 ;
        RECT 4.000 268.500 295.700 269.660 ;
        RECT 4.000 259.580 296.000 268.500 ;
        RECT 4.300 258.420 296.000 259.580 ;
        RECT 4.000 222.620 296.000 258.420 ;
        RECT 4.300 221.460 296.000 222.620 ;
        RECT 4.000 199.100 296.000 221.460 ;
        RECT 4.300 197.940 296.000 199.100 ;
        RECT 4.000 195.740 296.000 197.940 ;
        RECT 4.300 194.580 296.000 195.740 ;
        RECT 4.000 189.020 296.000 194.580 ;
        RECT 4.300 187.860 296.000 189.020 ;
        RECT 4.000 185.660 296.000 187.860 ;
        RECT 4.300 184.500 296.000 185.660 ;
        RECT 4.000 182.300 296.000 184.500 ;
        RECT 4.300 181.140 296.000 182.300 ;
        RECT 4.000 172.220 296.000 181.140 ;
        RECT 4.300 171.060 296.000 172.220 ;
        RECT 4.000 165.500 296.000 171.060 ;
        RECT 4.300 164.340 296.000 165.500 ;
        RECT 4.000 162.140 296.000 164.340 ;
        RECT 4.300 160.980 296.000 162.140 ;
        RECT 4.000 158.780 296.000 160.980 ;
        RECT 4.300 157.620 296.000 158.780 ;
        RECT 4.000 155.420 296.000 157.620 ;
        RECT 4.300 154.260 296.000 155.420 ;
        RECT 4.000 152.060 296.000 154.260 ;
        RECT 4.300 150.900 296.000 152.060 ;
        RECT 4.000 148.700 296.000 150.900 ;
        RECT 4.300 147.540 296.000 148.700 ;
        RECT 4.000 145.340 296.000 147.540 ;
        RECT 4.300 144.180 296.000 145.340 ;
        RECT 4.000 34.460 296.000 144.180 ;
        RECT 4.300 33.300 296.000 34.460 ;
        RECT 4.000 31.100 296.000 33.300 ;
        RECT 4.300 29.940 296.000 31.100 ;
        RECT 4.000 20.020 296.000 29.940 ;
      LAYER Metal4 ;
        RECT 117.740 75.690 175.540 219.430 ;
        RECT 177.740 75.690 191.380 219.430 ;
  END
END cells9
END LIBRARY

