* NGSPICE file created from loopback.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

.subckt loopback clk in[0] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17]
+ in[18] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] out[0] out[10] out[11]
+ out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] rst_n vdd vss
XPHY_EDGE_ROW_0_Left_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput31 net31 out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput32 net32 out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input11_I in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 net21 out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input3_I in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_4_Left_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput23 net23 out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_29_ net3 net4 net26 _09_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_1_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_28_ _08_ net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput24 net24 out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_2_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input1_I in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27_ net3 net26 _08_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput25 net25 out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_2_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_43_ clk net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26_ _07_ net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xoutput26 net26 out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_42_ _15_ net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Left_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25_ net19 net2 net24 _07_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_7_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput27 net27 out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_41_ net9 net10 net32 _15_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_10_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24_ _06_ net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput28 net28 out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input18_I in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_40_ _14_ net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_10_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23_ net19 net24 _06_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput29 net29 out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22_ _05_ net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21_ net17 _03_ _04_ _05_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_3_Left_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input8_I in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20_ net13 net15 _04_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xinput1 in[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 in[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_6_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_7_Left_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 in[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input14_I in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 in[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_10_Left_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput5 in[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput6 in[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput20 rst_n net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input12_I in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput7 in[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput10 in[18] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 in[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_2_Left_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_39_ net9 net32 _14_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xinput11 in[1] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput9 in[17] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput12 in[2] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_38_ _13_ net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_4_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_37_ net7 net8 net30 _13_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xinput13 in[3] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_6_Left_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput14 in[4] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_36_ _12_ net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19_ _00_ _01_ _02_ _03_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_9_Left_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_11_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_35_ net7 net30 _12_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xinput15 in[5] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18_ net14 net16 _02_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_34_ _11_ net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17_ net1 net20 _01_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xinput16 in[6] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input19_I in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_33_ net5 net6 net28 _11_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xinput17 in[7] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16_ net11 net12 net18 _00_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_9_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__43__I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_32_ _10_ net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput18 in[8] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_31_ net5 net28 _10_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_1_Left_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput19 in[9] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input17_I in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_30_ _09_ net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_5_Left_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input7_I in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input15_I in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input20_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input5_I in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input13_I in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput30 net30 out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
.ends

