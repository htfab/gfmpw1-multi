magic
tech gf180mcuD
magscale 1 10
timestamp 1702354384
<< metal1 >>
rect 1344 60394 62608 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 62608 60394
rect 1344 60308 62608 60342
rect 17950 60226 18002 60238
rect 17950 60162 18002 60174
rect 48974 60226 49026 60238
rect 48974 60162 49026 60174
rect 27570 60062 27582 60114
rect 27634 60062 27646 60114
rect 34974 60002 35026 60014
rect 15362 59950 15374 60002
rect 15426 59950 15438 60002
rect 16930 59950 16942 60002
rect 16994 59950 17006 60002
rect 28578 59950 28590 60002
rect 28642 59950 28654 60002
rect 33954 59950 33966 60002
rect 34018 59950 34030 60002
rect 47954 59950 47966 60002
rect 48018 59950 48030 60002
rect 34974 59938 35026 59950
rect 13582 59890 13634 59902
rect 13582 59826 13634 59838
rect 13806 59890 13858 59902
rect 13806 59826 13858 59838
rect 19966 59890 20018 59902
rect 19966 59826 20018 59838
rect 20862 59890 20914 59902
rect 20862 59826 20914 59838
rect 23214 59890 23266 59902
rect 23214 59826 23266 59838
rect 23774 59890 23826 59902
rect 23774 59826 23826 59838
rect 23886 59890 23938 59902
rect 23886 59826 23938 59838
rect 27358 59890 27410 59902
rect 27358 59826 27410 59838
rect 31166 59890 31218 59902
rect 31166 59826 31218 59838
rect 33070 59890 33122 59902
rect 33070 59826 33122 59838
rect 38558 59890 38610 59902
rect 38558 59826 38610 59838
rect 14142 59778 14194 59790
rect 14814 59778 14866 59790
rect 14466 59726 14478 59778
rect 14530 59726 14542 59778
rect 14142 59714 14194 59726
rect 14814 59714 14866 59726
rect 15374 59778 15426 59790
rect 15374 59714 15426 59726
rect 15934 59778 15986 59790
rect 15934 59714 15986 59726
rect 16158 59778 16210 59790
rect 16158 59714 16210 59726
rect 16270 59778 16322 59790
rect 16270 59714 16322 59726
rect 16382 59778 16434 59790
rect 16382 59714 16434 59726
rect 20078 59778 20130 59790
rect 20078 59714 20130 59726
rect 20302 59778 20354 59790
rect 20302 59714 20354 59726
rect 20974 59778 21026 59790
rect 20974 59714 21026 59726
rect 21198 59778 21250 59790
rect 24110 59778 24162 59790
rect 22082 59726 22094 59778
rect 22146 59726 22158 59778
rect 21198 59714 21250 59726
rect 24110 59714 24162 59726
rect 25006 59778 25058 59790
rect 32174 59778 32226 59790
rect 26338 59726 26350 59778
rect 26402 59726 26414 59778
rect 28354 59726 28366 59778
rect 28418 59726 28430 59778
rect 29810 59726 29822 59778
rect 29874 59726 29886 59778
rect 25006 59714 25058 59726
rect 32174 59714 32226 59726
rect 32286 59778 32338 59790
rect 32286 59714 32338 59726
rect 32398 59778 32450 59790
rect 32398 59714 32450 59726
rect 32622 59778 32674 59790
rect 32622 59714 32674 59726
rect 33182 59778 33234 59790
rect 34638 59778 34690 59790
rect 33730 59726 33742 59778
rect 33794 59726 33806 59778
rect 33182 59714 33234 59726
rect 34638 59714 34690 59726
rect 1344 59610 62608 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 62608 59610
rect 1344 59524 62608 59558
rect 14030 59442 14082 59454
rect 14030 59378 14082 59390
rect 16158 59442 16210 59454
rect 27470 59442 27522 59454
rect 22082 59390 22094 59442
rect 22146 59390 22158 59442
rect 16158 59378 16210 59390
rect 27470 59378 27522 59390
rect 30046 59442 30098 59454
rect 30046 59378 30098 59390
rect 49758 59442 49810 59454
rect 49758 59378 49810 59390
rect 62190 59330 62242 59342
rect 14914 59278 14926 59330
rect 14978 59278 14990 59330
rect 17938 59278 17950 59330
rect 18002 59278 18014 59330
rect 24322 59278 24334 59330
rect 24386 59278 24398 59330
rect 30818 59278 30830 59330
rect 30882 59278 30894 59330
rect 33730 59278 33742 59330
rect 33794 59278 33806 59330
rect 34178 59278 34190 59330
rect 34242 59278 34254 59330
rect 34738 59278 34750 59330
rect 34802 59278 34814 59330
rect 62190 59266 62242 59278
rect 35086 59218 35138 59230
rect 20514 59166 20526 59218
rect 20578 59166 20590 59218
rect 24546 59166 24558 59218
rect 24610 59166 24622 59218
rect 25554 59166 25566 59218
rect 25618 59166 25630 59218
rect 26450 59166 26462 59218
rect 26514 59166 26526 59218
rect 48738 59166 48750 59218
rect 48802 59166 48814 59218
rect 35086 59154 35138 59166
rect 16942 59106 16994 59118
rect 16942 59042 16994 59054
rect 23774 59106 23826 59118
rect 35534 59106 35586 59118
rect 29586 59054 29598 59106
rect 29650 59054 29662 59106
rect 23774 59042 23826 59054
rect 35534 59042 35586 59054
rect 36094 59106 36146 59118
rect 36094 59042 36146 59054
rect 19406 58994 19458 59006
rect 19406 58930 19458 58942
rect 23438 58994 23490 59006
rect 32622 58994 32674 59006
rect 26114 58942 26126 58994
rect 26178 58942 26190 58994
rect 23438 58930 23490 58942
rect 32622 58930 32674 58942
rect 33182 58994 33234 59006
rect 33182 58930 33234 58942
rect 33518 58994 33570 59006
rect 33518 58930 33570 58942
rect 1344 58826 62608 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 62608 58826
rect 1344 58740 62608 58774
rect 13470 58658 13522 58670
rect 13470 58594 13522 58606
rect 13806 58658 13858 58670
rect 24882 58606 24894 58658
rect 24946 58606 24958 58658
rect 29474 58606 29486 58658
rect 29538 58606 29550 58658
rect 33730 58606 33742 58658
rect 33794 58606 33806 58658
rect 13806 58594 13858 58606
rect 21982 58546 22034 58558
rect 20402 58494 20414 58546
rect 20466 58494 20478 58546
rect 21982 58482 22034 58494
rect 52110 58546 52162 58558
rect 52770 58494 52782 58546
rect 52834 58494 52846 58546
rect 52110 58482 52162 58494
rect 22542 58434 22594 58446
rect 24782 58434 24834 58446
rect 27022 58434 27074 58446
rect 31166 58434 31218 58446
rect 51326 58434 51378 58446
rect 17938 58382 17950 58434
rect 18002 58382 18014 58434
rect 18498 58382 18510 58434
rect 18562 58382 18574 58434
rect 19170 58382 19182 58434
rect 19234 58382 19246 58434
rect 19618 58382 19630 58434
rect 19682 58382 19694 58434
rect 22866 58382 22878 58434
rect 22930 58382 22942 58434
rect 24098 58382 24110 58434
rect 24162 58382 24174 58434
rect 24994 58382 25006 58434
rect 25058 58382 25070 58434
rect 27794 58382 27806 58434
rect 27858 58382 27870 58434
rect 29586 58382 29598 58434
rect 29650 58382 29662 58434
rect 31266 58382 31278 58434
rect 31330 58382 31342 58434
rect 22542 58370 22594 58382
rect 24782 58370 24834 58382
rect 27022 58370 27074 58382
rect 31166 58370 31218 58382
rect 51326 58370 51378 58382
rect 14030 58322 14082 58334
rect 50766 58322 50818 58334
rect 14690 58270 14702 58322
rect 14754 58270 14766 58322
rect 27682 58270 27694 58322
rect 27746 58270 27758 58322
rect 30146 58270 30158 58322
rect 30210 58270 30222 58322
rect 14030 58258 14082 58270
rect 50766 58258 50818 58270
rect 16494 58210 16546 58222
rect 16494 58146 16546 58158
rect 17166 58210 17218 58222
rect 17166 58146 17218 58158
rect 17838 58210 17890 58222
rect 17838 58146 17890 58158
rect 21310 58210 21362 58222
rect 26686 58210 26738 58222
rect 28590 58210 28642 58222
rect 36430 58210 36482 58222
rect 21634 58158 21646 58210
rect 21698 58158 21710 58210
rect 28242 58158 28254 58210
rect 28306 58158 28318 58210
rect 35186 58158 35198 58210
rect 35250 58158 35262 58210
rect 21310 58146 21362 58158
rect 26686 58146 26738 58158
rect 28590 58146 28642 58158
rect 36430 58146 36482 58158
rect 37102 58210 37154 58222
rect 37102 58146 37154 58158
rect 40798 58210 40850 58222
rect 40798 58146 40850 58158
rect 41134 58210 41186 58222
rect 41134 58146 41186 58158
rect 44382 58210 44434 58222
rect 44382 58146 44434 58158
rect 45166 58210 45218 58222
rect 45166 58146 45218 58158
rect 45614 58210 45666 58222
rect 45614 58146 45666 58158
rect 46062 58210 46114 58222
rect 46062 58146 46114 58158
rect 47630 58210 47682 58222
rect 47630 58146 47682 58158
rect 48078 58210 48130 58222
rect 48078 58146 48130 58158
rect 48526 58210 48578 58222
rect 48526 58146 48578 58158
rect 48974 58210 49026 58222
rect 48974 58146 49026 58158
rect 49422 58210 49474 58222
rect 49422 58146 49474 58158
rect 49870 58210 49922 58222
rect 49870 58146 49922 58158
rect 50206 58210 50258 58222
rect 50206 58146 50258 58158
rect 51662 58210 51714 58222
rect 51662 58146 51714 58158
rect 53230 58210 53282 58222
rect 53230 58146 53282 58158
rect 54462 58210 54514 58222
rect 54462 58146 54514 58158
rect 1344 58042 62608 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 62608 58042
rect 1344 57956 62608 57990
rect 14030 57874 14082 57886
rect 14030 57810 14082 57822
rect 14478 57874 14530 57886
rect 14478 57810 14530 57822
rect 14590 57874 14642 57886
rect 14590 57810 14642 57822
rect 24558 57874 24610 57886
rect 24558 57810 24610 57822
rect 24670 57874 24722 57886
rect 24670 57810 24722 57822
rect 40014 57874 40066 57886
rect 40014 57810 40066 57822
rect 42254 57874 42306 57886
rect 42254 57810 42306 57822
rect 43710 57874 43762 57886
rect 43710 57810 43762 57822
rect 47518 57874 47570 57886
rect 47518 57810 47570 57822
rect 48190 57874 48242 57886
rect 48190 57810 48242 57822
rect 49198 57874 49250 57886
rect 49198 57810 49250 57822
rect 14702 57762 14754 57774
rect 19406 57762 19458 57774
rect 15698 57710 15710 57762
rect 15762 57710 15774 57762
rect 16146 57710 16158 57762
rect 16210 57710 16222 57762
rect 14702 57698 14754 57710
rect 19406 57698 19458 57710
rect 24334 57762 24386 57774
rect 24334 57698 24386 57710
rect 24446 57762 24498 57774
rect 35198 57762 35250 57774
rect 33618 57710 33630 57762
rect 33682 57710 33694 57762
rect 24446 57698 24498 57710
rect 35198 57698 35250 57710
rect 36430 57762 36482 57774
rect 51886 57762 51938 57774
rect 44706 57710 44718 57762
rect 44770 57710 44782 57762
rect 49746 57710 49758 57762
rect 49810 57710 49822 57762
rect 36430 57698 36482 57710
rect 51886 57698 51938 57710
rect 52110 57762 52162 57774
rect 52110 57698 52162 57710
rect 56814 57762 56866 57774
rect 56814 57698 56866 57710
rect 14366 57650 14418 57662
rect 16382 57650 16434 57662
rect 19630 57650 19682 57662
rect 21870 57650 21922 57662
rect 25678 57650 25730 57662
rect 15026 57598 15038 57650
rect 15090 57598 15102 57650
rect 18834 57598 18846 57650
rect 18898 57598 18910 57650
rect 19170 57598 19182 57650
rect 19234 57598 19246 57650
rect 19954 57598 19966 57650
rect 20018 57598 20030 57650
rect 21186 57598 21198 57650
rect 21250 57598 21262 57650
rect 22082 57598 22094 57650
rect 22146 57598 22158 57650
rect 23874 57598 23886 57650
rect 23938 57598 23950 57650
rect 14366 57586 14418 57598
rect 16382 57586 16434 57598
rect 19630 57586 19682 57598
rect 21870 57586 21922 57598
rect 25678 57586 25730 57598
rect 26014 57650 26066 57662
rect 29598 57650 29650 57662
rect 34302 57650 34354 57662
rect 28130 57598 28142 57650
rect 28194 57598 28206 57650
rect 29250 57598 29262 57650
rect 29314 57598 29326 57650
rect 30146 57598 30158 57650
rect 30210 57598 30222 57650
rect 31154 57598 31166 57650
rect 31218 57598 31230 57650
rect 32386 57598 32398 57650
rect 32450 57598 32462 57650
rect 33730 57598 33742 57650
rect 33794 57598 33806 57650
rect 26014 57586 26066 57598
rect 29598 57586 29650 57598
rect 34302 57586 34354 57598
rect 35534 57650 35586 57662
rect 52558 57650 52610 57662
rect 47954 57598 47966 57650
rect 48018 57598 48030 57650
rect 49970 57598 49982 57650
rect 50034 57598 50046 57650
rect 51426 57598 51438 57650
rect 51490 57598 51502 57650
rect 52322 57598 52334 57650
rect 52386 57598 52398 57650
rect 35534 57586 35586 57598
rect 52558 57586 52610 57598
rect 52894 57650 52946 57662
rect 52894 57586 52946 57598
rect 53118 57650 53170 57662
rect 53118 57586 53170 57598
rect 53566 57650 53618 57662
rect 53566 57586 53618 57598
rect 53790 57650 53842 57662
rect 53790 57586 53842 57598
rect 54014 57650 54066 57662
rect 55794 57598 55806 57650
rect 55858 57598 55870 57650
rect 54014 57586 54066 57598
rect 12686 57538 12738 57550
rect 12686 57474 12738 57486
rect 13134 57538 13186 57550
rect 18174 57538 18226 57550
rect 26126 57538 26178 57550
rect 29822 57538 29874 57550
rect 36094 57538 36146 57550
rect 13570 57486 13582 57538
rect 13634 57486 13646 57538
rect 19282 57486 19294 57538
rect 19346 57486 19358 57538
rect 28466 57486 28478 57538
rect 28530 57486 28542 57538
rect 31714 57486 31726 57538
rect 31778 57486 31790 57538
rect 13134 57474 13186 57486
rect 18174 57474 18226 57486
rect 26126 57474 26178 57486
rect 29822 57474 29874 57486
rect 36094 57474 36146 57486
rect 36878 57538 36930 57550
rect 36878 57474 36930 57486
rect 37326 57538 37378 57550
rect 37326 57474 37378 57486
rect 37774 57538 37826 57550
rect 37774 57474 37826 57486
rect 41246 57538 41298 57550
rect 41246 57474 41298 57486
rect 41806 57538 41858 57550
rect 41806 57474 41858 57486
rect 46510 57538 46562 57550
rect 46510 57474 46562 57486
rect 47070 57538 47122 57550
rect 47070 57474 47122 57486
rect 50654 57538 50706 57550
rect 50654 57474 50706 57486
rect 50990 57538 51042 57550
rect 50990 57474 51042 57486
rect 52782 57538 52834 57550
rect 52782 57474 52834 57486
rect 53678 57538 53730 57550
rect 53678 57474 53730 57486
rect 55022 57538 55074 57550
rect 55458 57486 55470 57538
rect 55522 57486 55534 57538
rect 55022 57474 55074 57486
rect 16718 57426 16770 57438
rect 17950 57426 18002 57438
rect 34638 57426 34690 57438
rect 17602 57374 17614 57426
rect 17666 57374 17678 57426
rect 23202 57374 23214 57426
rect 23266 57374 23278 57426
rect 16718 57362 16770 57374
rect 17950 57362 18002 57374
rect 34638 57362 34690 57374
rect 45838 57426 45890 57438
rect 51774 57426 51826 57438
rect 46162 57374 46174 57426
rect 46226 57423 46238 57426
rect 46722 57423 46734 57426
rect 46226 57377 46734 57423
rect 46226 57374 46238 57377
rect 46722 57374 46734 57377
rect 46786 57374 46798 57426
rect 45838 57362 45890 57374
rect 51774 57362 51826 57374
rect 54462 57426 54514 57438
rect 54462 57362 54514 57374
rect 54798 57426 54850 57438
rect 54798 57362 54850 57374
rect 1344 57258 62608 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 62608 57258
rect 1344 57172 62608 57206
rect 15262 57090 15314 57102
rect 17166 57090 17218 57102
rect 32174 57090 32226 57102
rect 15586 57038 15598 57090
rect 15650 57038 15662 57090
rect 25666 57038 25678 57090
rect 25730 57038 25742 57090
rect 15262 57026 15314 57038
rect 17166 57026 17218 57038
rect 32174 57026 32226 57038
rect 32510 57090 32562 57102
rect 51438 57090 51490 57102
rect 37202 57038 37214 57090
rect 37266 57087 37278 57090
rect 38546 57087 38558 57090
rect 37266 57041 38558 57087
rect 37266 57038 37278 57041
rect 38546 57038 38558 57041
rect 38610 57038 38622 57090
rect 32510 57026 32562 57038
rect 51438 57026 51490 57038
rect 55022 57090 55074 57102
rect 55022 57026 55074 57038
rect 12126 56978 12178 56990
rect 12126 56914 12178 56926
rect 14030 56978 14082 56990
rect 14030 56914 14082 56926
rect 15038 56978 15090 56990
rect 21310 56978 21362 56990
rect 31166 56978 31218 56990
rect 19394 56926 19406 56978
rect 19458 56926 19470 56978
rect 26450 56926 26462 56978
rect 26514 56926 26526 56978
rect 15038 56914 15090 56926
rect 21310 56914 21362 56926
rect 31166 56914 31218 56926
rect 32734 56978 32786 56990
rect 38558 56978 38610 56990
rect 33394 56926 33406 56978
rect 33458 56926 33470 56978
rect 32734 56914 32786 56926
rect 38558 56914 38610 56926
rect 39566 56978 39618 56990
rect 44942 56978 44994 56990
rect 41346 56926 41358 56978
rect 41410 56926 41422 56978
rect 42690 56926 42702 56978
rect 42754 56926 42766 56978
rect 39566 56914 39618 56926
rect 44942 56914 44994 56926
rect 56366 56978 56418 56990
rect 56366 56914 56418 56926
rect 57822 56978 57874 56990
rect 57822 56914 57874 56926
rect 13022 56866 13074 56878
rect 13022 56802 13074 56814
rect 13582 56866 13634 56878
rect 16830 56866 16882 56878
rect 16034 56814 16046 56866
rect 16098 56814 16110 56866
rect 13582 56802 13634 56814
rect 16830 56802 16882 56814
rect 18510 56866 18562 56878
rect 20750 56866 20802 56878
rect 22766 56866 22818 56878
rect 40686 56866 40738 56878
rect 19506 56814 19518 56866
rect 19570 56814 19582 56866
rect 20514 56814 20526 56866
rect 20578 56814 20590 56866
rect 22082 56814 22094 56866
rect 22146 56814 22158 56866
rect 24098 56814 24110 56866
rect 24162 56814 24174 56866
rect 26674 56814 26686 56866
rect 26738 56814 26750 56866
rect 27570 56814 27582 56866
rect 27634 56814 27646 56866
rect 29586 56814 29598 56866
rect 29650 56814 29662 56866
rect 30370 56814 30382 56866
rect 30434 56814 30446 56866
rect 30594 56814 30606 56866
rect 30658 56814 30670 56866
rect 18510 56802 18562 56814
rect 20750 56802 20802 56814
rect 22766 56802 22818 56814
rect 40686 56802 40738 56814
rect 40910 56866 40962 56878
rect 55694 56866 55746 56878
rect 41458 56814 41470 56866
rect 41522 56814 41534 56866
rect 42578 56814 42590 56866
rect 42642 56814 42654 56866
rect 57250 56814 57262 56866
rect 57314 56814 57326 56866
rect 40910 56802 40962 56814
rect 55694 56802 55746 56814
rect 14366 56754 14418 56766
rect 14366 56690 14418 56702
rect 14702 56754 14754 56766
rect 17614 56754 17666 56766
rect 16258 56702 16270 56754
rect 16322 56702 16334 56754
rect 14702 56690 14754 56702
rect 17614 56690 17666 56702
rect 18174 56754 18226 56766
rect 18174 56690 18226 56702
rect 18734 56754 18786 56766
rect 18734 56690 18786 56702
rect 19742 56754 19794 56766
rect 19742 56690 19794 56702
rect 21422 56754 21474 56766
rect 24558 56754 24610 56766
rect 31278 56754 31330 56766
rect 21970 56702 21982 56754
rect 22034 56702 22046 56754
rect 23986 56702 23998 56754
rect 24050 56702 24062 56754
rect 28018 56702 28030 56754
rect 28082 56702 28094 56754
rect 29250 56702 29262 56754
rect 29314 56702 29326 56754
rect 29922 56702 29934 56754
rect 29986 56702 29998 56754
rect 21422 56690 21474 56702
rect 24558 56690 24610 56702
rect 31278 56690 31330 56702
rect 31390 56754 31442 56766
rect 33070 56754 33122 56766
rect 31490 56702 31502 56754
rect 31554 56702 31566 56754
rect 31390 56690 31442 56702
rect 33070 56690 33122 56702
rect 33742 56754 33794 56766
rect 37102 56754 37154 56766
rect 35074 56702 35086 56754
rect 35138 56702 35150 56754
rect 33742 56690 33794 56702
rect 37102 56690 37154 56702
rect 40462 56754 40514 56766
rect 40462 56690 40514 56702
rect 42254 56754 42306 56766
rect 42254 56690 42306 56702
rect 45838 56754 45890 56766
rect 55470 56754 55522 56766
rect 46498 56702 46510 56754
rect 46562 56702 46574 56754
rect 47618 56702 47630 56754
rect 47682 56702 47694 56754
rect 53778 56702 53790 56754
rect 53842 56702 53854 56754
rect 45838 56690 45890 56702
rect 55470 56690 55522 56702
rect 57038 56754 57090 56766
rect 57038 56690 57090 56702
rect 58270 56754 58322 56766
rect 58270 56690 58322 56702
rect 11678 56642 11730 56654
rect 11678 56578 11730 56590
rect 12574 56642 12626 56654
rect 12574 56578 12626 56590
rect 17726 56642 17778 56654
rect 17726 56578 17778 56590
rect 17950 56642 18002 56654
rect 17950 56578 18002 56590
rect 18286 56642 18338 56654
rect 18286 56578 18338 56590
rect 23102 56642 23154 56654
rect 23102 56578 23154 56590
rect 24334 56642 24386 56654
rect 24334 56578 24386 56590
rect 24446 56642 24498 56654
rect 24446 56578 24498 56590
rect 31054 56642 31106 56654
rect 31054 56578 31106 56590
rect 33294 56642 33346 56654
rect 33294 56578 33346 56590
rect 33854 56642 33906 56654
rect 33854 56578 33906 56590
rect 33966 56642 34018 56654
rect 33966 56578 34018 56590
rect 36206 56642 36258 56654
rect 36206 56578 36258 56590
rect 37662 56642 37714 56654
rect 37662 56578 37714 56590
rect 37998 56642 38050 56654
rect 37998 56578 38050 56590
rect 38894 56642 38946 56654
rect 38894 56578 38946 56590
rect 40126 56642 40178 56654
rect 40126 56578 40178 56590
rect 40798 56642 40850 56654
rect 40798 56578 40850 56590
rect 43486 56642 43538 56654
rect 43486 56578 43538 56590
rect 44046 56642 44098 56654
rect 44046 56578 44098 56590
rect 45502 56642 45554 56654
rect 45502 56578 45554 56590
rect 46174 56642 46226 56654
rect 46174 56578 46226 56590
rect 48974 56642 49026 56654
rect 52222 56642 52274 56654
rect 50082 56590 50094 56642
rect 50146 56590 50158 56642
rect 48974 56578 49026 56590
rect 52222 56578 52274 56590
rect 52894 56642 52946 56654
rect 56478 56642 56530 56654
rect 56018 56590 56030 56642
rect 56082 56590 56094 56642
rect 52894 56578 52946 56590
rect 56478 56578 56530 56590
rect 1344 56474 62608 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 62608 56474
rect 1344 56388 62608 56422
rect 15598 56306 15650 56318
rect 30382 56306 30434 56318
rect 32062 56306 32114 56318
rect 21186 56254 21198 56306
rect 21250 56254 21262 56306
rect 23650 56254 23662 56306
rect 23714 56254 23726 56306
rect 31378 56254 31390 56306
rect 31442 56254 31454 56306
rect 15598 56242 15650 56254
rect 30382 56242 30434 56254
rect 32062 56242 32114 56254
rect 32398 56306 32450 56318
rect 32398 56242 32450 56254
rect 38446 56306 38498 56318
rect 38446 56242 38498 56254
rect 38558 56306 38610 56318
rect 38558 56242 38610 56254
rect 46734 56306 46786 56318
rect 46734 56242 46786 56254
rect 48078 56306 48130 56318
rect 48078 56242 48130 56254
rect 48862 56306 48914 56318
rect 55358 56306 55410 56318
rect 51650 56254 51662 56306
rect 51714 56254 51726 56306
rect 48862 56242 48914 56254
rect 55358 56242 55410 56254
rect 58382 56306 58434 56318
rect 58382 56242 58434 56254
rect 59278 56306 59330 56318
rect 59278 56242 59330 56254
rect 22990 56194 23042 56206
rect 25566 56194 25618 56206
rect 16146 56142 16158 56194
rect 16210 56142 16222 56194
rect 16594 56142 16606 56194
rect 16658 56142 16670 56194
rect 21858 56142 21870 56194
rect 21922 56142 21934 56194
rect 23538 56142 23550 56194
rect 23602 56142 23614 56194
rect 24322 56142 24334 56194
rect 24386 56142 24398 56194
rect 22990 56130 23042 56142
rect 25566 56130 25618 56142
rect 27022 56194 27074 56206
rect 27022 56130 27074 56142
rect 27470 56194 27522 56206
rect 29150 56194 29202 56206
rect 28130 56142 28142 56194
rect 28194 56142 28206 56194
rect 28802 56142 28814 56194
rect 28866 56142 28878 56194
rect 27470 56130 27522 56142
rect 29150 56130 29202 56142
rect 30494 56194 30546 56206
rect 30494 56130 30546 56142
rect 31614 56194 31666 56206
rect 31614 56130 31666 56142
rect 32174 56194 32226 56206
rect 55582 56194 55634 56206
rect 34626 56142 34638 56194
rect 34690 56142 34702 56194
rect 42914 56142 42926 56194
rect 42978 56142 42990 56194
rect 45266 56142 45278 56194
rect 45330 56142 45342 56194
rect 45602 56142 45614 56194
rect 45666 56142 45678 56194
rect 47058 56142 47070 56194
rect 47122 56142 47134 56194
rect 49858 56142 49870 56194
rect 49922 56142 49934 56194
rect 57810 56142 57822 56194
rect 57874 56142 57886 56194
rect 32174 56130 32226 56142
rect 55582 56130 55634 56142
rect 15934 56082 15986 56094
rect 20190 56082 20242 56094
rect 22430 56082 22482 56094
rect 23438 56082 23490 56094
rect 25790 56082 25842 56094
rect 15026 56030 15038 56082
rect 15090 56030 15102 56082
rect 17490 56030 17502 56082
rect 17554 56030 17566 56082
rect 18498 56030 18510 56082
rect 18562 56030 18574 56082
rect 19730 56030 19742 56082
rect 19794 56030 19806 56082
rect 20626 56030 20638 56082
rect 20690 56030 20702 56082
rect 21074 56030 21086 56082
rect 21138 56030 21150 56082
rect 22082 56030 22094 56082
rect 22146 56030 22158 56082
rect 22754 56030 22766 56082
rect 22818 56030 22830 56082
rect 25218 56030 25230 56082
rect 25282 56030 25294 56082
rect 15934 56018 15986 56030
rect 20190 56018 20242 56030
rect 22430 56018 22482 56030
rect 23438 56018 23490 56030
rect 25790 56018 25842 56030
rect 25902 56082 25954 56094
rect 25902 56018 25954 56030
rect 27582 56082 27634 56094
rect 29374 56082 29426 56094
rect 27906 56030 27918 56082
rect 27970 56030 27982 56082
rect 27582 56018 27634 56030
rect 29374 56018 29426 56030
rect 29598 56082 29650 56094
rect 31278 56082 31330 56094
rect 29922 56030 29934 56082
rect 29986 56030 29998 56082
rect 30818 56030 30830 56082
rect 30882 56030 30894 56082
rect 29598 56018 29650 56030
rect 31278 56018 31330 56030
rect 31950 56082 32002 56094
rect 31950 56018 32002 56030
rect 33182 56082 33234 56094
rect 33182 56018 33234 56030
rect 33630 56082 33682 56094
rect 33630 56018 33682 56030
rect 33854 56082 33906 56094
rect 37102 56082 37154 56094
rect 35410 56030 35422 56082
rect 35474 56030 35486 56082
rect 36194 56030 36206 56082
rect 36258 56030 36270 56082
rect 33854 56018 33906 56030
rect 37102 56018 37154 56030
rect 37886 56082 37938 56094
rect 37886 56018 37938 56030
rect 38334 56082 38386 56094
rect 38334 56018 38386 56030
rect 45950 56082 46002 56094
rect 50542 56082 50594 56094
rect 57038 56082 57090 56094
rect 48178 56030 48190 56082
rect 48242 56030 48254 56082
rect 49746 56030 49758 56082
rect 49810 56030 49822 56082
rect 54898 56030 54910 56082
rect 54962 56030 54974 56082
rect 55122 56030 55134 56082
rect 55186 56030 55198 56082
rect 57698 56030 57710 56082
rect 57762 56030 57774 56082
rect 58258 56030 58270 56082
rect 58322 56030 58334 56082
rect 45950 56018 46002 56030
rect 50542 56018 50594 56030
rect 57038 56018 57090 56030
rect 11230 55970 11282 55982
rect 11230 55906 11282 55918
rect 11678 55970 11730 55982
rect 11678 55906 11730 55918
rect 12126 55970 12178 55982
rect 12126 55906 12178 55918
rect 12574 55970 12626 55982
rect 12574 55906 12626 55918
rect 13022 55970 13074 55982
rect 13022 55906 13074 55918
rect 13470 55970 13522 55982
rect 13470 55906 13522 55918
rect 13806 55970 13858 55982
rect 13806 55906 13858 55918
rect 14366 55970 14418 55982
rect 37662 55970 37714 55982
rect 14690 55918 14702 55970
rect 14754 55918 14766 55970
rect 18162 55918 18174 55970
rect 18226 55918 18238 55970
rect 33394 55918 33406 55970
rect 33458 55918 33470 55970
rect 34626 55918 34638 55970
rect 34690 55918 34702 55970
rect 14366 55906 14418 55918
rect 37662 55906 37714 55918
rect 39006 55970 39058 55982
rect 39006 55906 39058 55918
rect 39454 55970 39506 55982
rect 39454 55906 39506 55918
rect 40126 55970 40178 55982
rect 40126 55906 40178 55918
rect 41022 55970 41074 55982
rect 41022 55906 41074 55918
rect 41470 55970 41522 55982
rect 41470 55906 41522 55918
rect 42254 55970 42306 55982
rect 42254 55906 42306 55918
rect 47630 55970 47682 55982
rect 47630 55906 47682 55918
rect 54238 55970 54290 55982
rect 56142 55970 56194 55982
rect 55346 55918 55358 55970
rect 55410 55918 55422 55970
rect 54238 55906 54290 55918
rect 56142 55906 56194 55918
rect 23102 55858 23154 55870
rect 13010 55806 13022 55858
rect 13074 55855 13086 55858
rect 14354 55855 14366 55858
rect 13074 55809 14366 55855
rect 13074 55806 13086 55809
rect 14354 55806 14366 55809
rect 14418 55806 14430 55858
rect 23102 55794 23154 55806
rect 27470 55858 27522 55870
rect 27470 55794 27522 55806
rect 30382 55858 30434 55870
rect 30382 55794 30434 55806
rect 31166 55858 31218 55870
rect 31166 55794 31218 55806
rect 33070 55858 33122 55870
rect 33070 55794 33122 55806
rect 44830 55858 44882 55870
rect 44830 55794 44882 55806
rect 46286 55858 46338 55870
rect 46286 55794 46338 55806
rect 49198 55858 49250 55870
rect 49198 55794 49250 55806
rect 50430 55858 50482 55870
rect 56702 55858 56754 55870
rect 53106 55806 53118 55858
rect 53170 55806 53182 55858
rect 50430 55794 50482 55806
rect 56702 55794 56754 55806
rect 1344 55690 62608 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 62608 55690
rect 1344 55604 62608 55638
rect 20638 55522 20690 55534
rect 20638 55458 20690 55470
rect 31054 55522 31106 55534
rect 31054 55458 31106 55470
rect 35310 55522 35362 55534
rect 41010 55470 41022 55522
rect 41074 55470 41086 55522
rect 55794 55470 55806 55522
rect 55858 55470 55870 55522
rect 35310 55458 35362 55470
rect 15486 55410 15538 55422
rect 15486 55346 15538 55358
rect 18398 55410 18450 55422
rect 25342 55410 25394 55422
rect 23762 55358 23774 55410
rect 23826 55358 23838 55410
rect 18398 55346 18450 55358
rect 25342 55346 25394 55358
rect 29598 55410 29650 55422
rect 29598 55346 29650 55358
rect 30158 55410 30210 55422
rect 30158 55346 30210 55358
rect 32734 55410 32786 55422
rect 46174 55410 46226 55422
rect 38882 55358 38894 55410
rect 38946 55358 38958 55410
rect 42914 55358 42926 55410
rect 42978 55358 42990 55410
rect 32734 55346 32786 55358
rect 46174 55346 46226 55358
rect 47742 55410 47794 55422
rect 47742 55346 47794 55358
rect 25230 55298 25282 55310
rect 23426 55246 23438 55298
rect 23490 55246 23502 55298
rect 24210 55246 24222 55298
rect 24274 55246 24286 55298
rect 24770 55246 24782 55298
rect 24834 55246 24846 55298
rect 25230 55234 25282 55246
rect 25678 55298 25730 55310
rect 25678 55234 25730 55246
rect 26574 55298 26626 55310
rect 26574 55234 26626 55246
rect 27134 55298 27186 55310
rect 29262 55298 29314 55310
rect 27682 55246 27694 55298
rect 27746 55246 27758 55298
rect 28466 55246 28478 55298
rect 28530 55246 28542 55298
rect 27134 55234 27186 55246
rect 29262 55234 29314 55246
rect 29486 55298 29538 55310
rect 29486 55234 29538 55246
rect 29822 55298 29874 55310
rect 29822 55234 29874 55246
rect 30046 55298 30098 55310
rect 30046 55234 30098 55246
rect 30718 55298 30770 55310
rect 30718 55234 30770 55246
rect 31390 55298 31442 55310
rect 32622 55298 32674 55310
rect 36990 55298 37042 55310
rect 39678 55298 39730 55310
rect 42590 55298 42642 55310
rect 47966 55298 48018 55310
rect 52670 55298 52722 55310
rect 32162 55246 32174 55298
rect 32226 55246 32238 55298
rect 35634 55246 35646 55298
rect 35698 55246 35710 55298
rect 38994 55246 39006 55298
rect 39058 55246 39070 55298
rect 40562 55246 40574 55298
rect 40626 55246 40638 55298
rect 43362 55246 43374 55298
rect 43426 55246 43438 55298
rect 45714 55246 45726 55298
rect 45778 55246 45790 55298
rect 48738 55246 48750 55298
rect 48802 55246 48814 55298
rect 49298 55246 49310 55298
rect 49362 55246 49374 55298
rect 50306 55246 50318 55298
rect 50370 55246 50382 55298
rect 31390 55234 31442 55246
rect 32622 55234 32674 55246
rect 36990 55234 37042 55246
rect 39678 55234 39730 55246
rect 42590 55234 42642 55246
rect 47966 55234 48018 55246
rect 52670 55234 52722 55246
rect 53230 55298 53282 55310
rect 53230 55234 53282 55246
rect 53902 55298 53954 55310
rect 55570 55246 55582 55298
rect 55634 55246 55646 55298
rect 56690 55246 56702 55298
rect 56754 55246 56766 55298
rect 58146 55246 58158 55298
rect 58210 55246 58222 55298
rect 53902 55234 53954 55246
rect 1710 55186 1762 55198
rect 25566 55186 25618 55198
rect 14130 55134 14142 55186
rect 14194 55134 14206 55186
rect 16482 55134 16494 55186
rect 16546 55134 16558 55186
rect 19170 55134 19182 55186
rect 19234 55134 19246 55186
rect 1710 55122 1762 55134
rect 25566 55122 25618 55134
rect 26686 55186 26738 55198
rect 30270 55186 30322 55198
rect 42814 55186 42866 55198
rect 27794 55134 27806 55186
rect 27858 55134 27870 55186
rect 31938 55134 31950 55186
rect 32002 55134 32014 55186
rect 33394 55134 33406 55186
rect 33458 55134 33470 55186
rect 37314 55134 37326 55186
rect 37378 55134 37390 55186
rect 26686 55122 26738 55134
rect 30270 55122 30322 55134
rect 42814 55122 42866 55134
rect 42926 55186 42978 55198
rect 46510 55186 46562 55198
rect 54126 55186 54178 55198
rect 58718 55186 58770 55198
rect 45490 55134 45502 55186
rect 45554 55134 45566 55186
rect 48402 55134 48414 55186
rect 48466 55134 48478 55186
rect 55458 55134 55470 55186
rect 55522 55134 55534 55186
rect 42926 55122 42978 55134
rect 46510 55122 46562 55134
rect 54126 55122 54178 55134
rect 58718 55122 58770 55134
rect 58942 55186 58994 55198
rect 58942 55122 58994 55134
rect 59278 55186 59330 55198
rect 59278 55122 59330 55134
rect 59614 55186 59666 55198
rect 59614 55122 59666 55134
rect 61070 55186 61122 55198
rect 61070 55122 61122 55134
rect 2046 55074 2098 55086
rect 2046 55010 2098 55022
rect 2494 55074 2546 55086
rect 2494 55010 2546 55022
rect 9998 55074 10050 55086
rect 9998 55010 10050 55022
rect 10558 55074 10610 55086
rect 10558 55010 10610 55022
rect 11006 55074 11058 55086
rect 11006 55010 11058 55022
rect 11454 55074 11506 55086
rect 11454 55010 11506 55022
rect 11902 55074 11954 55086
rect 11902 55010 11954 55022
rect 12350 55074 12402 55086
rect 12350 55010 12402 55022
rect 13022 55074 13074 55086
rect 23102 55074 23154 55086
rect 21970 55022 21982 55074
rect 22034 55022 22046 55074
rect 13022 55010 13074 55022
rect 23102 55010 23154 55022
rect 26910 55074 26962 55086
rect 35870 55074 35922 55086
rect 28242 55022 28254 55074
rect 28306 55022 28318 55074
rect 26910 55010 26962 55022
rect 35870 55010 35922 55022
rect 36318 55074 36370 55086
rect 36318 55010 36370 55022
rect 41918 55074 41970 55086
rect 41918 55010 41970 55022
rect 42254 55074 42306 55086
rect 42254 55010 42306 55022
rect 43934 55074 43986 55086
rect 43934 55010 43986 55022
rect 44270 55074 44322 55086
rect 44270 55010 44322 55022
rect 44942 55074 44994 55086
rect 44942 55010 44994 55022
rect 47182 55074 47234 55086
rect 51214 55074 51266 55086
rect 47394 55022 47406 55074
rect 47458 55022 47470 55074
rect 47182 55010 47234 55022
rect 51214 55010 51266 55022
rect 51662 55074 51714 55086
rect 51662 55010 51714 55022
rect 51886 55074 51938 55086
rect 51886 55010 51938 55022
rect 51998 55074 52050 55086
rect 51998 55010 52050 55022
rect 52110 55074 52162 55086
rect 58382 55074 58434 55086
rect 53554 55022 53566 55074
rect 53618 55022 53630 55074
rect 52110 55010 52162 55022
rect 58382 55010 58434 55022
rect 58494 55074 58546 55086
rect 58494 55010 58546 55022
rect 60734 55074 60786 55086
rect 60734 55010 60786 55022
rect 1344 54906 62608 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 62608 54906
rect 1344 54820 62608 54854
rect 12686 54738 12738 54750
rect 12686 54674 12738 54686
rect 13246 54738 13298 54750
rect 15038 54738 15090 54750
rect 14578 54686 14590 54738
rect 14642 54686 14654 54738
rect 13246 54674 13298 54686
rect 15038 54674 15090 54686
rect 20862 54738 20914 54750
rect 20862 54674 20914 54686
rect 29486 54738 29538 54750
rect 39342 54738 39394 54750
rect 36306 54686 36318 54738
rect 36370 54686 36382 54738
rect 37762 54686 37774 54738
rect 37826 54686 37838 54738
rect 29486 54674 29538 54686
rect 39342 54674 39394 54686
rect 44718 54738 44770 54750
rect 44718 54674 44770 54686
rect 47070 54738 47122 54750
rect 48738 54686 48750 54738
rect 48802 54686 48814 54738
rect 59378 54686 59390 54738
rect 59442 54686 59454 54738
rect 47070 54674 47122 54686
rect 13806 54626 13858 54638
rect 16718 54626 16770 54638
rect 15922 54574 15934 54626
rect 15986 54574 15998 54626
rect 13806 54562 13858 54574
rect 16718 54562 16770 54574
rect 17390 54626 17442 54638
rect 18510 54626 18562 54638
rect 20974 54626 21026 54638
rect 21870 54626 21922 54638
rect 23886 54626 23938 54638
rect 17602 54574 17614 54626
rect 17666 54574 17678 54626
rect 20290 54574 20302 54626
rect 20354 54574 20366 54626
rect 21522 54574 21534 54626
rect 21586 54574 21598 54626
rect 22530 54574 22542 54626
rect 22594 54574 22606 54626
rect 17390 54562 17442 54574
rect 18510 54562 18562 54574
rect 20974 54562 21026 54574
rect 21870 54562 21922 54574
rect 23886 54562 23938 54574
rect 24558 54626 24610 54638
rect 24558 54562 24610 54574
rect 28478 54626 28530 54638
rect 32174 54626 32226 54638
rect 30930 54574 30942 54626
rect 30994 54574 31006 54626
rect 31378 54574 31390 54626
rect 31442 54574 31454 54626
rect 28478 54562 28530 54574
rect 32174 54562 32226 54574
rect 32510 54626 32562 54638
rect 32510 54562 32562 54574
rect 37214 54626 37266 54638
rect 37214 54562 37266 54574
rect 38446 54626 38498 54638
rect 47406 54626 47458 54638
rect 45602 54574 45614 54626
rect 45666 54574 45678 54626
rect 38446 54562 38498 54574
rect 47406 54562 47458 54574
rect 47630 54626 47682 54638
rect 49858 54574 49870 54626
rect 49922 54574 49934 54626
rect 52098 54574 52110 54626
rect 52162 54574 52174 54626
rect 52770 54574 52782 54626
rect 52834 54574 52846 54626
rect 53218 54574 53230 54626
rect 53282 54574 53294 54626
rect 55906 54574 55918 54626
rect 55970 54574 55982 54626
rect 47630 54562 47682 54574
rect 12462 54514 12514 54526
rect 12462 54450 12514 54462
rect 12798 54514 12850 54526
rect 12798 54450 12850 54462
rect 13134 54514 13186 54526
rect 13134 54450 13186 54462
rect 13694 54514 13746 54526
rect 13694 54450 13746 54462
rect 14254 54514 14306 54526
rect 14254 54450 14306 54462
rect 15374 54514 15426 54526
rect 16830 54514 16882 54526
rect 18622 54514 18674 54526
rect 22094 54514 22146 54526
rect 24334 54514 24386 54526
rect 29262 54514 29314 54526
rect 16146 54462 16158 54514
rect 16210 54462 16222 54514
rect 17938 54462 17950 54514
rect 18002 54462 18014 54514
rect 18946 54462 18958 54514
rect 19010 54462 19022 54514
rect 19506 54462 19518 54514
rect 19570 54462 19582 54514
rect 20178 54462 20190 54514
rect 20242 54462 20254 54514
rect 21634 54462 21646 54514
rect 21698 54462 21710 54514
rect 23426 54462 23438 54514
rect 23490 54462 23502 54514
rect 28018 54462 28030 54514
rect 28082 54462 28094 54514
rect 28690 54462 28702 54514
rect 28754 54462 28766 54514
rect 15374 54450 15426 54462
rect 16830 54450 16882 54462
rect 18622 54450 18674 54462
rect 22094 54450 22146 54462
rect 24334 54450 24386 54462
rect 29262 54450 29314 54462
rect 29486 54514 29538 54526
rect 29486 54450 29538 54462
rect 29710 54514 29762 54526
rect 36654 54514 36706 54526
rect 30146 54462 30158 54514
rect 30210 54462 30222 54514
rect 30594 54462 30606 54514
rect 30658 54462 30670 54514
rect 31266 54462 31278 54514
rect 31330 54462 31342 54514
rect 33170 54462 33182 54514
rect 33234 54462 33246 54514
rect 29710 54450 29762 54462
rect 36654 54450 36706 54462
rect 36878 54514 36930 54526
rect 36878 54450 36930 54462
rect 37438 54514 37490 54526
rect 37438 54450 37490 54462
rect 38110 54514 38162 54526
rect 45054 54514 45106 54526
rect 46286 54514 46338 54526
rect 41346 54462 41358 54514
rect 41410 54462 41422 54514
rect 45714 54462 45726 54514
rect 45778 54462 45790 54514
rect 38110 54450 38162 54462
rect 45054 54450 45106 54462
rect 46286 54450 46338 54462
rect 46622 54514 46674 54526
rect 53454 54514 53506 54526
rect 46946 54462 46958 54514
rect 47010 54462 47022 54514
rect 50418 54462 50430 54514
rect 50482 54462 50494 54514
rect 51650 54462 51662 54514
rect 51714 54462 51726 54514
rect 46622 54450 46674 54462
rect 53454 54450 53506 54462
rect 53790 54514 53842 54526
rect 53790 54450 53842 54462
rect 54462 54514 54514 54526
rect 54462 54450 54514 54462
rect 54686 54514 54738 54526
rect 56578 54462 56590 54514
rect 56642 54462 56654 54514
rect 54686 54450 54738 54462
rect 9662 54402 9714 54414
rect 9662 54338 9714 54350
rect 10222 54402 10274 54414
rect 10222 54338 10274 54350
rect 10670 54402 10722 54414
rect 10670 54338 10722 54350
rect 11006 54402 11058 54414
rect 11006 54338 11058 54350
rect 11790 54402 11842 54414
rect 11790 54338 11842 54350
rect 12126 54402 12178 54414
rect 12126 54338 12178 54350
rect 17502 54402 17554 54414
rect 17502 54338 17554 54350
rect 17838 54402 17890 54414
rect 17838 54338 17890 54350
rect 19854 54402 19906 54414
rect 38894 54402 38946 54414
rect 21298 54350 21310 54402
rect 21362 54350 21374 54402
rect 25218 54350 25230 54402
rect 25282 54350 25294 54402
rect 27346 54350 27358 54402
rect 27410 54350 27422 54402
rect 33842 54350 33854 54402
rect 33906 54350 33918 54402
rect 35970 54350 35982 54402
rect 36034 54350 36046 54402
rect 19854 54338 19906 54350
rect 38894 54338 38946 54350
rect 39790 54402 39842 54414
rect 39790 54338 39842 54350
rect 40238 54402 40290 54414
rect 40238 54338 40290 54350
rect 41134 54402 41186 54414
rect 47518 54402 47570 54414
rect 42130 54350 42142 54402
rect 42194 54350 42206 54402
rect 44258 54350 44270 54402
rect 44322 54350 44334 54402
rect 41134 54338 41186 54350
rect 47518 54338 47570 54350
rect 48190 54402 48242 54414
rect 48190 54338 48242 54350
rect 49310 54402 49362 54414
rect 60510 54402 60562 54414
rect 55682 54350 55694 54402
rect 55746 54350 55758 54402
rect 49310 54338 49362 54350
rect 60510 54338 60562 54350
rect 61070 54402 61122 54414
rect 61070 54338 61122 54350
rect 61518 54402 61570 54414
rect 61518 54338 61570 54350
rect 61854 54402 61906 54414
rect 61854 54338 61906 54350
rect 12238 54290 12290 54302
rect 12238 54226 12290 54238
rect 13246 54290 13298 54302
rect 13246 54226 13298 54238
rect 13806 54290 13858 54302
rect 13806 54226 13858 54238
rect 16718 54290 16770 54302
rect 24670 54290 24722 54302
rect 48078 54290 48130 54302
rect 22978 54238 22990 54290
rect 23042 54238 23054 54290
rect 38770 54238 38782 54290
rect 38834 54287 38846 54290
rect 39330 54287 39342 54290
rect 38834 54241 39342 54287
rect 38834 54238 38846 54241
rect 39330 54238 39342 54241
rect 39394 54238 39406 54290
rect 46834 54238 46846 54290
rect 46898 54238 46910 54290
rect 16718 54226 16770 54238
rect 24670 54226 24722 54238
rect 48078 54226 48130 54238
rect 49086 54290 49138 54302
rect 49086 54226 49138 54238
rect 54350 54290 54402 54302
rect 54350 54226 54402 54238
rect 56702 54290 56754 54302
rect 57922 54238 57934 54290
rect 57986 54238 57998 54290
rect 56702 54226 56754 54238
rect 1344 54122 62608 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 62608 54122
rect 1344 54036 62608 54070
rect 13806 53954 13858 53966
rect 27694 53954 27746 53966
rect 10658 53902 10670 53954
rect 10722 53951 10734 53954
rect 10722 53905 11727 53951
rect 10722 53902 10734 53905
rect 11681 53842 11727 53905
rect 16258 53902 16270 53954
rect 16322 53902 16334 53954
rect 23986 53902 23998 53954
rect 24050 53902 24062 53954
rect 13806 53890 13858 53902
rect 27694 53890 27746 53902
rect 30158 53954 30210 53966
rect 30158 53890 30210 53902
rect 30382 53954 30434 53966
rect 30382 53890 30434 53902
rect 30830 53954 30882 53966
rect 30830 53890 30882 53902
rect 31278 53954 31330 53966
rect 31278 53890 31330 53902
rect 44942 53954 44994 53966
rect 44942 53890 44994 53902
rect 52894 53954 52946 53966
rect 56914 53902 56926 53954
rect 56978 53902 56990 53954
rect 57698 53902 57710 53954
rect 57762 53902 57774 53954
rect 52894 53890 52946 53902
rect 18846 53842 18898 53854
rect 11666 53790 11678 53842
rect 11730 53790 11742 53842
rect 18846 53778 18898 53790
rect 20750 53842 20802 53854
rect 31502 53842 31554 53854
rect 21970 53790 21982 53842
rect 22034 53790 22046 53842
rect 22194 53790 22206 53842
rect 22258 53790 22270 53842
rect 25106 53790 25118 53842
rect 25170 53790 25182 53842
rect 20750 53778 20802 53790
rect 31502 53778 31554 53790
rect 31838 53842 31890 53854
rect 31838 53778 31890 53790
rect 45390 53842 45442 53854
rect 61294 53842 61346 53854
rect 51090 53790 51102 53842
rect 51154 53790 51166 53842
rect 58146 53790 58158 53842
rect 58210 53790 58222 53842
rect 45390 53778 45442 53790
rect 61294 53778 61346 53790
rect 10110 53730 10162 53742
rect 10110 53666 10162 53678
rect 10894 53730 10946 53742
rect 10894 53666 10946 53678
rect 12910 53730 12962 53742
rect 12910 53666 12962 53678
rect 13694 53730 13746 53742
rect 13694 53666 13746 53678
rect 14142 53730 14194 53742
rect 14142 53666 14194 53678
rect 14814 53730 14866 53742
rect 14814 53666 14866 53678
rect 15150 53730 15202 53742
rect 15150 53666 15202 53678
rect 15486 53730 15538 53742
rect 15486 53666 15538 53678
rect 15710 53730 15762 53742
rect 15710 53666 15762 53678
rect 16046 53730 16098 53742
rect 17278 53730 17330 53742
rect 16258 53678 16270 53730
rect 16322 53678 16334 53730
rect 16046 53666 16098 53678
rect 17278 53666 17330 53678
rect 18174 53730 18226 53742
rect 19070 53730 19122 53742
rect 25454 53730 25506 53742
rect 27246 53730 27298 53742
rect 30718 53730 30770 53742
rect 18722 53678 18734 53730
rect 18786 53678 18798 53730
rect 19842 53678 19854 53730
rect 19906 53678 19918 53730
rect 21522 53678 21534 53730
rect 21586 53678 21598 53730
rect 22306 53678 22318 53730
rect 22370 53678 22382 53730
rect 24770 53678 24782 53730
rect 24834 53678 24846 53730
rect 26674 53678 26686 53730
rect 26738 53678 26750 53730
rect 27458 53678 27470 53730
rect 27522 53678 27534 53730
rect 27906 53678 27918 53730
rect 27970 53678 27982 53730
rect 29250 53678 29262 53730
rect 29314 53678 29326 53730
rect 18174 53666 18226 53678
rect 19070 53666 19122 53678
rect 25454 53666 25506 53678
rect 27246 53666 27298 53678
rect 30718 53666 30770 53678
rect 31950 53730 32002 53742
rect 31950 53666 32002 53678
rect 36094 53730 36146 53742
rect 36094 53666 36146 53678
rect 36206 53730 36258 53742
rect 40014 53730 40066 53742
rect 43710 53730 43762 53742
rect 39442 53678 39454 53730
rect 39506 53678 39518 53730
rect 43250 53678 43262 53730
rect 43314 53678 43326 53730
rect 36206 53666 36258 53678
rect 40014 53666 40066 53678
rect 43710 53666 43762 53678
rect 44270 53730 44322 53742
rect 44270 53666 44322 53678
rect 45614 53730 45666 53742
rect 45614 53666 45666 53678
rect 48862 53730 48914 53742
rect 48862 53666 48914 53678
rect 49086 53730 49138 53742
rect 49086 53666 49138 53678
rect 49534 53730 49586 53742
rect 49534 53666 49586 53678
rect 49758 53730 49810 53742
rect 55582 53730 55634 53742
rect 59054 53730 59106 53742
rect 50978 53678 50990 53730
rect 51042 53678 51054 53730
rect 51986 53678 51998 53730
rect 52050 53678 52062 53730
rect 53666 53678 53678 53730
rect 53730 53678 53742 53730
rect 55122 53678 55134 53730
rect 55186 53678 55198 53730
rect 55906 53678 55918 53730
rect 55970 53678 55982 53730
rect 58034 53678 58046 53730
rect 58098 53678 58110 53730
rect 58370 53678 58382 53730
rect 58434 53678 58446 53730
rect 49758 53666 49810 53678
rect 55582 53666 55634 53678
rect 59054 53666 59106 53678
rect 9662 53618 9714 53630
rect 9662 53554 9714 53566
rect 11454 53618 11506 53630
rect 11454 53554 11506 53566
rect 12350 53618 12402 53630
rect 16830 53618 16882 53630
rect 12562 53566 12574 53618
rect 12626 53566 12638 53618
rect 12350 53554 12402 53566
rect 16830 53554 16882 53566
rect 17166 53618 17218 53630
rect 17166 53554 17218 53566
rect 17838 53618 17890 53630
rect 17838 53554 17890 53566
rect 28478 53618 28530 53630
rect 28478 53554 28530 53566
rect 28590 53618 28642 53630
rect 28590 53554 28642 53566
rect 30942 53618 30994 53630
rect 30942 53554 30994 53566
rect 32398 53618 32450 53630
rect 40910 53618 40962 53630
rect 34290 53566 34302 53618
rect 34354 53566 34366 53618
rect 37650 53566 37662 53618
rect 37714 53566 37726 53618
rect 32398 53554 32450 53566
rect 40910 53554 40962 53566
rect 41246 53618 41298 53630
rect 44046 53618 44098 53630
rect 41570 53566 41582 53618
rect 41634 53566 41646 53618
rect 41246 53554 41298 53566
rect 44046 53554 44098 53566
rect 44830 53618 44882 53630
rect 44830 53554 44882 53566
rect 45054 53618 45106 53630
rect 52670 53618 52722 53630
rect 46498 53566 46510 53618
rect 46562 53566 46574 53618
rect 50082 53566 50094 53618
rect 50146 53566 50158 53618
rect 51202 53566 51214 53618
rect 51266 53566 51278 53618
rect 51650 53566 51662 53618
rect 51714 53566 51726 53618
rect 45054 53554 45106 53566
rect 52670 53554 52722 53566
rect 8654 53506 8706 53518
rect 8654 53442 8706 53454
rect 9102 53506 9154 53518
rect 9102 53442 9154 53454
rect 10558 53506 10610 53518
rect 10558 53442 10610 53454
rect 11790 53506 11842 53518
rect 11790 53442 11842 53454
rect 13582 53506 13634 53518
rect 15262 53506 15314 53518
rect 14466 53454 14478 53506
rect 14530 53454 14542 53506
rect 13582 53442 13634 53454
rect 15262 53442 15314 53454
rect 15822 53506 15874 53518
rect 15822 53442 15874 53454
rect 16942 53506 16994 53518
rect 16942 53442 16994 53454
rect 18510 53506 18562 53518
rect 20190 53506 20242 53518
rect 28254 53506 28306 53518
rect 31726 53506 31778 53518
rect 19282 53454 19294 53506
rect 19346 53454 19358 53506
rect 27570 53454 27582 53506
rect 27634 53454 27646 53506
rect 29698 53454 29710 53506
rect 29762 53454 29774 53506
rect 18510 53442 18562 53454
rect 20190 53442 20242 53454
rect 28254 53442 28306 53454
rect 31726 53442 31778 53454
rect 32510 53506 32562 53518
rect 32510 53442 32562 53454
rect 32846 53506 32898 53518
rect 35422 53506 35474 53518
rect 33170 53454 33182 53506
rect 33234 53454 33246 53506
rect 32846 53442 32898 53454
rect 35422 53442 35474 53454
rect 38782 53506 38834 53518
rect 40686 53506 40738 53518
rect 39218 53454 39230 53506
rect 39282 53454 39294 53506
rect 38782 53442 38834 53454
rect 40686 53442 40738 53454
rect 41918 53506 41970 53518
rect 41918 53442 41970 53454
rect 42366 53506 42418 53518
rect 42366 53442 42418 53454
rect 43038 53506 43090 53518
rect 43038 53442 43090 53454
rect 43934 53506 43986 53518
rect 43934 53442 43986 53454
rect 48302 53506 48354 53518
rect 48302 53442 48354 53454
rect 48974 53506 49026 53518
rect 59614 53506 59666 53518
rect 53218 53454 53230 53506
rect 53282 53454 53294 53506
rect 48974 53442 49026 53454
rect 59614 53442 59666 53454
rect 60734 53506 60786 53518
rect 60734 53442 60786 53454
rect 61854 53506 61906 53518
rect 61854 53442 61906 53454
rect 62190 53506 62242 53518
rect 62190 53442 62242 53454
rect 1344 53338 62608 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 62608 53338
rect 1344 53252 62608 53286
rect 9102 53170 9154 53182
rect 9102 53106 9154 53118
rect 9886 53170 9938 53182
rect 9886 53106 9938 53118
rect 19966 53170 20018 53182
rect 19966 53106 20018 53118
rect 25342 53170 25394 53182
rect 25342 53106 25394 53118
rect 25790 53170 25842 53182
rect 25790 53106 25842 53118
rect 25902 53170 25954 53182
rect 25902 53106 25954 53118
rect 27022 53170 27074 53182
rect 29262 53170 29314 53182
rect 28130 53118 28142 53170
rect 28194 53118 28206 53170
rect 27022 53106 27074 53118
rect 29262 53106 29314 53118
rect 29710 53170 29762 53182
rect 46398 53170 46450 53182
rect 45490 53118 45502 53170
rect 45554 53118 45566 53170
rect 29710 53106 29762 53118
rect 46398 53106 46450 53118
rect 53566 53170 53618 53182
rect 53566 53106 53618 53118
rect 53790 53170 53842 53182
rect 53790 53106 53842 53118
rect 60734 53170 60786 53182
rect 60734 53106 60786 53118
rect 15038 53058 15090 53070
rect 17838 53058 17890 53070
rect 25230 53058 25282 53070
rect 32398 53058 32450 53070
rect 40910 53058 40962 53070
rect 46510 53058 46562 53070
rect 16594 53006 16606 53058
rect 16658 53006 16670 53058
rect 18722 53006 18734 53058
rect 18786 53006 18798 53058
rect 22194 53006 22206 53058
rect 22258 53006 22270 53058
rect 26674 53006 26686 53058
rect 26738 53006 26750 53058
rect 38994 53006 39006 53058
rect 39058 53006 39070 53058
rect 39330 53006 39342 53058
rect 39394 53006 39406 53058
rect 42690 53006 42702 53058
rect 42754 53006 42766 53058
rect 45266 53006 45278 53058
rect 45330 53006 45342 53058
rect 15038 52994 15090 53006
rect 17838 52994 17890 53006
rect 25230 52994 25282 53006
rect 32398 52994 32450 53006
rect 40910 52994 40962 53006
rect 46510 52994 46562 53006
rect 46734 53058 46786 53070
rect 46734 52994 46786 53006
rect 47966 53058 48018 53070
rect 53902 53058 53954 53070
rect 57486 53058 57538 53070
rect 49970 53006 49982 53058
rect 50034 53006 50046 53058
rect 55010 53006 55022 53058
rect 55074 53006 55086 53058
rect 58818 53006 58830 53058
rect 58882 53006 58894 53058
rect 47966 52994 48018 53006
rect 53902 52994 53954 53006
rect 57486 52994 57538 53006
rect 7758 52946 7810 52958
rect 15150 52946 15202 52958
rect 14354 52894 14366 52946
rect 14418 52894 14430 52946
rect 7758 52882 7810 52894
rect 15150 52882 15202 52894
rect 15598 52946 15650 52958
rect 15598 52882 15650 52894
rect 15822 52946 15874 52958
rect 20414 52946 20466 52958
rect 16370 52894 16382 52946
rect 16434 52894 16446 52946
rect 15822 52882 15874 52894
rect 20414 52882 20466 52894
rect 20638 52946 20690 52958
rect 20638 52882 20690 52894
rect 21086 52946 21138 52958
rect 25566 52946 25618 52958
rect 21522 52894 21534 52946
rect 21586 52894 21598 52946
rect 23202 52894 23214 52946
rect 23266 52894 23278 52946
rect 21086 52882 21138 52894
rect 25566 52882 25618 52894
rect 26014 52946 26066 52958
rect 26014 52882 26066 52894
rect 26462 52946 26514 52958
rect 32174 52946 32226 52958
rect 30482 52894 30494 52946
rect 30546 52894 30558 52946
rect 31266 52894 31278 52946
rect 31330 52894 31342 52946
rect 26462 52882 26514 52894
rect 32174 52882 32226 52894
rect 32510 52946 32562 52958
rect 32510 52882 32562 52894
rect 33294 52946 33346 52958
rect 33294 52882 33346 52894
rect 33518 52946 33570 52958
rect 33518 52882 33570 52894
rect 33966 52946 34018 52958
rect 33966 52882 34018 52894
rect 34526 52946 34578 52958
rect 45054 52946 45106 52958
rect 46062 52946 46114 52958
rect 48190 52946 48242 52958
rect 49422 52946 49474 52958
rect 50990 52946 51042 52958
rect 35074 52894 35086 52946
rect 35138 52894 35150 52946
rect 40114 52894 40126 52946
rect 40178 52894 40190 52946
rect 41122 52894 41134 52946
rect 41186 52894 41198 52946
rect 45826 52894 45838 52946
rect 45890 52894 45902 52946
rect 47506 52894 47518 52946
rect 47570 52894 47582 52946
rect 47730 52894 47742 52946
rect 47794 52894 47806 52946
rect 49186 52894 49198 52946
rect 49250 52894 49262 52946
rect 49858 52894 49870 52946
rect 49922 52894 49934 52946
rect 34526 52882 34578 52894
rect 45054 52882 45106 52894
rect 46062 52882 46114 52894
rect 48190 52882 48242 52894
rect 49422 52882 49474 52894
rect 50990 52882 51042 52894
rect 51326 52946 51378 52958
rect 51326 52882 51378 52894
rect 51550 52946 51602 52958
rect 56814 52946 56866 52958
rect 51986 52894 51998 52946
rect 52050 52894 52062 52946
rect 52546 52894 52558 52946
rect 52610 52894 52622 52946
rect 54226 52894 54238 52946
rect 54290 52894 54302 52946
rect 54786 52894 54798 52946
rect 54850 52894 54862 52946
rect 51550 52882 51602 52894
rect 56814 52882 56866 52894
rect 57822 52946 57874 52958
rect 59042 52894 59054 52946
rect 59106 52894 59118 52946
rect 59602 52894 59614 52946
rect 59666 52894 59678 52946
rect 57822 52882 57874 52894
rect 8094 52834 8146 52846
rect 8094 52770 8146 52782
rect 8542 52834 8594 52846
rect 8542 52770 8594 52782
rect 10446 52834 10498 52846
rect 10446 52770 10498 52782
rect 10894 52834 10946 52846
rect 10894 52770 10946 52782
rect 11230 52834 11282 52846
rect 20526 52834 20578 52846
rect 33406 52834 33458 52846
rect 11554 52782 11566 52834
rect 11618 52782 11630 52834
rect 13682 52782 13694 52834
rect 13746 52782 13758 52834
rect 17490 52782 17502 52834
rect 17554 52782 17566 52834
rect 23314 52782 23326 52834
rect 23378 52782 23390 52834
rect 30146 52782 30158 52834
rect 30210 52782 30222 52834
rect 31490 52782 31502 52834
rect 31554 52782 31566 52834
rect 11230 52770 11282 52782
rect 20526 52770 20578 52782
rect 33406 52770 33458 52782
rect 34750 52834 34802 52846
rect 41694 52834 41746 52846
rect 35858 52782 35870 52834
rect 35922 52782 35934 52834
rect 37986 52782 37998 52834
rect 38050 52782 38062 52834
rect 40002 52782 40014 52834
rect 40066 52782 40078 52834
rect 34750 52770 34802 52782
rect 41694 52770 41746 52782
rect 44270 52834 44322 52846
rect 51102 52834 51154 52846
rect 56590 52834 56642 52846
rect 44594 52782 44606 52834
rect 44658 52782 44670 52834
rect 47842 52782 47854 52834
rect 47906 52782 47918 52834
rect 50194 52782 50206 52834
rect 50258 52782 50270 52834
rect 52098 52782 52110 52834
rect 52162 52782 52174 52834
rect 52434 52782 52446 52834
rect 52498 52782 52510 52834
rect 54338 52782 54350 52834
rect 54402 52782 54414 52834
rect 44270 52770 44322 52782
rect 51102 52770 51154 52782
rect 56590 52770 56642 52782
rect 58382 52834 58434 52846
rect 60286 52834 60338 52846
rect 58930 52782 58942 52834
rect 58994 52782 59006 52834
rect 58382 52770 58434 52782
rect 60286 52770 60338 52782
rect 61294 52834 61346 52846
rect 61294 52770 61346 52782
rect 61966 52834 62018 52846
rect 61966 52770 62018 52782
rect 15150 52722 15202 52734
rect 38446 52722 38498 52734
rect 10098 52670 10110 52722
rect 10162 52719 10174 52722
rect 11330 52719 11342 52722
rect 10162 52673 11342 52719
rect 10162 52670 10174 52673
rect 11330 52670 11342 52673
rect 11394 52670 11406 52722
rect 21410 52670 21422 52722
rect 21474 52670 21486 52722
rect 31602 52670 31614 52722
rect 31666 52670 31678 52722
rect 34178 52670 34190 52722
rect 34242 52670 34254 52722
rect 15150 52658 15202 52670
rect 38446 52658 38498 52670
rect 38782 52722 38834 52734
rect 38782 52658 38834 52670
rect 43822 52722 43874 52734
rect 55582 52722 55634 52734
rect 45602 52670 45614 52722
rect 45666 52670 45678 52722
rect 43822 52658 43874 52670
rect 55582 52658 55634 52670
rect 55918 52722 55970 52734
rect 57138 52670 57150 52722
rect 57202 52670 57214 52722
rect 55918 52658 55970 52670
rect 1344 52554 62608 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 62608 52554
rect 1344 52468 62608 52502
rect 37102 52386 37154 52398
rect 7858 52334 7870 52386
rect 7922 52383 7934 52386
rect 8306 52383 8318 52386
rect 7922 52337 8318 52383
rect 7922 52334 7934 52337
rect 8306 52334 8318 52337
rect 8370 52334 8382 52386
rect 23090 52334 23102 52386
rect 23154 52334 23166 52386
rect 50082 52334 50094 52386
rect 50146 52334 50158 52386
rect 37102 52322 37154 52334
rect 6862 52274 6914 52286
rect 6862 52210 6914 52222
rect 8318 52274 8370 52286
rect 8318 52210 8370 52222
rect 9102 52274 9154 52286
rect 9102 52210 9154 52222
rect 9550 52274 9602 52286
rect 9550 52210 9602 52222
rect 14366 52274 14418 52286
rect 22206 52274 22258 52286
rect 44270 52274 44322 52286
rect 15250 52222 15262 52274
rect 15314 52222 15326 52274
rect 15698 52222 15710 52274
rect 15762 52222 15774 52274
rect 17602 52222 17614 52274
rect 17666 52222 17678 52274
rect 19730 52222 19742 52274
rect 19794 52222 19806 52274
rect 23314 52222 23326 52274
rect 23378 52222 23390 52274
rect 23986 52222 23998 52274
rect 24050 52222 24062 52274
rect 28242 52222 28254 52274
rect 28306 52222 28318 52274
rect 32722 52222 32734 52274
rect 32786 52222 32798 52274
rect 43138 52222 43150 52274
rect 43202 52222 43214 52274
rect 14366 52210 14418 52222
rect 22206 52210 22258 52222
rect 44270 52210 44322 52222
rect 45390 52274 45442 52286
rect 55694 52274 55746 52286
rect 60734 52274 60786 52286
rect 47282 52222 47294 52274
rect 47346 52222 47358 52274
rect 58258 52222 58270 52274
rect 58322 52222 58334 52274
rect 45390 52210 45442 52222
rect 55694 52210 55746 52222
rect 60734 52210 60786 52222
rect 61070 52274 61122 52286
rect 61070 52210 61122 52222
rect 61518 52274 61570 52286
rect 61518 52210 61570 52222
rect 7422 52162 7474 52174
rect 7422 52098 7474 52110
rect 10110 52162 10162 52174
rect 10110 52098 10162 52110
rect 13694 52162 13746 52174
rect 13694 52098 13746 52110
rect 13806 52162 13858 52174
rect 15822 52162 15874 52174
rect 21198 52162 21250 52174
rect 23662 52162 23714 52174
rect 32510 52162 32562 52174
rect 35086 52162 35138 52174
rect 35758 52162 35810 52174
rect 45166 52162 45218 52174
rect 15138 52110 15150 52162
rect 15202 52110 15214 52162
rect 16034 52110 16046 52162
rect 16098 52110 16110 52162
rect 20514 52110 20526 52162
rect 20578 52110 20590 52162
rect 21858 52110 21870 52162
rect 21922 52110 21934 52162
rect 24322 52110 24334 52162
rect 24386 52110 24398 52162
rect 25330 52110 25342 52162
rect 25394 52110 25406 52162
rect 29922 52110 29934 52162
rect 29986 52110 29998 52162
rect 32162 52110 32174 52162
rect 32226 52110 32238 52162
rect 32834 52110 32846 52162
rect 32898 52110 32910 52162
rect 34850 52110 34862 52162
rect 34914 52110 34926 52162
rect 35410 52110 35422 52162
rect 35474 52110 35486 52162
rect 36194 52110 36206 52162
rect 36258 52110 36270 52162
rect 36978 52110 36990 52162
rect 37042 52110 37054 52162
rect 40338 52110 40350 52162
rect 40402 52110 40414 52162
rect 43698 52110 43710 52162
rect 43762 52110 43774 52162
rect 13806 52098 13858 52110
rect 15822 52098 15874 52110
rect 21198 52098 21250 52110
rect 23662 52098 23714 52110
rect 32510 52098 32562 52110
rect 35086 52098 35138 52110
rect 35758 52098 35810 52110
rect 45166 52098 45218 52110
rect 45726 52162 45778 52174
rect 45726 52098 45778 52110
rect 45950 52162 46002 52174
rect 45950 52098 46002 52110
rect 46734 52162 46786 52174
rect 52558 52162 52610 52174
rect 48290 52110 48302 52162
rect 48354 52110 48366 52162
rect 48850 52110 48862 52162
rect 48914 52110 48926 52162
rect 49970 52110 49982 52162
rect 50034 52110 50046 52162
rect 51874 52110 51886 52162
rect 51938 52110 51950 52162
rect 46734 52098 46786 52110
rect 52558 52098 52610 52110
rect 52782 52162 52834 52174
rect 52782 52098 52834 52110
rect 52894 52162 52946 52174
rect 52894 52098 52946 52110
rect 53118 52162 53170 52174
rect 53118 52098 53170 52110
rect 53454 52162 53506 52174
rect 53454 52098 53506 52110
rect 53902 52162 53954 52174
rect 59614 52162 59666 52174
rect 54786 52110 54798 52162
rect 54850 52110 54862 52162
rect 55458 52110 55470 52162
rect 55522 52110 55534 52162
rect 57698 52110 57710 52162
rect 57762 52110 57774 52162
rect 58818 52110 58830 52162
rect 58882 52110 58894 52162
rect 53902 52098 53954 52110
rect 59614 52098 59666 52110
rect 12574 52050 12626 52062
rect 11666 51998 11678 52050
rect 11730 51998 11742 52050
rect 12574 51986 12626 51998
rect 12910 52050 12962 52062
rect 12910 51986 12962 51998
rect 14478 52050 14530 52062
rect 14478 51986 14530 51998
rect 17278 52050 17330 52062
rect 17278 51986 17330 51998
rect 21534 52050 21586 52062
rect 24558 52050 24610 52062
rect 24210 51998 24222 52050
rect 24274 51998 24286 52050
rect 21534 51986 21586 51998
rect 24558 51986 24610 51998
rect 24782 52050 24834 52062
rect 29150 52050 29202 52062
rect 26114 51998 26126 52050
rect 26178 51998 26190 52050
rect 24782 51986 24834 51998
rect 29150 51986 29202 51998
rect 30270 52050 30322 52062
rect 30270 51986 30322 51998
rect 30382 52050 30434 52062
rect 30382 51986 30434 51998
rect 30606 52050 30658 52062
rect 34638 52050 34690 52062
rect 43486 52050 43538 52062
rect 31826 51998 31838 52050
rect 31890 51998 31902 52050
rect 38434 51998 38446 52050
rect 38498 51998 38510 52050
rect 41010 51998 41022 52050
rect 41074 51998 41086 52050
rect 30606 51986 30658 51998
rect 34638 51986 34690 51998
rect 43486 51986 43538 51998
rect 48078 52050 48130 52062
rect 54126 52050 54178 52062
rect 51538 51998 51550 52050
rect 51602 51998 51614 52050
rect 48078 51986 48130 51998
rect 54126 51986 54178 51998
rect 7870 51938 7922 51950
rect 7870 51874 7922 51886
rect 8766 51938 8818 51950
rect 8766 51874 8818 51886
rect 10446 51938 10498 51950
rect 10446 51874 10498 51886
rect 14254 51938 14306 51950
rect 14254 51874 14306 51886
rect 16942 51938 16994 51950
rect 16942 51874 16994 51886
rect 21422 51938 21474 51950
rect 21422 51874 21474 51886
rect 29262 51938 29314 51950
rect 29262 51874 29314 51886
rect 30494 51938 30546 51950
rect 30494 51874 30546 51886
rect 35422 51938 35474 51950
rect 35422 51874 35474 51886
rect 39790 51938 39842 51950
rect 47742 51938 47794 51950
rect 44818 51886 44830 51938
rect 44882 51886 44894 51938
rect 46274 51886 46286 51938
rect 46338 51886 46350 51938
rect 39790 51874 39842 51886
rect 47742 51874 47794 51886
rect 53678 51938 53730 51950
rect 53678 51874 53730 51886
rect 58830 51938 58882 51950
rect 58830 51874 58882 51886
rect 60062 51938 60114 51950
rect 60062 51874 60114 51886
rect 61966 51938 62018 51950
rect 61966 51874 62018 51886
rect 1344 51770 62608 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 62608 51770
rect 1344 51684 62608 51718
rect 4846 51602 4898 51614
rect 4846 51538 4898 51550
rect 5854 51602 5906 51614
rect 5854 51538 5906 51550
rect 7198 51602 7250 51614
rect 7198 51538 7250 51550
rect 8206 51602 8258 51614
rect 8206 51538 8258 51550
rect 8654 51602 8706 51614
rect 13470 51602 13522 51614
rect 10210 51550 10222 51602
rect 10274 51550 10286 51602
rect 8654 51538 8706 51550
rect 13470 51538 13522 51550
rect 17502 51602 17554 51614
rect 23438 51602 23490 51614
rect 26350 51602 26402 51614
rect 18946 51550 18958 51602
rect 19010 51550 19022 51602
rect 20066 51550 20078 51602
rect 20130 51550 20142 51602
rect 25218 51550 25230 51602
rect 25282 51550 25294 51602
rect 17502 51538 17554 51550
rect 23438 51538 23490 51550
rect 26350 51538 26402 51550
rect 26574 51602 26626 51614
rect 28926 51602 28978 51614
rect 27794 51550 27806 51602
rect 27858 51550 27870 51602
rect 26574 51538 26626 51550
rect 28926 51538 28978 51550
rect 29374 51602 29426 51614
rect 29374 51538 29426 51550
rect 29598 51602 29650 51614
rect 29598 51538 29650 51550
rect 32398 51602 32450 51614
rect 32398 51538 32450 51550
rect 39790 51602 39842 51614
rect 39790 51538 39842 51550
rect 40238 51602 40290 51614
rect 40238 51538 40290 51550
rect 43150 51602 43202 51614
rect 43150 51538 43202 51550
rect 44718 51602 44770 51614
rect 44718 51538 44770 51550
rect 44942 51602 44994 51614
rect 47742 51602 47794 51614
rect 45826 51550 45838 51602
rect 45890 51550 45902 51602
rect 44942 51538 44994 51550
rect 47742 51538 47794 51550
rect 61294 51602 61346 51614
rect 61294 51538 61346 51550
rect 17390 51490 17442 51502
rect 31614 51490 31666 51502
rect 36766 51490 36818 51502
rect 44606 51490 44658 51502
rect 60846 51490 60898 51502
rect 18274 51438 18286 51490
rect 18338 51438 18350 51490
rect 21522 51438 21534 51490
rect 21586 51438 21598 51490
rect 24546 51438 24558 51490
rect 24610 51438 24622 51490
rect 30258 51438 30270 51490
rect 30322 51438 30334 51490
rect 33954 51438 33966 51490
rect 34018 51438 34030 51490
rect 38098 51438 38110 51490
rect 38162 51438 38174 51490
rect 38322 51438 38334 51490
rect 38386 51438 38398 51490
rect 39442 51438 39454 51490
rect 39506 51438 39518 51490
rect 41906 51438 41918 51490
rect 41970 51438 41982 51490
rect 53330 51438 53342 51490
rect 53394 51438 53406 51490
rect 17390 51426 17442 51438
rect 31614 51426 31666 51438
rect 36766 51426 36818 51438
rect 44606 51426 44658 51438
rect 60846 51426 60898 51438
rect 13358 51378 13410 51390
rect 13358 51314 13410 51326
rect 13694 51378 13746 51390
rect 23774 51378 23826 51390
rect 26686 51378 26738 51390
rect 14018 51326 14030 51378
rect 14082 51326 14094 51378
rect 17938 51326 17950 51378
rect 18002 51326 18014 51378
rect 18834 51326 18846 51378
rect 18898 51326 18910 51378
rect 22978 51326 22990 51378
rect 23042 51326 23054 51378
rect 24434 51326 24446 51378
rect 24498 51326 24510 51378
rect 25442 51326 25454 51378
rect 25506 51326 25518 51378
rect 13694 51314 13746 51326
rect 23774 51314 23826 51326
rect 26686 51314 26738 51326
rect 26798 51378 26850 51390
rect 31278 51378 31330 51390
rect 29810 51326 29822 51378
rect 29874 51326 29886 51378
rect 26798 51314 26850 51326
rect 31278 51314 31330 51326
rect 32062 51378 32114 51390
rect 32062 51314 32114 51326
rect 32174 51378 32226 51390
rect 32174 51314 32226 51326
rect 32510 51378 32562 51390
rect 38670 51378 38722 51390
rect 54350 51378 54402 51390
rect 33506 51326 33518 51378
rect 33570 51326 33582 51378
rect 34962 51326 34974 51378
rect 35026 51326 35038 51378
rect 36418 51326 36430 51378
rect 36482 51326 36494 51378
rect 37090 51326 37102 51378
rect 37154 51326 37166 51378
rect 43810 51326 43822 51378
rect 43874 51326 43886 51378
rect 49186 51326 49198 51378
rect 49250 51326 49262 51378
rect 53554 51326 53566 51378
rect 53618 51326 53630 51378
rect 54562 51326 54574 51378
rect 54626 51326 54638 51378
rect 57026 51326 57038 51378
rect 57090 51326 57102 51378
rect 32510 51314 32562 51326
rect 38670 51314 38722 51326
rect 54350 51314 54402 51326
rect 2942 51266 2994 51278
rect 2942 51202 2994 51214
rect 4174 51266 4226 51278
rect 4174 51202 4226 51214
rect 6414 51266 6466 51278
rect 6414 51202 6466 51214
rect 6862 51266 6914 51278
rect 6862 51202 6914 51214
rect 7646 51266 7698 51278
rect 7646 51202 7698 51214
rect 9102 51266 9154 51278
rect 9102 51202 9154 51214
rect 12686 51266 12738 51278
rect 29710 51266 29762 51278
rect 12898 51214 12910 51266
rect 12962 51214 12974 51266
rect 14690 51214 14702 51266
rect 14754 51214 14766 51266
rect 16818 51214 16830 51266
rect 16882 51214 16894 51266
rect 22642 51214 22654 51266
rect 22706 51214 22718 51266
rect 12686 51202 12738 51214
rect 29710 51202 29762 51214
rect 41022 51266 41074 51278
rect 41022 51202 41074 51214
rect 44270 51266 44322 51278
rect 44270 51202 44322 51214
rect 48974 51266 49026 51278
rect 56702 51266 56754 51278
rect 60398 51266 60450 51278
rect 49970 51214 49982 51266
rect 50034 51214 50046 51266
rect 52098 51214 52110 51266
rect 52162 51214 52174 51266
rect 57810 51214 57822 51266
rect 57874 51214 57886 51266
rect 59938 51214 59950 51266
rect 60002 51214 60014 51266
rect 48974 51202 49026 51214
rect 56702 51202 56754 51214
rect 60398 51202 60450 51214
rect 61742 51266 61794 51278
rect 61742 51202 61794 51214
rect 62190 51266 62242 51278
rect 62190 51202 62242 51214
rect 12126 51154 12178 51166
rect 12126 51090 12178 51102
rect 17502 51154 17554 51166
rect 37102 51154 37154 51166
rect 30594 51102 30606 51154
rect 30658 51102 30670 51154
rect 33618 51102 33630 51154
rect 33682 51102 33694 51154
rect 17502 51090 17554 51102
rect 37102 51090 37154 51102
rect 39006 51154 39058 51166
rect 55010 51102 55022 51154
rect 55074 51102 55086 51154
rect 60386 51102 60398 51154
rect 60450 51151 60462 51154
rect 61954 51151 61966 51154
rect 60450 51105 61966 51151
rect 60450 51102 60462 51105
rect 61954 51102 61966 51105
rect 62018 51102 62030 51154
rect 39006 51090 39058 51102
rect 1344 50986 62608 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 62608 50986
rect 1344 50900 62608 50934
rect 22542 50818 22594 50830
rect 3602 50766 3614 50818
rect 3666 50815 3678 50818
rect 4498 50815 4510 50818
rect 3666 50769 4510 50815
rect 3666 50766 3678 50769
rect 4498 50766 4510 50769
rect 4562 50766 4574 50818
rect 22542 50754 22594 50766
rect 22878 50818 22930 50830
rect 22878 50754 22930 50766
rect 24334 50818 24386 50830
rect 24334 50754 24386 50766
rect 34526 50818 34578 50830
rect 34526 50754 34578 50766
rect 36094 50818 36146 50830
rect 36094 50754 36146 50766
rect 47630 50818 47682 50830
rect 47630 50754 47682 50766
rect 49422 50818 49474 50830
rect 50866 50766 50878 50818
rect 50930 50766 50942 50818
rect 60498 50766 60510 50818
rect 60562 50815 60574 50818
rect 61282 50815 61294 50818
rect 60562 50769 61294 50815
rect 60562 50766 60574 50769
rect 61282 50766 61294 50769
rect 61346 50766 61358 50818
rect 49422 50754 49474 50766
rect 6190 50706 6242 50718
rect 6190 50642 6242 50654
rect 7870 50706 7922 50718
rect 7870 50642 7922 50654
rect 15822 50706 15874 50718
rect 36318 50706 36370 50718
rect 31378 50654 31390 50706
rect 31442 50654 31454 50706
rect 33506 50654 33518 50706
rect 33570 50654 33582 50706
rect 34738 50654 34750 50706
rect 34802 50654 34814 50706
rect 15822 50642 15874 50654
rect 36318 50642 36370 50654
rect 39790 50706 39842 50718
rect 39790 50642 39842 50654
rect 40350 50706 40402 50718
rect 40350 50642 40402 50654
rect 41694 50706 41746 50718
rect 41694 50642 41746 50654
rect 46398 50706 46450 50718
rect 59950 50706 60002 50718
rect 47506 50654 47518 50706
rect 47570 50654 47582 50706
rect 49746 50654 49758 50706
rect 49810 50654 49822 50706
rect 53218 50654 53230 50706
rect 53282 50654 53294 50706
rect 46398 50642 46450 50654
rect 59950 50642 60002 50654
rect 60622 50706 60674 50718
rect 60622 50642 60674 50654
rect 61518 50706 61570 50718
rect 61518 50642 61570 50654
rect 61966 50706 62018 50718
rect 61966 50642 62018 50654
rect 5182 50594 5234 50606
rect 5182 50530 5234 50542
rect 7086 50594 7138 50606
rect 9886 50594 9938 50606
rect 9314 50542 9326 50594
rect 9378 50542 9390 50594
rect 7086 50530 7138 50542
rect 9886 50530 9938 50542
rect 10110 50594 10162 50606
rect 10110 50530 10162 50542
rect 13022 50594 13074 50606
rect 14366 50594 14418 50606
rect 13794 50542 13806 50594
rect 13858 50542 13870 50594
rect 13022 50530 13074 50542
rect 14366 50530 14418 50542
rect 15150 50594 15202 50606
rect 15150 50530 15202 50542
rect 15486 50594 15538 50606
rect 15486 50530 15538 50542
rect 15934 50594 15986 50606
rect 15934 50530 15986 50542
rect 20526 50594 20578 50606
rect 23326 50594 23378 50606
rect 25790 50594 25842 50606
rect 28030 50594 28082 50606
rect 21858 50542 21870 50594
rect 21922 50542 21934 50594
rect 24434 50542 24446 50594
rect 24498 50542 24510 50594
rect 26226 50542 26238 50594
rect 26290 50542 26302 50594
rect 20526 50530 20578 50542
rect 23326 50530 23378 50542
rect 25790 50530 25842 50542
rect 28030 50530 28082 50542
rect 28590 50594 28642 50606
rect 34638 50594 34690 50606
rect 29698 50542 29710 50594
rect 29762 50542 29774 50594
rect 30594 50542 30606 50594
rect 30658 50542 30670 50594
rect 30930 50542 30942 50594
rect 30994 50542 31006 50594
rect 33394 50542 33406 50594
rect 33458 50542 33470 50594
rect 28590 50530 28642 50542
rect 34638 50530 34690 50542
rect 35086 50594 35138 50606
rect 35086 50530 35138 50542
rect 35310 50594 35362 50606
rect 35310 50530 35362 50542
rect 40014 50594 40066 50606
rect 40014 50530 40066 50542
rect 41246 50594 41298 50606
rect 41246 50530 41298 50542
rect 42478 50594 42530 50606
rect 42478 50530 42530 50542
rect 42702 50594 42754 50606
rect 43710 50594 43762 50606
rect 43250 50542 43262 50594
rect 43314 50542 43326 50594
rect 42702 50530 42754 50542
rect 43710 50530 43762 50542
rect 44270 50594 44322 50606
rect 49198 50594 49250 50606
rect 45938 50542 45950 50594
rect 46002 50542 46014 50594
rect 47170 50542 47182 50594
rect 47234 50542 47246 50594
rect 48066 50542 48078 50594
rect 48130 50542 48142 50594
rect 48514 50542 48526 50594
rect 48578 50542 48590 50594
rect 44270 50530 44322 50542
rect 49198 50530 49250 50542
rect 50318 50594 50370 50606
rect 50318 50530 50370 50542
rect 50654 50594 50706 50606
rect 51438 50594 51490 50606
rect 50978 50542 50990 50594
rect 51042 50542 51054 50594
rect 50654 50530 50706 50542
rect 51438 50530 51490 50542
rect 51662 50594 51714 50606
rect 55694 50594 55746 50606
rect 52994 50542 53006 50594
rect 53058 50542 53070 50594
rect 54226 50542 54238 50594
rect 54290 50542 54302 50594
rect 55234 50542 55246 50594
rect 55298 50542 55310 50594
rect 58034 50542 58046 50594
rect 58098 50542 58110 50594
rect 58706 50542 58718 50594
rect 58770 50542 58782 50594
rect 59378 50542 59390 50594
rect 59442 50542 59454 50594
rect 51662 50530 51714 50542
rect 55694 50530 55746 50542
rect 3614 50482 3666 50494
rect 3614 50418 3666 50430
rect 4398 50482 4450 50494
rect 4398 50418 4450 50430
rect 6638 50482 6690 50494
rect 6638 50418 6690 50430
rect 8430 50482 8482 50494
rect 8430 50418 8482 50430
rect 8654 50482 8706 50494
rect 8654 50418 8706 50430
rect 8766 50482 8818 50494
rect 8766 50418 8818 50430
rect 8990 50482 9042 50494
rect 8990 50418 9042 50430
rect 9550 50482 9602 50494
rect 15262 50482 15314 50494
rect 11218 50430 11230 50482
rect 11282 50430 11294 50482
rect 13570 50430 13582 50482
rect 13634 50430 13646 50482
rect 9550 50418 9602 50430
rect 15262 50418 15314 50430
rect 15710 50482 15762 50494
rect 15710 50418 15762 50430
rect 16158 50482 16210 50494
rect 20638 50482 20690 50494
rect 18722 50430 18734 50482
rect 18786 50430 18798 50482
rect 16158 50418 16210 50430
rect 20638 50418 20690 50430
rect 20750 50482 20802 50494
rect 29374 50482 29426 50494
rect 40798 50482 40850 50494
rect 21746 50430 21758 50482
rect 21810 50430 21822 50482
rect 24994 50430 25006 50482
rect 25058 50430 25070 50482
rect 37314 50430 37326 50482
rect 37378 50430 37390 50482
rect 20750 50418 20802 50430
rect 29374 50418 29426 50430
rect 40798 50418 40850 50430
rect 41022 50482 41074 50494
rect 41022 50418 41074 50430
rect 43038 50482 43090 50494
rect 48414 50482 48466 50494
rect 45042 50430 45054 50482
rect 45106 50430 45118 50482
rect 45826 50430 45838 50482
rect 45890 50430 45902 50482
rect 43038 50418 43090 50430
rect 48414 50418 48466 50430
rect 49758 50482 49810 50494
rect 49758 50418 49810 50430
rect 49982 50482 50034 50494
rect 49982 50418 50034 50430
rect 51886 50482 51938 50494
rect 58494 50482 58546 50494
rect 56914 50430 56926 50482
rect 56978 50430 56990 50482
rect 51886 50418 51938 50430
rect 58494 50418 58546 50430
rect 59166 50482 59218 50494
rect 59166 50418 59218 50430
rect 61182 50482 61234 50494
rect 61182 50418 61234 50430
rect 1934 50370 1986 50382
rect 1934 50306 1986 50318
rect 2382 50370 2434 50382
rect 2382 50306 2434 50318
rect 2830 50370 2882 50382
rect 2830 50306 2882 50318
rect 4062 50370 4114 50382
rect 4062 50306 4114 50318
rect 7534 50370 7586 50382
rect 14702 50370 14754 50382
rect 10434 50318 10446 50370
rect 10498 50318 10510 50370
rect 7534 50306 7586 50318
rect 14702 50306 14754 50318
rect 16830 50370 16882 50382
rect 16830 50306 16882 50318
rect 19966 50370 20018 50382
rect 19966 50306 20018 50318
rect 20302 50370 20354 50382
rect 39118 50370 39170 50382
rect 23650 50318 23662 50370
rect 23714 50318 23726 50370
rect 35746 50318 35758 50370
rect 35810 50318 35822 50370
rect 20302 50306 20354 50318
rect 39118 50306 39170 50318
rect 41134 50370 41186 50382
rect 50430 50370 50482 50382
rect 42130 50318 42142 50370
rect 42194 50318 42206 50370
rect 45154 50318 45166 50370
rect 45218 50318 45230 50370
rect 41134 50306 41186 50318
rect 50430 50306 50482 50318
rect 51550 50370 51602 50382
rect 57810 50318 57822 50370
rect 57874 50318 57886 50370
rect 51550 50306 51602 50318
rect 1344 50202 62608 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 62608 50202
rect 1344 50116 62608 50150
rect 3054 50034 3106 50046
rect 3054 49970 3106 49982
rect 5966 50034 6018 50046
rect 5966 49970 6018 49982
rect 6414 50034 6466 50046
rect 6414 49970 6466 49982
rect 6750 50034 6802 50046
rect 6750 49970 6802 49982
rect 7310 50034 7362 50046
rect 7310 49970 7362 49982
rect 8094 50034 8146 50046
rect 11566 50034 11618 50046
rect 10210 49982 10222 50034
rect 10274 49982 10286 50034
rect 8094 49970 8146 49982
rect 11566 49970 11618 49982
rect 16718 50034 16770 50046
rect 16718 49970 16770 49982
rect 25678 50034 25730 50046
rect 30718 50034 30770 50046
rect 27122 49982 27134 50034
rect 27186 49982 27198 50034
rect 25678 49970 25730 49982
rect 30718 49970 30770 49982
rect 30830 50034 30882 50046
rect 30830 49970 30882 49982
rect 31278 50034 31330 50046
rect 31278 49970 31330 49982
rect 33406 50034 33458 50046
rect 33406 49970 33458 49982
rect 38446 50034 38498 50046
rect 51214 50034 51266 50046
rect 49746 49982 49758 50034
rect 49810 49982 49822 50034
rect 38446 49970 38498 49982
rect 51214 49970 51266 49982
rect 51438 50034 51490 50046
rect 51438 49970 51490 49982
rect 54798 50034 54850 50046
rect 61854 50034 61906 50046
rect 56578 49982 56590 50034
rect 56642 49982 56654 50034
rect 54798 49970 54850 49982
rect 61854 49970 61906 49982
rect 2382 49922 2434 49934
rect 16494 49922 16546 49934
rect 3378 49870 3390 49922
rect 3442 49870 3454 49922
rect 12674 49870 12686 49922
rect 12738 49870 12750 49922
rect 16370 49870 16382 49922
rect 16434 49870 16446 49922
rect 2382 49858 2434 49870
rect 16494 49858 16546 49870
rect 16606 49922 16658 49934
rect 22430 49922 22482 49934
rect 30494 49922 30546 49934
rect 18386 49870 18398 49922
rect 18450 49870 18462 49922
rect 21410 49870 21422 49922
rect 21474 49870 21486 49922
rect 30258 49870 30270 49922
rect 30322 49870 30334 49922
rect 16606 49858 16658 49870
rect 22430 49858 22482 49870
rect 30494 49858 30546 49870
rect 30606 49922 30658 49934
rect 33070 49922 33122 49934
rect 31938 49870 31950 49922
rect 32002 49870 32014 49922
rect 32386 49870 32398 49922
rect 32450 49870 32462 49922
rect 30606 49858 30658 49870
rect 33070 49858 33122 49870
rect 33182 49922 33234 49934
rect 38894 49922 38946 49934
rect 33730 49870 33742 49922
rect 33794 49870 33806 49922
rect 36642 49870 36654 49922
rect 36706 49870 36718 49922
rect 33182 49858 33234 49870
rect 38894 49858 38946 49870
rect 40350 49922 40402 49934
rect 51662 49922 51714 49934
rect 48850 49870 48862 49922
rect 48914 49870 48926 49922
rect 40350 49858 40402 49870
rect 51662 49858 51714 49870
rect 51774 49922 51826 49934
rect 52882 49870 52894 49922
rect 52946 49870 52958 49922
rect 55682 49870 55694 49922
rect 55746 49870 55758 49922
rect 51774 49858 51826 49870
rect 2718 49810 2770 49822
rect 2718 49746 2770 49758
rect 8430 49810 8482 49822
rect 8430 49746 8482 49758
rect 8654 49810 8706 49822
rect 8654 49746 8706 49758
rect 9102 49810 9154 49822
rect 13246 49810 13298 49822
rect 12450 49758 12462 49810
rect 12514 49758 12526 49810
rect 9102 49746 9154 49758
rect 13246 49746 13298 49758
rect 13918 49810 13970 49822
rect 13918 49746 13970 49758
rect 14366 49810 14418 49822
rect 14366 49746 14418 49758
rect 14590 49810 14642 49822
rect 16830 49810 16882 49822
rect 15698 49758 15710 49810
rect 15762 49758 15774 49810
rect 14590 49746 14642 49758
rect 16830 49746 16882 49758
rect 19518 49810 19570 49822
rect 25566 49810 25618 49822
rect 20290 49758 20302 49810
rect 20354 49758 20366 49810
rect 21746 49758 21758 49810
rect 21810 49758 21822 49810
rect 22754 49758 22766 49810
rect 22818 49758 22830 49810
rect 24098 49758 24110 49810
rect 24162 49758 24174 49810
rect 25218 49758 25230 49810
rect 25282 49758 25294 49810
rect 19518 49746 19570 49758
rect 25566 49746 25618 49758
rect 25790 49810 25842 49822
rect 25790 49746 25842 49758
rect 31614 49810 31666 49822
rect 39902 49810 39954 49822
rect 42814 49810 42866 49822
rect 47406 49810 47458 49822
rect 34178 49758 34190 49810
rect 34242 49758 34254 49810
rect 34738 49758 34750 49810
rect 34802 49758 34814 49810
rect 35522 49758 35534 49810
rect 35586 49758 35598 49810
rect 41010 49758 41022 49810
rect 41074 49758 41086 49810
rect 42130 49758 42142 49810
rect 42194 49758 42206 49810
rect 43586 49758 43598 49810
rect 43650 49758 43662 49810
rect 44818 49758 44830 49810
rect 44882 49758 44894 49810
rect 45714 49758 45726 49810
rect 45778 49758 45790 49810
rect 31614 49746 31666 49758
rect 39902 49746 39954 49758
rect 42814 49746 42866 49758
rect 47406 49746 47458 49758
rect 47742 49810 47794 49822
rect 50430 49810 50482 49822
rect 49186 49758 49198 49810
rect 49250 49758 49262 49810
rect 49634 49758 49646 49810
rect 49698 49758 49710 49810
rect 47742 49746 47794 49758
rect 50430 49746 50482 49758
rect 50766 49810 50818 49822
rect 54238 49810 54290 49822
rect 56926 49810 56978 49822
rect 50978 49758 50990 49810
rect 51042 49758 51054 49810
rect 55794 49758 55806 49810
rect 55858 49758 55870 49810
rect 50766 49746 50818 49758
rect 54238 49746 54290 49758
rect 56926 49746 56978 49758
rect 57150 49810 57202 49822
rect 57150 49746 57202 49758
rect 58046 49810 58098 49822
rect 58046 49746 58098 49758
rect 58270 49810 58322 49822
rect 58270 49746 58322 49758
rect 58718 49810 58770 49822
rect 58718 49746 58770 49758
rect 58942 49810 58994 49822
rect 58942 49746 58994 49758
rect 59838 49810 59890 49822
rect 61282 49758 61294 49810
rect 61346 49758 61358 49810
rect 59838 49746 59890 49758
rect 1822 49698 1874 49710
rect 1822 49634 1874 49646
rect 3950 49698 4002 49710
rect 3950 49634 4002 49646
rect 4510 49698 4562 49710
rect 4510 49634 4562 49646
rect 4958 49698 5010 49710
rect 4958 49634 5010 49646
rect 5518 49698 5570 49710
rect 5518 49634 5570 49646
rect 7758 49698 7810 49710
rect 7758 49634 7810 49646
rect 8878 49698 8930 49710
rect 8878 49634 8930 49646
rect 14478 49698 14530 49710
rect 24670 49698 24722 49710
rect 15474 49646 15486 49698
rect 15538 49646 15550 49698
rect 14478 49634 14530 49646
rect 24670 49634 24722 49646
rect 29822 49698 29874 49710
rect 29822 49634 29874 49646
rect 45502 49698 45554 49710
rect 45502 49634 45554 49646
rect 57486 49698 57538 49710
rect 57486 49634 57538 49646
rect 58494 49698 58546 49710
rect 60286 49698 60338 49710
rect 59378 49646 59390 49698
rect 59442 49646 59454 49698
rect 58494 49634 58546 49646
rect 60286 49634 60338 49646
rect 60846 49698 60898 49710
rect 60846 49634 60898 49646
rect 13582 49586 13634 49598
rect 29038 49586 29090 49598
rect 1810 49534 1822 49586
rect 1874 49583 1886 49586
rect 2146 49583 2158 49586
rect 1874 49537 2158 49583
rect 1874 49534 1886 49537
rect 2146 49534 2158 49537
rect 2210 49534 2222 49586
rect 19954 49534 19966 49586
rect 20018 49534 20030 49586
rect 13582 49522 13634 49534
rect 29038 49522 29090 49534
rect 38782 49586 38834 49598
rect 39678 49586 39730 49598
rect 50878 49586 50930 49598
rect 39330 49534 39342 49586
rect 39394 49534 39406 49586
rect 44146 49534 44158 49586
rect 44210 49534 44222 49586
rect 38782 49522 38834 49534
rect 39678 49522 39730 49534
rect 50878 49522 50930 49534
rect 55134 49586 55186 49598
rect 55134 49522 55186 49534
rect 1344 49418 62608 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 62608 49418
rect 1344 49332 62608 49366
rect 11006 49250 11058 49262
rect 11006 49186 11058 49198
rect 21310 49250 21362 49262
rect 21310 49186 21362 49198
rect 21758 49250 21810 49262
rect 34974 49250 35026 49262
rect 30930 49198 30942 49250
rect 30994 49198 31006 49250
rect 21758 49186 21810 49198
rect 34974 49186 35026 49198
rect 42702 49250 42754 49262
rect 42702 49186 42754 49198
rect 48078 49250 48130 49262
rect 48078 49186 48130 49198
rect 51438 49250 51490 49262
rect 51438 49186 51490 49198
rect 54574 49250 54626 49262
rect 54574 49186 54626 49198
rect 4510 49138 4562 49150
rect 4510 49074 4562 49086
rect 5630 49138 5682 49150
rect 5630 49074 5682 49086
rect 6862 49138 6914 49150
rect 10446 49138 10498 49150
rect 21422 49138 21474 49150
rect 10098 49086 10110 49138
rect 10162 49086 10174 49138
rect 11330 49086 11342 49138
rect 11394 49086 11406 49138
rect 6862 49074 6914 49086
rect 10446 49074 10498 49086
rect 21422 49074 21474 49086
rect 27694 49138 27746 49150
rect 35870 49138 35922 49150
rect 32610 49086 32622 49138
rect 32674 49086 32686 49138
rect 27694 49074 27746 49086
rect 35870 49074 35922 49086
rect 37102 49138 37154 49150
rect 37102 49074 37154 49086
rect 44046 49138 44098 49150
rect 47070 49138 47122 49150
rect 45938 49086 45950 49138
rect 46002 49086 46014 49138
rect 44046 49074 44098 49086
rect 47070 49074 47122 49086
rect 49310 49138 49362 49150
rect 58382 49138 58434 49150
rect 52770 49086 52782 49138
rect 52834 49086 52846 49138
rect 49310 49074 49362 49086
rect 58382 49074 58434 49086
rect 59278 49138 59330 49150
rect 60510 49138 60562 49150
rect 59938 49086 59950 49138
rect 60002 49086 60014 49138
rect 59278 49074 59330 49086
rect 60510 49074 60562 49086
rect 4062 49026 4114 49038
rect 2482 48974 2494 49026
rect 2546 48974 2558 49026
rect 4062 48962 4114 48974
rect 4734 49026 4786 49038
rect 4734 48962 4786 48974
rect 5854 49026 5906 49038
rect 10670 49026 10722 49038
rect 12126 49026 12178 49038
rect 7186 48974 7198 49026
rect 7250 48974 7262 49026
rect 11666 48974 11678 49026
rect 11730 48974 11742 49026
rect 5854 48962 5906 48974
rect 10670 48962 10722 48974
rect 12126 48962 12178 48974
rect 14142 49026 14194 49038
rect 14142 48962 14194 48974
rect 14366 49026 14418 49038
rect 14366 48962 14418 48974
rect 15598 49026 15650 49038
rect 20078 49026 20130 49038
rect 17602 48974 17614 49026
rect 17666 48974 17678 49026
rect 18498 48974 18510 49026
rect 18562 48974 18574 49026
rect 19730 48974 19742 49026
rect 19794 48974 19806 49026
rect 15598 48962 15650 48974
rect 20078 48962 20130 48974
rect 22094 49026 22146 49038
rect 28254 49026 28306 49038
rect 30046 49026 30098 49038
rect 35646 49026 35698 49038
rect 22754 48974 22766 49026
rect 22818 48974 22830 49026
rect 24098 48974 24110 49026
rect 24162 48974 24174 49026
rect 24434 48974 24446 49026
rect 24498 48974 24510 49026
rect 29586 48974 29598 49026
rect 29650 48974 29662 49026
rect 31490 48974 31502 49026
rect 31554 48974 31566 49026
rect 32274 48974 32286 49026
rect 32338 48974 32350 49026
rect 34290 48974 34302 49026
rect 34354 48974 34366 49026
rect 22094 48962 22146 48974
rect 28254 48962 28306 48974
rect 30046 48962 30098 48974
rect 35646 48962 35698 48974
rect 36206 49026 36258 49038
rect 36206 48962 36258 48974
rect 36878 49026 36930 49038
rect 36878 48962 36930 48974
rect 37438 49026 37490 49038
rect 38558 49026 38610 49038
rect 42366 49026 42418 49038
rect 46958 49026 47010 49038
rect 38098 48974 38110 49026
rect 38162 48974 38174 49026
rect 39330 48974 39342 49026
rect 39394 48974 39406 49026
rect 40562 48974 40574 49026
rect 40626 48974 40638 49026
rect 43474 48974 43486 49026
rect 43538 48974 43550 49026
rect 37438 48962 37490 48974
rect 38558 48962 38610 48974
rect 42366 48962 42418 48974
rect 46958 48962 47010 48974
rect 47182 49026 47234 49038
rect 58158 49026 58210 49038
rect 48962 48974 48974 49026
rect 49026 48974 49038 49026
rect 49858 48974 49870 49026
rect 49922 48974 49934 49026
rect 50194 48974 50206 49026
rect 50258 48974 50270 49026
rect 50754 48974 50766 49026
rect 50818 48974 50830 49026
rect 52882 48974 52894 49026
rect 52946 48974 52958 49026
rect 53778 48974 53790 49026
rect 53842 48974 53854 49026
rect 47182 48962 47234 48974
rect 58158 48962 58210 48974
rect 59054 49026 59106 49038
rect 59054 48962 59106 48974
rect 59614 49026 59666 49038
rect 59614 48962 59666 48974
rect 60734 49026 60786 49038
rect 61618 48974 61630 49026
rect 61682 48974 61694 49026
rect 60734 48962 60786 48974
rect 2046 48914 2098 48926
rect 3502 48914 3554 48926
rect 17950 48914 18002 48926
rect 2706 48862 2718 48914
rect 2770 48862 2782 48914
rect 7970 48862 7982 48914
rect 8034 48862 8046 48914
rect 11554 48862 11566 48914
rect 11618 48862 11630 48914
rect 12898 48862 12910 48914
rect 12962 48862 12974 48914
rect 14802 48862 14814 48914
rect 14866 48862 14878 48914
rect 15250 48862 15262 48914
rect 15314 48862 15326 48914
rect 16930 48862 16942 48914
rect 16994 48862 17006 48914
rect 2046 48850 2098 48862
rect 3502 48850 3554 48862
rect 17950 48850 18002 48862
rect 20638 48914 20690 48926
rect 20638 48850 20690 48862
rect 22318 48914 22370 48926
rect 28030 48914 28082 48926
rect 36094 48914 36146 48926
rect 24546 48862 24558 48914
rect 24610 48862 24622 48914
rect 26674 48862 26686 48914
rect 26738 48862 26750 48914
rect 30930 48862 30942 48914
rect 30994 48862 31006 48914
rect 34402 48862 34414 48914
rect 34466 48862 34478 48914
rect 22318 48850 22370 48862
rect 28030 48850 28082 48862
rect 36094 48850 36146 48862
rect 37326 48914 37378 48926
rect 45278 48914 45330 48926
rect 47742 48914 47794 48926
rect 39442 48862 39454 48914
rect 39506 48862 39518 48914
rect 41122 48862 41134 48914
rect 41186 48862 41198 48914
rect 43250 48862 43262 48914
rect 43314 48862 43326 48914
rect 45714 48862 45726 48914
rect 45778 48862 45790 48914
rect 37326 48850 37378 48862
rect 45278 48850 45330 48862
rect 47742 48850 47794 48862
rect 48190 48914 48242 48926
rect 48738 48862 48750 48914
rect 48802 48862 48814 48914
rect 50642 48862 50654 48914
rect 50706 48862 50718 48914
rect 54002 48862 54014 48914
rect 54066 48862 54078 48914
rect 56802 48862 56814 48914
rect 56866 48862 56878 48914
rect 48190 48850 48242 48862
rect 1710 48802 1762 48814
rect 1710 48738 1762 48750
rect 3166 48802 3218 48814
rect 3166 48738 3218 48750
rect 4174 48802 4226 48814
rect 11902 48802 11954 48814
rect 5058 48750 5070 48802
rect 5122 48750 5134 48802
rect 6178 48750 6190 48802
rect 6242 48750 6254 48802
rect 4174 48738 4226 48750
rect 11902 48738 11954 48750
rect 12574 48802 12626 48814
rect 15934 48802 15986 48814
rect 13794 48750 13806 48802
rect 13858 48750 13870 48802
rect 12574 48738 12626 48750
rect 15934 48738 15986 48750
rect 25454 48802 25506 48814
rect 35310 48802 35362 48814
rect 28578 48750 28590 48802
rect 28642 48750 28654 48802
rect 25454 48738 25506 48750
rect 35310 48738 35362 48750
rect 37886 48802 37938 48814
rect 37886 48738 37938 48750
rect 38894 48802 38946 48814
rect 38894 48738 38946 48750
rect 44942 48802 44994 48814
rect 44942 48738 44994 48750
rect 47966 48802 48018 48814
rect 47966 48738 48018 48750
rect 51774 48802 51826 48814
rect 51774 48738 51826 48750
rect 54910 48802 54962 48814
rect 54910 48738 54962 48750
rect 55470 48802 55522 48814
rect 61742 48802 61794 48814
rect 57810 48750 57822 48802
rect 57874 48750 57886 48802
rect 58706 48750 58718 48802
rect 58770 48750 58782 48802
rect 61058 48750 61070 48802
rect 61122 48750 61134 48802
rect 55470 48738 55522 48750
rect 61742 48738 61794 48750
rect 1344 48634 62608 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 62608 48634
rect 1344 48548 62608 48582
rect 4174 48466 4226 48478
rect 1698 48414 1710 48466
rect 1762 48414 1774 48466
rect 4174 48402 4226 48414
rect 4958 48466 5010 48478
rect 4958 48402 5010 48414
rect 8094 48466 8146 48478
rect 8094 48402 8146 48414
rect 8766 48466 8818 48478
rect 8766 48402 8818 48414
rect 12798 48466 12850 48478
rect 12798 48402 12850 48414
rect 23326 48466 23378 48478
rect 31614 48466 31666 48478
rect 24322 48414 24334 48466
rect 24386 48414 24398 48466
rect 27234 48414 27246 48466
rect 27298 48414 27310 48466
rect 23326 48402 23378 48414
rect 31614 48402 31666 48414
rect 36542 48466 36594 48478
rect 36542 48402 36594 48414
rect 37662 48466 37714 48478
rect 37662 48402 37714 48414
rect 40126 48466 40178 48478
rect 40126 48402 40178 48414
rect 54350 48466 54402 48478
rect 54350 48402 54402 48414
rect 56702 48466 56754 48478
rect 56702 48402 56754 48414
rect 30046 48354 30098 48366
rect 36654 48354 36706 48366
rect 3042 48302 3054 48354
rect 3106 48302 3118 48354
rect 4610 48302 4622 48354
rect 4674 48302 4686 48354
rect 5730 48302 5742 48354
rect 5794 48302 5806 48354
rect 10658 48302 10670 48354
rect 10722 48302 10734 48354
rect 13122 48302 13134 48354
rect 13186 48302 13198 48354
rect 22194 48302 22206 48354
rect 22258 48302 22270 48354
rect 30594 48302 30606 48354
rect 30658 48302 30670 48354
rect 31042 48302 31054 48354
rect 31106 48302 31118 48354
rect 33170 48302 33182 48354
rect 33234 48302 33246 48354
rect 33730 48302 33742 48354
rect 33794 48302 33806 48354
rect 35298 48302 35310 48354
rect 35362 48302 35374 48354
rect 35746 48302 35758 48354
rect 35810 48302 35822 48354
rect 30046 48290 30098 48302
rect 36654 48290 36706 48302
rect 36766 48354 36818 48366
rect 36766 48290 36818 48302
rect 40014 48354 40066 48366
rect 40014 48290 40066 48302
rect 41582 48354 41634 48366
rect 50878 48354 50930 48366
rect 62078 48354 62130 48366
rect 44146 48302 44158 48354
rect 44210 48302 44222 48354
rect 47730 48302 47742 48354
rect 47794 48302 47806 48354
rect 49970 48302 49982 48354
rect 50034 48302 50046 48354
rect 52434 48302 52446 48354
rect 52498 48302 52510 48354
rect 59602 48302 59614 48354
rect 59666 48302 59678 48354
rect 41582 48290 41634 48302
rect 50878 48290 50930 48302
rect 62078 48290 62130 48302
rect 8318 48242 8370 48254
rect 1922 48190 1934 48242
rect 1986 48190 1998 48242
rect 5282 48190 5294 48242
rect 5346 48190 5358 48242
rect 6290 48190 6302 48242
rect 6354 48190 6366 48242
rect 6738 48190 6750 48242
rect 6802 48190 6814 48242
rect 8318 48178 8370 48190
rect 8990 48242 9042 48254
rect 15374 48242 15426 48254
rect 18062 48242 18114 48254
rect 23774 48242 23826 48254
rect 13570 48190 13582 48242
rect 13634 48190 13646 48242
rect 14690 48190 14702 48242
rect 14754 48190 14766 48242
rect 16594 48190 16606 48242
rect 16658 48190 16670 48242
rect 18274 48190 18286 48242
rect 18338 48190 18350 48242
rect 20066 48190 20078 48242
rect 20130 48190 20142 48242
rect 20514 48190 20526 48242
rect 20578 48190 20590 48242
rect 8990 48178 9042 48190
rect 15374 48178 15426 48190
rect 18062 48178 18114 48190
rect 23774 48178 23826 48190
rect 23998 48242 24050 48254
rect 29038 48242 29090 48254
rect 31278 48242 31330 48254
rect 34862 48242 34914 48254
rect 36430 48242 36482 48254
rect 37438 48242 37490 48254
rect 28578 48190 28590 48242
rect 28642 48190 28654 48242
rect 29810 48190 29822 48242
rect 29874 48190 29886 48242
rect 33058 48190 33070 48242
rect 33122 48190 33134 48242
rect 34290 48190 34302 48242
rect 34354 48190 34366 48242
rect 36082 48190 36094 48242
rect 36146 48190 36158 48242
rect 37202 48190 37214 48242
rect 37266 48190 37278 48242
rect 23998 48178 24050 48190
rect 29038 48178 29090 48190
rect 31278 48178 31330 48190
rect 34862 48178 34914 48190
rect 36430 48178 36482 48190
rect 37438 48178 37490 48190
rect 37774 48242 37826 48254
rect 37774 48178 37826 48190
rect 38110 48242 38162 48254
rect 40350 48242 40402 48254
rect 42590 48242 42642 48254
rect 51214 48242 51266 48254
rect 39554 48190 39566 48242
rect 39618 48190 39630 48242
rect 41122 48190 41134 48242
rect 41186 48190 41198 48242
rect 42018 48190 42030 48242
rect 42082 48190 42094 48242
rect 44594 48190 44606 48242
rect 44658 48190 44670 48242
rect 45490 48190 45502 48242
rect 45554 48190 45566 48242
rect 47058 48190 47070 48242
rect 47122 48190 47134 48242
rect 47618 48190 47630 48242
rect 47682 48190 47694 48242
rect 49410 48190 49422 48242
rect 49474 48190 49486 48242
rect 50642 48190 50654 48242
rect 50706 48190 50718 48242
rect 38110 48178 38162 48190
rect 40350 48178 40402 48190
rect 42590 48178 42642 48190
rect 51214 48178 51266 48190
rect 51438 48242 51490 48254
rect 54574 48242 54626 48254
rect 51762 48190 51774 48242
rect 51826 48190 51838 48242
rect 51438 48178 51490 48190
rect 54574 48178 54626 48190
rect 54798 48242 54850 48254
rect 54798 48178 54850 48190
rect 55246 48242 55298 48254
rect 57934 48242 57986 48254
rect 55458 48190 55470 48242
rect 55522 48190 55534 48242
rect 57138 48190 57150 48242
rect 57202 48190 57214 48242
rect 57698 48190 57710 48242
rect 57762 48190 57774 48242
rect 55246 48178 55298 48190
rect 57934 48178 57986 48190
rect 58270 48242 58322 48254
rect 58270 48178 58322 48190
rect 58494 48242 58546 48254
rect 58494 48178 58546 48190
rect 58942 48242 58994 48254
rect 61842 48190 61854 48242
rect 61906 48190 61918 48242
rect 58942 48178 58994 48190
rect 8878 48130 8930 48142
rect 8878 48066 8930 48078
rect 9550 48130 9602 48142
rect 25342 48130 25394 48142
rect 9762 48078 9774 48130
rect 9826 48078 9838 48130
rect 21074 48078 21086 48130
rect 21138 48078 21150 48130
rect 9550 48066 9602 48078
rect 25342 48066 25394 48078
rect 32622 48130 32674 48142
rect 32622 48066 32674 48078
rect 33854 48130 33906 48142
rect 33854 48066 33906 48078
rect 38446 48130 38498 48142
rect 39230 48130 39282 48142
rect 43038 48130 43090 48142
rect 48862 48130 48914 48142
rect 51326 48130 51378 48142
rect 38770 48078 38782 48130
rect 38834 48078 38846 48130
rect 40002 48078 40014 48130
rect 40066 48078 40078 48130
rect 41458 48078 41470 48130
rect 41522 48078 41534 48130
rect 45602 48078 45614 48130
rect 45666 48078 45678 48130
rect 48066 48078 48078 48130
rect 48130 48078 48142 48130
rect 49858 48078 49870 48130
rect 49922 48078 49934 48130
rect 38446 48066 38498 48078
rect 39230 48066 39282 48078
rect 43038 48066 43090 48078
rect 48862 48066 48914 48078
rect 51326 48066 51378 48078
rect 54686 48130 54738 48142
rect 54686 48066 54738 48078
rect 57822 48130 57874 48142
rect 57822 48066 57874 48078
rect 58382 48130 58434 48142
rect 58382 48066 58434 48078
rect 12462 48018 12514 48030
rect 25902 48018 25954 48030
rect 61518 48018 61570 48030
rect 16706 47966 16718 48018
rect 16770 47966 16782 48018
rect 28914 47966 28926 48018
rect 28978 47966 28990 48018
rect 46274 47966 46286 48018
rect 46338 47966 46350 48018
rect 56018 47966 56030 48018
rect 56082 47966 56094 48018
rect 57362 47966 57374 48018
rect 57426 47966 57438 48018
rect 12462 47954 12514 47966
rect 25902 47954 25954 47966
rect 61518 47954 61570 47966
rect 1344 47850 62608 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 62608 47850
rect 1344 47764 62608 47798
rect 8542 47682 8594 47694
rect 8542 47618 8594 47630
rect 24110 47682 24162 47694
rect 24110 47618 24162 47630
rect 26574 47682 26626 47694
rect 46062 47682 46114 47694
rect 30930 47630 30942 47682
rect 30994 47630 31006 47682
rect 33618 47630 33630 47682
rect 33682 47630 33694 47682
rect 35634 47630 35646 47682
rect 35698 47630 35710 47682
rect 41570 47630 41582 47682
rect 41634 47630 41646 47682
rect 26574 47618 26626 47630
rect 46062 47618 46114 47630
rect 51774 47682 51826 47694
rect 51774 47618 51826 47630
rect 53566 47682 53618 47694
rect 61966 47682 62018 47694
rect 59266 47630 59278 47682
rect 59330 47630 59342 47682
rect 53566 47618 53618 47630
rect 61966 47618 62018 47630
rect 16158 47570 16210 47582
rect 4610 47518 4622 47570
rect 4674 47518 4686 47570
rect 9202 47518 9214 47570
rect 9266 47518 9278 47570
rect 16158 47506 16210 47518
rect 19854 47570 19906 47582
rect 19854 47506 19906 47518
rect 22542 47570 22594 47582
rect 22542 47506 22594 47518
rect 23662 47570 23714 47582
rect 51326 47570 51378 47582
rect 53678 47570 53730 47582
rect 27794 47518 27806 47570
rect 27858 47518 27870 47570
rect 37986 47518 37998 47570
rect 38050 47518 38062 47570
rect 43026 47518 43038 47570
rect 43090 47518 43102 47570
rect 53106 47518 53118 47570
rect 53170 47518 53182 47570
rect 23662 47506 23714 47518
rect 51326 47506 51378 47518
rect 53678 47506 53730 47518
rect 60958 47570 61010 47582
rect 60958 47506 61010 47518
rect 11230 47458 11282 47470
rect 16046 47458 16098 47470
rect 19966 47458 20018 47470
rect 1698 47406 1710 47458
rect 1762 47406 1774 47458
rect 9314 47406 9326 47458
rect 9378 47406 9390 47458
rect 10322 47406 10334 47458
rect 10386 47406 10398 47458
rect 10546 47406 10558 47458
rect 10610 47406 10622 47458
rect 12002 47406 12014 47458
rect 12066 47406 12078 47458
rect 12674 47406 12686 47458
rect 12738 47406 12750 47458
rect 14018 47406 14030 47458
rect 14082 47406 14094 47458
rect 14242 47406 14254 47458
rect 14306 47406 14318 47458
rect 15474 47406 15486 47458
rect 15538 47406 15550 47458
rect 16482 47406 16494 47458
rect 16546 47406 16558 47458
rect 17490 47406 17502 47458
rect 17554 47406 17566 47458
rect 11230 47394 11282 47406
rect 16046 47394 16098 47406
rect 19966 47394 20018 47406
rect 20302 47458 20354 47470
rect 24446 47458 24498 47470
rect 35086 47458 35138 47470
rect 43822 47458 43874 47470
rect 51438 47458 51490 47470
rect 57598 47458 57650 47470
rect 58942 47458 58994 47470
rect 60622 47458 60674 47470
rect 21298 47406 21310 47458
rect 21362 47406 21374 47458
rect 25778 47406 25790 47458
rect 25842 47406 25854 47458
rect 29362 47406 29374 47458
rect 29426 47406 29438 47458
rect 30594 47406 30606 47458
rect 30658 47406 30670 47458
rect 31490 47406 31502 47458
rect 31554 47406 31566 47458
rect 33282 47406 33294 47458
rect 33346 47406 33358 47458
rect 34290 47406 34302 47458
rect 34354 47406 34366 47458
rect 35298 47406 35310 47458
rect 35362 47406 35374 47458
rect 35858 47406 35870 47458
rect 35922 47406 35934 47458
rect 37650 47406 37662 47458
rect 37714 47406 37726 47458
rect 41794 47406 41806 47458
rect 41858 47406 41870 47458
rect 45826 47406 45838 47458
rect 45890 47406 45902 47458
rect 47506 47406 47518 47458
rect 47570 47406 47582 47458
rect 48850 47406 48862 47458
rect 48914 47406 48926 47458
rect 49522 47406 49534 47458
rect 49586 47406 49598 47458
rect 52098 47406 52110 47458
rect 52162 47406 52174 47458
rect 55010 47406 55022 47458
rect 55074 47406 55086 47458
rect 55458 47406 55470 47458
rect 55522 47406 55534 47458
rect 56354 47406 56366 47458
rect 56418 47406 56430 47458
rect 56802 47406 56814 47458
rect 56866 47406 56878 47458
rect 58482 47406 58494 47458
rect 58546 47406 58558 47458
rect 59714 47406 59726 47458
rect 59778 47406 59790 47458
rect 20302 47394 20354 47406
rect 24446 47394 24498 47406
rect 35086 47394 35138 47406
rect 43822 47394 43874 47406
rect 51438 47394 51490 47406
rect 57598 47394 57650 47406
rect 58942 47394 58994 47406
rect 60622 47394 60674 47406
rect 60734 47458 60786 47470
rect 60734 47394 60786 47406
rect 4958 47346 5010 47358
rect 13582 47346 13634 47358
rect 16270 47346 16322 47358
rect 18062 47346 18114 47358
rect 26910 47346 26962 47358
rect 28254 47346 28306 47358
rect 2482 47294 2494 47346
rect 2546 47294 2558 47346
rect 6514 47294 6526 47346
rect 6578 47294 6590 47346
rect 9202 47294 9214 47346
rect 9266 47294 9278 47346
rect 12786 47294 12798 47346
rect 12850 47294 12862 47346
rect 14690 47294 14702 47346
rect 14754 47294 14766 47346
rect 15362 47294 15374 47346
rect 15426 47294 15438 47346
rect 16594 47294 16606 47346
rect 16658 47294 16670 47346
rect 21410 47294 21422 47346
rect 21474 47294 21486 47346
rect 21970 47294 21982 47346
rect 22034 47294 22046 47346
rect 23314 47294 23326 47346
rect 23378 47294 23390 47346
rect 24770 47294 24782 47346
rect 24834 47294 24846 47346
rect 24994 47294 25006 47346
rect 25058 47294 25070 47346
rect 26002 47294 26014 47346
rect 26066 47294 26078 47346
rect 28130 47294 28142 47346
rect 28194 47294 28206 47346
rect 4958 47282 5010 47294
rect 13582 47282 13634 47294
rect 16270 47282 16322 47294
rect 18062 47282 18114 47294
rect 26910 47282 26962 47294
rect 28254 47282 28306 47294
rect 28366 47346 28418 47358
rect 28366 47282 28418 47294
rect 28590 47346 28642 47358
rect 33070 47346 33122 47358
rect 31938 47294 31950 47346
rect 32002 47294 32014 47346
rect 28590 47282 28642 47294
rect 33070 47282 33122 47294
rect 34078 47346 34130 47358
rect 34078 47282 34130 47294
rect 37214 47346 37266 47358
rect 42590 47346 42642 47358
rect 39106 47294 39118 47346
rect 39170 47294 39182 47346
rect 37214 47282 37266 47294
rect 42590 47282 42642 47294
rect 42702 47346 42754 47358
rect 43486 47346 43538 47358
rect 43362 47294 43374 47346
rect 43426 47294 43438 47346
rect 42702 47282 42754 47294
rect 43486 47282 43538 47294
rect 43598 47346 43650 47358
rect 49982 47346 50034 47358
rect 46162 47294 46174 47346
rect 46226 47294 46238 47346
rect 43598 47282 43650 47294
rect 49982 47282 50034 47294
rect 50094 47346 50146 47358
rect 50094 47282 50146 47294
rect 50206 47346 50258 47358
rect 51102 47346 51154 47358
rect 62190 47346 62242 47358
rect 50866 47294 50878 47346
rect 50930 47294 50942 47346
rect 55794 47294 55806 47346
rect 55858 47294 55870 47346
rect 56914 47294 56926 47346
rect 56978 47294 56990 47346
rect 50206 47282 50258 47294
rect 51102 47282 51154 47294
rect 62190 47282 62242 47294
rect 5070 47234 5122 47246
rect 5070 47170 5122 47182
rect 10894 47234 10946 47246
rect 10894 47170 10946 47182
rect 11118 47234 11170 47246
rect 13470 47234 13522 47246
rect 11890 47182 11902 47234
rect 11954 47182 11966 47234
rect 11118 47170 11170 47182
rect 13470 47170 13522 47182
rect 22990 47234 23042 47246
rect 22990 47170 23042 47182
rect 27582 47234 27634 47246
rect 36318 47234 36370 47246
rect 42366 47234 42418 47246
rect 35410 47182 35422 47234
rect 35474 47182 35486 47234
rect 40562 47182 40574 47234
rect 40626 47182 40638 47234
rect 27582 47170 27634 47182
rect 36318 47170 36370 47182
rect 42366 47170 42418 47182
rect 44270 47234 44322 47246
rect 45166 47234 45218 47246
rect 44818 47182 44830 47234
rect 44882 47182 44894 47234
rect 44270 47170 44322 47182
rect 45166 47170 45218 47182
rect 50318 47234 50370 47246
rect 50318 47170 50370 47182
rect 51214 47234 51266 47246
rect 51214 47170 51266 47182
rect 51886 47234 51938 47246
rect 51886 47170 51938 47182
rect 52670 47234 52722 47246
rect 52670 47170 52722 47182
rect 57934 47234 57986 47246
rect 57934 47170 57986 47182
rect 60622 47234 60674 47246
rect 61618 47182 61630 47234
rect 61682 47182 61694 47234
rect 60622 47170 60674 47182
rect 1344 47066 62608 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 62608 47066
rect 1344 46980 62608 47014
rect 5294 46898 5346 46910
rect 5294 46834 5346 46846
rect 8542 46898 8594 46910
rect 8542 46834 8594 46846
rect 12798 46898 12850 46910
rect 12798 46834 12850 46846
rect 13022 46898 13074 46910
rect 13022 46834 13074 46846
rect 13134 46898 13186 46910
rect 13134 46834 13186 46846
rect 13246 46898 13298 46910
rect 13246 46834 13298 46846
rect 18622 46898 18674 46910
rect 18622 46834 18674 46846
rect 27470 46898 27522 46910
rect 42254 46898 42306 46910
rect 38210 46846 38222 46898
rect 38274 46846 38286 46898
rect 27470 46834 27522 46846
rect 42254 46834 42306 46846
rect 43822 46898 43874 46910
rect 43822 46834 43874 46846
rect 44046 46898 44098 46910
rect 44046 46834 44098 46846
rect 45726 46898 45778 46910
rect 45726 46834 45778 46846
rect 45838 46898 45890 46910
rect 45838 46834 45890 46846
rect 45950 46898 46002 46910
rect 45950 46834 46002 46846
rect 46398 46898 46450 46910
rect 50430 46898 50482 46910
rect 49298 46846 49310 46898
rect 49362 46846 49374 46898
rect 46398 46834 46450 46846
rect 50430 46834 50482 46846
rect 53342 46898 53394 46910
rect 53342 46834 53394 46846
rect 53678 46898 53730 46910
rect 53678 46834 53730 46846
rect 2270 46786 2322 46798
rect 2270 46722 2322 46734
rect 3614 46786 3666 46798
rect 3614 46722 3666 46734
rect 3950 46786 4002 46798
rect 6862 46786 6914 46798
rect 6626 46734 6638 46786
rect 6690 46734 6702 46786
rect 3950 46722 4002 46734
rect 6862 46722 6914 46734
rect 8430 46786 8482 46798
rect 8430 46722 8482 46734
rect 10446 46786 10498 46798
rect 10446 46722 10498 46734
rect 10670 46786 10722 46798
rect 10670 46722 10722 46734
rect 10782 46786 10834 46798
rect 10782 46722 10834 46734
rect 11790 46786 11842 46798
rect 22878 46786 22930 46798
rect 24558 46786 24610 46798
rect 32510 46786 32562 46798
rect 14466 46734 14478 46786
rect 14530 46734 14542 46786
rect 15362 46734 15374 46786
rect 15426 46734 15438 46786
rect 15922 46734 15934 46786
rect 15986 46734 15998 46786
rect 17714 46734 17726 46786
rect 17778 46734 17790 46786
rect 17938 46734 17950 46786
rect 18002 46734 18014 46786
rect 19730 46734 19742 46786
rect 19794 46734 19806 46786
rect 23986 46734 23998 46786
rect 24050 46734 24062 46786
rect 25554 46734 25566 46786
rect 25618 46734 25630 46786
rect 28802 46734 28814 46786
rect 28866 46734 28878 46786
rect 31602 46734 31614 46786
rect 31666 46734 31678 46786
rect 32162 46734 32174 46786
rect 32226 46734 32238 46786
rect 11790 46722 11842 46734
rect 22878 46722 22930 46734
rect 24558 46722 24610 46734
rect 32510 46722 32562 46734
rect 33406 46786 33458 46798
rect 33406 46722 33458 46734
rect 33854 46786 33906 46798
rect 33854 46722 33906 46734
rect 40910 46786 40962 46798
rect 45614 46786 45666 46798
rect 48078 46786 48130 46798
rect 42802 46734 42814 46786
rect 42866 46734 42878 46786
rect 43362 46734 43374 46786
rect 43426 46734 43438 46786
rect 45378 46734 45390 46786
rect 45442 46734 45454 46786
rect 47506 46734 47518 46786
rect 47570 46734 47582 46786
rect 40910 46722 40962 46734
rect 45614 46722 45666 46734
rect 48078 46722 48130 46734
rect 48190 46786 48242 46798
rect 53902 46786 53954 46798
rect 56702 46786 56754 46798
rect 49410 46734 49422 46786
rect 49474 46734 49486 46786
rect 49858 46734 49870 46786
rect 49922 46734 49934 46786
rect 51538 46734 51550 46786
rect 51602 46734 51614 46786
rect 54450 46734 54462 46786
rect 54514 46734 54526 46786
rect 48190 46722 48242 46734
rect 53902 46722 53954 46734
rect 56702 46722 56754 46734
rect 56814 46786 56866 46798
rect 57474 46734 57486 46786
rect 57538 46734 57550 46786
rect 56814 46722 56866 46734
rect 2494 46674 2546 46686
rect 2494 46610 2546 46622
rect 2718 46674 2770 46686
rect 2718 46610 2770 46622
rect 3838 46674 3890 46686
rect 8318 46674 8370 46686
rect 6066 46622 6078 46674
rect 6130 46622 6142 46674
rect 7298 46622 7310 46674
rect 7362 46622 7374 46674
rect 3838 46610 3890 46622
rect 8318 46610 8370 46622
rect 9550 46674 9602 46686
rect 9550 46610 9602 46622
rect 9774 46674 9826 46686
rect 16158 46674 16210 46686
rect 22766 46674 22818 46686
rect 13794 46622 13806 46674
rect 13858 46622 13870 46674
rect 14690 46622 14702 46674
rect 14754 46622 14766 46674
rect 19282 46622 19294 46674
rect 19346 46622 19358 46674
rect 21074 46622 21086 46674
rect 21138 46622 21150 46674
rect 9774 46610 9826 46622
rect 16158 46610 16210 46622
rect 22766 46610 22818 46622
rect 22990 46674 23042 46686
rect 33630 46674 33682 46686
rect 42590 46674 42642 46686
rect 44830 46674 44882 46686
rect 23314 46622 23326 46674
rect 23378 46622 23390 46674
rect 23762 46622 23774 46674
rect 23826 46622 23838 46674
rect 24322 46622 24334 46674
rect 24386 46622 24398 46674
rect 27794 46622 27806 46674
rect 27858 46622 27870 46674
rect 28578 46622 28590 46674
rect 28642 46622 28654 46674
rect 29698 46622 29710 46674
rect 29762 46622 29774 46674
rect 29922 46622 29934 46674
rect 29986 46622 29998 46674
rect 31378 46622 31390 46674
rect 31442 46622 31454 46674
rect 34178 46622 34190 46674
rect 34242 46622 34254 46674
rect 40002 46622 40014 46674
rect 40066 46622 40078 46674
rect 44370 46622 44382 46674
rect 44434 46622 44446 46674
rect 22990 46610 23042 46622
rect 33630 46610 33682 46622
rect 42590 46610 42642 46622
rect 44830 46610 44882 46622
rect 46734 46674 46786 46686
rect 48974 46674 49026 46686
rect 55246 46674 55298 46686
rect 61518 46674 61570 46686
rect 47282 46622 47294 46674
rect 47346 46622 47358 46674
rect 50530 46622 50542 46674
rect 50594 46622 50606 46674
rect 54786 46622 54798 46674
rect 54850 46622 54862 46674
rect 55682 46622 55694 46674
rect 55746 46622 55758 46674
rect 58146 46622 58158 46674
rect 58210 46622 58222 46674
rect 59042 46622 59054 46674
rect 59106 46622 59118 46674
rect 60274 46622 60286 46674
rect 60338 46622 60350 46674
rect 46734 46610 46786 46622
rect 48974 46610 49026 46622
rect 55246 46610 55298 46622
rect 61518 46610 61570 46622
rect 61966 46674 62018 46686
rect 61966 46610 62018 46622
rect 62190 46674 62242 46686
rect 62190 46610 62242 46622
rect 1934 46562 1986 46574
rect 1934 46498 1986 46510
rect 2606 46562 2658 46574
rect 2606 46498 2658 46510
rect 4510 46562 4562 46574
rect 8766 46562 8818 46574
rect 16270 46562 16322 46574
rect 16830 46562 16882 46574
rect 4834 46510 4846 46562
rect 4898 46510 4910 46562
rect 6290 46510 6302 46562
rect 6354 46510 6366 46562
rect 14018 46510 14030 46562
rect 14082 46510 14094 46562
rect 16482 46510 16494 46562
rect 16546 46510 16558 46562
rect 4510 46498 4562 46510
rect 8766 46498 8818 46510
rect 16270 46498 16322 46510
rect 16830 46498 16882 46510
rect 18286 46562 18338 46574
rect 24670 46562 24722 46574
rect 33742 46562 33794 46574
rect 43934 46562 43986 46574
rect 61294 46562 61346 46574
rect 21298 46510 21310 46562
rect 21362 46510 21374 46562
rect 28130 46510 28142 46562
rect 28194 46510 28206 46562
rect 34962 46510 34974 46562
rect 35026 46510 35038 46562
rect 37090 46510 37102 46562
rect 37154 46510 37166 46562
rect 54338 46510 54350 46562
rect 54402 46510 54414 46562
rect 57250 46510 57262 46562
rect 57314 46510 57326 46562
rect 18286 46498 18338 46510
rect 24670 46498 24722 46510
rect 33742 46498 33794 46510
rect 43934 46498 43986 46510
rect 61294 46498 61346 46510
rect 61742 46562 61794 46574
rect 61742 46498 61794 46510
rect 3166 46450 3218 46462
rect 3166 46386 3218 46398
rect 3390 46450 3442 46462
rect 3390 46386 3442 46398
rect 8990 46450 9042 46462
rect 11006 46450 11058 46462
rect 10098 46398 10110 46450
rect 10162 46398 10174 46450
rect 8990 46386 9042 46398
rect 11006 46386 11058 46398
rect 11230 46450 11282 46462
rect 11230 46386 11282 46398
rect 12014 46450 12066 46462
rect 12014 46386 12066 46398
rect 12350 46450 12402 46462
rect 41134 46450 41186 46462
rect 21410 46398 21422 46450
rect 21474 46398 21486 46450
rect 12350 46386 12402 46398
rect 41134 46386 41186 46398
rect 41470 46450 41522 46462
rect 41470 46386 41522 46398
rect 48078 46450 48130 46462
rect 48078 46386 48130 46398
rect 53566 46450 53618 46462
rect 53566 46386 53618 46398
rect 56702 46450 56754 46462
rect 56702 46386 56754 46398
rect 1344 46282 62608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 62608 46282
rect 1344 46196 62608 46230
rect 7422 46114 7474 46126
rect 7422 46050 7474 46062
rect 9774 46114 9826 46126
rect 9774 46050 9826 46062
rect 9998 46114 10050 46126
rect 18174 46114 18226 46126
rect 28254 46114 28306 46126
rect 37102 46114 37154 46126
rect 11778 46062 11790 46114
rect 11842 46062 11854 46114
rect 24770 46062 24782 46114
rect 24834 46062 24846 46114
rect 28578 46062 28590 46114
rect 28642 46062 28654 46114
rect 9998 46050 10050 46062
rect 18174 46050 18226 46062
rect 28254 46050 28306 46062
rect 37102 46050 37154 46062
rect 39678 46114 39730 46126
rect 46050 46062 46062 46114
rect 46114 46062 46126 46114
rect 55682 46062 55694 46114
rect 55746 46062 55758 46114
rect 39678 46050 39730 46062
rect 11342 46002 11394 46014
rect 28030 46002 28082 46014
rect 5730 45950 5742 46002
rect 5794 45950 5806 46002
rect 8642 45950 8654 46002
rect 8706 45950 8718 46002
rect 18946 45950 18958 46002
rect 19010 45950 19022 46002
rect 20066 45950 20078 46002
rect 20130 45950 20142 46002
rect 24210 45950 24222 46002
rect 24274 45950 24286 46002
rect 11342 45938 11394 45950
rect 28030 45938 28082 45950
rect 29598 46002 29650 46014
rect 29598 45938 29650 45950
rect 30382 46002 30434 46014
rect 30382 45938 30434 45950
rect 31278 46002 31330 46014
rect 51550 46002 51602 46014
rect 60622 46002 60674 46014
rect 44258 45950 44270 46002
rect 44322 45950 44334 46002
rect 44930 45950 44942 46002
rect 44994 45950 45006 46002
rect 47954 45950 47966 46002
rect 48018 45950 48030 46002
rect 55458 45950 55470 46002
rect 55522 45950 55534 46002
rect 31278 45938 31330 45950
rect 51550 45938 51602 45950
rect 60622 45938 60674 45950
rect 5182 45890 5234 45902
rect 10446 45890 10498 45902
rect 6066 45838 6078 45890
rect 6130 45838 6142 45890
rect 8530 45838 8542 45890
rect 8594 45838 8606 45890
rect 9202 45838 9214 45890
rect 9266 45838 9278 45890
rect 5182 45826 5234 45838
rect 10446 45826 10498 45838
rect 11230 45890 11282 45902
rect 12350 45890 12402 45902
rect 18622 45890 18674 45902
rect 25790 45890 25842 45902
rect 11778 45838 11790 45890
rect 11842 45838 11854 45890
rect 13458 45838 13470 45890
rect 13522 45838 13534 45890
rect 14354 45838 14366 45890
rect 14418 45838 14430 45890
rect 15138 45838 15150 45890
rect 15202 45838 15214 45890
rect 18834 45838 18846 45890
rect 18898 45838 18910 45890
rect 19730 45838 19742 45890
rect 19794 45838 19806 45890
rect 21410 45838 21422 45890
rect 21474 45838 21486 45890
rect 24546 45838 24558 45890
rect 24610 45838 24622 45890
rect 11230 45826 11282 45838
rect 12350 45826 12402 45838
rect 18622 45826 18674 45838
rect 25790 45826 25842 45838
rect 26014 45890 26066 45902
rect 26014 45826 26066 45838
rect 26350 45890 26402 45902
rect 26350 45826 26402 45838
rect 26798 45890 26850 45902
rect 26798 45826 26850 45838
rect 27022 45890 27074 45902
rect 27022 45826 27074 45838
rect 27470 45890 27522 45902
rect 29486 45890 29538 45902
rect 29138 45838 29150 45890
rect 29202 45838 29214 45890
rect 27470 45826 27522 45838
rect 29486 45826 29538 45838
rect 29710 45890 29762 45902
rect 29710 45826 29762 45838
rect 31166 45890 31218 45902
rect 31166 45826 31218 45838
rect 35534 45890 35586 45902
rect 50542 45890 50594 45902
rect 40226 45838 40238 45890
rect 40290 45838 40302 45890
rect 41346 45838 41358 45890
rect 41410 45838 41422 45890
rect 46834 45838 46846 45890
rect 46898 45838 46910 45890
rect 47842 45838 47854 45890
rect 47906 45838 47918 45890
rect 50082 45838 50094 45890
rect 50146 45838 50158 45890
rect 35534 45826 35586 45838
rect 50542 45826 50594 45838
rect 51326 45890 51378 45902
rect 51326 45826 51378 45838
rect 53118 45890 53170 45902
rect 60510 45890 60562 45902
rect 61966 45890 62018 45902
rect 55570 45838 55582 45890
rect 55634 45838 55646 45890
rect 56466 45838 56478 45890
rect 56530 45838 56542 45890
rect 61282 45838 61294 45890
rect 61346 45838 61358 45890
rect 53118 45826 53170 45838
rect 60510 45826 60562 45838
rect 61966 45826 62018 45838
rect 62190 45890 62242 45902
rect 62190 45826 62242 45838
rect 4510 45778 4562 45790
rect 3042 45726 3054 45778
rect 3106 45726 3118 45778
rect 4510 45714 4562 45726
rect 4734 45778 4786 45790
rect 10558 45778 10610 45790
rect 12910 45778 12962 45790
rect 25342 45778 25394 45790
rect 6738 45726 6750 45778
rect 6802 45726 6814 45778
rect 7186 45726 7198 45778
rect 7250 45726 7262 45778
rect 8642 45726 8654 45778
rect 8706 45726 8718 45778
rect 11442 45726 11454 45778
rect 11506 45726 11518 45778
rect 14242 45726 14254 45778
rect 14306 45726 14318 45778
rect 16706 45726 16718 45778
rect 16770 45726 16782 45778
rect 22082 45726 22094 45778
rect 22146 45726 22158 45778
rect 25106 45726 25118 45778
rect 25170 45726 25182 45778
rect 4734 45714 4786 45726
rect 10558 45714 10610 45726
rect 12910 45714 12962 45726
rect 25342 45714 25394 45726
rect 26574 45778 26626 45790
rect 26574 45714 26626 45726
rect 30942 45778 30994 45790
rect 30942 45714 30994 45726
rect 33966 45778 34018 45790
rect 45390 45778 45442 45790
rect 60846 45778 60898 45790
rect 34850 45726 34862 45778
rect 34914 45726 34926 45778
rect 35186 45726 35198 45778
rect 35250 45726 35262 45778
rect 38210 45726 38222 45778
rect 38274 45726 38286 45778
rect 40338 45726 40350 45778
rect 40402 45726 40414 45778
rect 42130 45726 42142 45778
rect 42194 45726 42206 45778
rect 46610 45726 46622 45778
rect 46674 45726 46686 45778
rect 49746 45726 49758 45778
rect 49810 45726 49822 45778
rect 53330 45726 53342 45778
rect 53394 45726 53406 45778
rect 53890 45726 53902 45778
rect 53954 45726 53966 45778
rect 57026 45726 57038 45778
rect 57090 45726 57102 45778
rect 58706 45726 58718 45778
rect 58770 45726 58782 45778
rect 33966 45714 34018 45726
rect 45390 45714 45442 45726
rect 60846 45714 60898 45726
rect 1822 45666 1874 45678
rect 1822 45602 1874 45614
rect 4286 45666 4338 45678
rect 4286 45602 4338 45614
rect 4846 45666 4898 45678
rect 4846 45602 4898 45614
rect 7758 45666 7810 45678
rect 7758 45602 7810 45614
rect 9662 45666 9714 45678
rect 9662 45602 9714 45614
rect 20862 45666 20914 45678
rect 20862 45602 20914 45614
rect 24558 45666 24610 45678
rect 24558 45602 24610 45614
rect 26014 45666 26066 45678
rect 26014 45602 26066 45614
rect 26686 45666 26738 45678
rect 26686 45602 26738 45614
rect 27582 45666 27634 45678
rect 27582 45602 27634 45614
rect 27806 45666 27858 45678
rect 27806 45602 27858 45614
rect 31390 45666 31442 45678
rect 33518 45666 33570 45678
rect 32386 45614 32398 45666
rect 32450 45614 32462 45666
rect 31390 45602 31442 45614
rect 33518 45602 33570 45614
rect 34302 45666 34354 45678
rect 34302 45602 34354 45614
rect 35870 45666 35922 45678
rect 35870 45602 35922 45614
rect 36542 45666 36594 45678
rect 36542 45602 36594 45614
rect 39342 45666 39394 45678
rect 39342 45602 39394 45614
rect 41134 45666 41186 45678
rect 41134 45602 41186 45614
rect 50878 45666 50930 45678
rect 52782 45666 52834 45678
rect 51874 45614 51886 45666
rect 51938 45614 51950 45666
rect 50878 45602 50930 45614
rect 52782 45602 52834 45614
rect 59838 45666 59890 45678
rect 59838 45602 59890 45614
rect 60734 45666 60786 45678
rect 61618 45614 61630 45666
rect 61682 45614 61694 45666
rect 60734 45602 60786 45614
rect 1344 45498 62608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 62608 45498
rect 1344 45412 62608 45446
rect 4174 45330 4226 45342
rect 4174 45266 4226 45278
rect 7086 45330 7138 45342
rect 7086 45266 7138 45278
rect 7310 45330 7362 45342
rect 7310 45266 7362 45278
rect 8542 45330 8594 45342
rect 8542 45266 8594 45278
rect 10670 45330 10722 45342
rect 10670 45266 10722 45278
rect 11230 45330 11282 45342
rect 11230 45266 11282 45278
rect 12798 45330 12850 45342
rect 12798 45266 12850 45278
rect 17390 45330 17442 45342
rect 17390 45266 17442 45278
rect 17614 45330 17666 45342
rect 17614 45266 17666 45278
rect 26350 45330 26402 45342
rect 40910 45330 40962 45342
rect 46846 45330 46898 45342
rect 35186 45278 35198 45330
rect 35250 45278 35262 45330
rect 40226 45278 40238 45330
rect 40290 45278 40302 45330
rect 45714 45278 45726 45330
rect 45778 45278 45790 45330
rect 26350 45266 26402 45278
rect 40910 45266 40962 45278
rect 46846 45266 46898 45278
rect 53790 45330 53842 45342
rect 53790 45266 53842 45278
rect 7422 45218 7474 45230
rect 2594 45166 2606 45218
rect 2658 45166 2670 45218
rect 3154 45166 3166 45218
rect 3218 45166 3230 45218
rect 6626 45166 6638 45218
rect 6690 45166 6702 45218
rect 7422 45154 7474 45166
rect 8206 45218 8258 45230
rect 8206 45154 8258 45166
rect 10558 45218 10610 45230
rect 10558 45154 10610 45166
rect 10782 45218 10834 45230
rect 17726 45218 17778 45230
rect 23886 45218 23938 45230
rect 35646 45218 35698 45230
rect 41694 45218 41746 45230
rect 43822 45218 43874 45230
rect 47630 45218 47682 45230
rect 12226 45166 12238 45218
rect 12290 45166 12302 45218
rect 21746 45166 21758 45218
rect 21810 45166 21822 45218
rect 24098 45166 24110 45218
rect 24162 45166 24174 45218
rect 28130 45166 28142 45218
rect 28194 45166 28206 45218
rect 36530 45166 36542 45218
rect 36594 45166 36606 45218
rect 43250 45166 43262 45218
rect 43314 45166 43326 45218
rect 43922 45166 43934 45218
rect 43986 45166 43998 45218
rect 10782 45154 10834 45166
rect 17726 45154 17778 45166
rect 23886 45154 23938 45166
rect 35646 45154 35698 45166
rect 41694 45154 41746 45166
rect 43822 45154 43874 45166
rect 47630 45154 47682 45166
rect 48862 45218 48914 45230
rect 53678 45218 53730 45230
rect 49970 45166 49982 45218
rect 50034 45166 50046 45218
rect 55906 45166 55918 45218
rect 55970 45166 55982 45218
rect 56914 45166 56926 45218
rect 56978 45166 56990 45218
rect 61618 45166 61630 45218
rect 61682 45166 61694 45218
rect 48862 45154 48914 45166
rect 53678 45154 53730 45166
rect 8430 45106 8482 45118
rect 2370 45054 2382 45106
rect 2434 45054 2446 45106
rect 3042 45054 3054 45106
rect 3106 45054 3118 45106
rect 5282 45054 5294 45106
rect 5346 45054 5358 45106
rect 6290 45054 6302 45106
rect 6354 45054 6366 45106
rect 7858 45054 7870 45106
rect 7922 45054 7934 45106
rect 8430 45042 8482 45054
rect 8766 45106 8818 45118
rect 8766 45042 8818 45054
rect 9550 45106 9602 45118
rect 9550 45042 9602 45054
rect 11566 45106 11618 45118
rect 15374 45106 15426 45118
rect 20638 45106 20690 45118
rect 22878 45106 22930 45118
rect 12338 45054 12350 45106
rect 12402 45054 12414 45106
rect 13010 45054 13022 45106
rect 13074 45054 13086 45106
rect 13570 45054 13582 45106
rect 13634 45054 13646 45106
rect 14690 45054 14702 45106
rect 14754 45054 14766 45106
rect 16258 45054 16270 45106
rect 16322 45054 16334 45106
rect 18050 45054 18062 45106
rect 18114 45054 18126 45106
rect 20178 45054 20190 45106
rect 20242 45054 20254 45106
rect 21074 45054 21086 45106
rect 21138 45054 21150 45106
rect 11566 45042 11618 45054
rect 15374 45042 15426 45054
rect 20638 45042 20690 45054
rect 22878 45042 22930 45054
rect 23214 45106 23266 45118
rect 23214 45042 23266 45054
rect 23438 45106 23490 45118
rect 23438 45042 23490 45054
rect 23998 45106 24050 45118
rect 33742 45106 33794 45118
rect 43710 45106 43762 45118
rect 47182 45106 47234 45118
rect 24658 45054 24670 45106
rect 24722 45054 24734 45106
rect 26002 45054 26014 45106
rect 26066 45054 26078 45106
rect 29250 45054 29262 45106
rect 29314 45054 29326 45106
rect 33394 45054 33406 45106
rect 33458 45054 33470 45106
rect 37202 45054 37214 45106
rect 37266 45054 37278 45106
rect 38098 45054 38110 45106
rect 38162 45054 38174 45106
rect 39218 45054 39230 45106
rect 39282 45054 39294 45106
rect 41122 45054 41134 45106
rect 41186 45054 41198 45106
rect 42130 45054 42142 45106
rect 42194 45054 42206 45106
rect 43026 45054 43038 45106
rect 43090 45054 43102 45106
rect 44482 45054 44494 45106
rect 44546 45054 44558 45106
rect 23998 45042 24050 45054
rect 33742 45042 33794 45054
rect 43710 45042 43762 45054
rect 47182 45042 47234 45054
rect 47742 45106 47794 45118
rect 47742 45042 47794 45054
rect 48974 45106 49026 45118
rect 54014 45106 54066 45118
rect 50306 45054 50318 45106
rect 50370 45054 50382 45106
rect 51202 45054 51214 45106
rect 51266 45054 51278 45106
rect 53330 45054 53342 45106
rect 53394 45054 53406 45106
rect 54786 45054 54798 45106
rect 54850 45054 54862 45106
rect 55570 45054 55582 45106
rect 55634 45054 55646 45106
rect 60162 45054 60174 45106
rect 60226 45054 60238 45106
rect 60722 45054 60734 45106
rect 60786 45054 60798 45106
rect 61170 45054 61182 45106
rect 61234 45054 61246 45106
rect 48974 45042 49026 45054
rect 54014 45042 54066 45054
rect 2046 44994 2098 45006
rect 2046 44930 2098 44942
rect 4846 44994 4898 45006
rect 18622 44994 18674 45006
rect 5730 44942 5742 44994
rect 5794 44942 5806 44994
rect 6514 44942 6526 44994
rect 6578 44942 6590 44994
rect 7298 44942 7310 44994
rect 7362 44942 7374 44994
rect 9986 44942 9998 44994
rect 10050 44942 10062 44994
rect 17714 44942 17726 44994
rect 17778 44942 17790 44994
rect 4846 44930 4898 44942
rect 18622 44930 18674 44942
rect 22654 44994 22706 45006
rect 33966 44994 34018 45006
rect 25666 44942 25678 44994
rect 25730 44942 25742 44994
rect 30034 44942 30046 44994
rect 30098 44942 30110 44994
rect 32162 44942 32174 44994
rect 32226 44942 32238 44994
rect 22654 44930 22706 44942
rect 33966 44930 34018 44942
rect 34638 44994 34690 45006
rect 34638 44930 34690 44942
rect 34862 44994 34914 45006
rect 34862 44930 34914 44942
rect 39678 44994 39730 45006
rect 47406 44994 47458 45006
rect 55246 44994 55298 45006
rect 62190 44994 62242 45006
rect 43138 44942 43150 44994
rect 43202 44942 43214 44994
rect 51426 44942 51438 44994
rect 51490 44942 51502 44994
rect 53218 44942 53230 44994
rect 53282 44942 53294 44994
rect 55906 44942 55918 44994
rect 55970 44942 55982 44994
rect 39678 44930 39730 44942
rect 47406 44930 47458 44942
rect 55246 44930 55298 44942
rect 62190 44930 62242 44942
rect 3838 44882 3890 44894
rect 22766 44882 22818 44894
rect 33294 44882 33346 44894
rect 39902 44882 39954 44894
rect 48862 44882 48914 44894
rect 58830 44882 58882 44894
rect 16706 44830 16718 44882
rect 16770 44830 16782 44882
rect 20290 44830 20302 44882
rect 20354 44830 20366 44882
rect 24434 44830 24446 44882
rect 24498 44830 24510 44882
rect 34290 44830 34302 44882
rect 34354 44830 34366 44882
rect 38322 44830 38334 44882
rect 38386 44830 38398 44882
rect 44258 44830 44270 44882
rect 44322 44830 44334 44882
rect 50642 44830 50654 44882
rect 50706 44830 50718 44882
rect 3838 44818 3890 44830
rect 22766 44818 22818 44830
rect 33294 44818 33346 44830
rect 39902 44818 39954 44830
rect 48862 44818 48914 44830
rect 58830 44818 58882 44830
rect 1344 44714 62608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 62608 44714
rect 1344 44628 62608 44662
rect 2718 44546 2770 44558
rect 32846 44546 32898 44558
rect 41358 44546 41410 44558
rect 29250 44494 29262 44546
rect 29314 44543 29326 44546
rect 29698 44543 29710 44546
rect 29314 44497 29710 44543
rect 29314 44494 29326 44497
rect 29698 44494 29710 44497
rect 29762 44494 29774 44546
rect 36306 44494 36318 44546
rect 36370 44494 36382 44546
rect 2718 44482 2770 44494
rect 32846 44482 32898 44494
rect 41358 44482 41410 44494
rect 42590 44546 42642 44558
rect 42590 44482 42642 44494
rect 42702 44546 42754 44558
rect 42702 44482 42754 44494
rect 43374 44546 43426 44558
rect 43374 44482 43426 44494
rect 43934 44546 43986 44558
rect 59838 44546 59890 44558
rect 51762 44494 51774 44546
rect 51826 44494 51838 44546
rect 54450 44494 54462 44546
rect 54514 44494 54526 44546
rect 43934 44482 43986 44494
rect 59838 44482 59890 44494
rect 60622 44546 60674 44558
rect 60622 44482 60674 44494
rect 60958 44546 61010 44558
rect 60958 44482 61010 44494
rect 3502 44434 3554 44446
rect 3502 44370 3554 44382
rect 4622 44434 4674 44446
rect 12238 44434 12290 44446
rect 26798 44434 26850 44446
rect 5730 44382 5742 44434
rect 5794 44382 5806 44434
rect 8642 44382 8654 44434
rect 8706 44382 8718 44434
rect 10322 44382 10334 44434
rect 10386 44382 10398 44434
rect 16706 44382 16718 44434
rect 16770 44382 16782 44434
rect 23986 44382 23998 44434
rect 24050 44382 24062 44434
rect 24546 44382 24558 44434
rect 24610 44382 24622 44434
rect 4622 44370 4674 44382
rect 12238 44370 12290 44382
rect 26798 44370 26850 44382
rect 28030 44434 28082 44446
rect 28030 44370 28082 44382
rect 29262 44434 29314 44446
rect 29262 44370 29314 44382
rect 29710 44434 29762 44446
rect 29710 44370 29762 44382
rect 30158 44434 30210 44446
rect 39342 44434 39394 44446
rect 41022 44434 41074 44446
rect 34402 44382 34414 44434
rect 34466 44382 34478 44434
rect 37874 44382 37886 44434
rect 37938 44382 37950 44434
rect 40114 44382 40126 44434
rect 40178 44382 40190 44434
rect 46162 44382 46174 44434
rect 46226 44382 46238 44434
rect 53218 44382 53230 44434
rect 53282 44382 53294 44434
rect 30158 44370 30210 44382
rect 39342 44370 39394 44382
rect 41022 44370 41074 44382
rect 3390 44322 3442 44334
rect 4286 44322 4338 44334
rect 8318 44322 8370 44334
rect 12126 44322 12178 44334
rect 18062 44322 18114 44334
rect 21758 44322 21810 44334
rect 1810 44270 1822 44322
rect 1874 44270 1886 44322
rect 3602 44270 3614 44322
rect 3666 44270 3678 44322
rect 4386 44270 4398 44322
rect 4450 44270 4462 44322
rect 4722 44270 4734 44322
rect 4786 44270 4798 44322
rect 6066 44270 6078 44322
rect 6130 44270 6142 44322
rect 6850 44270 6862 44322
rect 6914 44270 6926 44322
rect 7186 44270 7198 44322
rect 7250 44270 7262 44322
rect 7634 44270 7646 44322
rect 7698 44270 7710 44322
rect 10882 44270 10894 44322
rect 10946 44270 10958 44322
rect 13794 44270 13806 44322
rect 13858 44270 13870 44322
rect 18946 44270 18958 44322
rect 19010 44270 19022 44322
rect 20514 44270 20526 44322
rect 20578 44270 20590 44322
rect 3390 44258 3442 44270
rect 4286 44258 4338 44270
rect 8318 44258 8370 44270
rect 12126 44258 12178 44270
rect 18062 44258 18114 44270
rect 21758 44258 21810 44270
rect 21982 44322 22034 44334
rect 21982 44258 22034 44270
rect 22318 44322 22370 44334
rect 34974 44322 35026 44334
rect 37102 44322 37154 44334
rect 38670 44322 38722 44334
rect 23090 44270 23102 44322
rect 23154 44270 23166 44322
rect 23650 44270 23662 44322
rect 23714 44270 23726 44322
rect 24882 44270 24894 44322
rect 24946 44270 24958 44322
rect 25666 44270 25678 44322
rect 25730 44270 25742 44322
rect 34290 44270 34302 44322
rect 34354 44270 34366 44322
rect 36194 44270 36206 44322
rect 36258 44270 36270 44322
rect 37762 44270 37774 44322
rect 37826 44270 37838 44322
rect 22318 44258 22370 44270
rect 34974 44258 35026 44270
rect 37102 44258 37154 44270
rect 38670 44258 38722 44270
rect 43150 44322 43202 44334
rect 44718 44322 44770 44334
rect 43810 44270 43822 44322
rect 43874 44270 43886 44322
rect 43150 44258 43202 44270
rect 44718 44258 44770 44270
rect 44942 44322 44994 44334
rect 44942 44258 44994 44270
rect 45166 44322 45218 44334
rect 50990 44322 51042 44334
rect 46946 44270 46958 44322
rect 47010 44270 47022 44322
rect 47394 44270 47406 44322
rect 47458 44270 47470 44322
rect 48290 44270 48302 44322
rect 48354 44270 48366 44322
rect 48626 44270 48638 44322
rect 48690 44270 48702 44322
rect 49186 44270 49198 44322
rect 49250 44270 49262 44322
rect 50418 44270 50430 44322
rect 50482 44270 50494 44322
rect 52658 44270 52670 44322
rect 52722 44270 52734 44322
rect 54114 44270 54126 44322
rect 54178 44270 54190 44322
rect 55346 44270 55358 44322
rect 55410 44270 55422 44322
rect 56130 44270 56142 44322
rect 56194 44270 56206 44322
rect 45166 44258 45218 44270
rect 50990 44258 51042 44270
rect 2046 44210 2098 44222
rect 2046 44146 2098 44158
rect 2382 44210 2434 44222
rect 2382 44146 2434 44158
rect 2606 44210 2658 44222
rect 2606 44146 2658 44158
rect 3054 44210 3106 44222
rect 3054 44146 3106 44158
rect 4174 44210 4226 44222
rect 11790 44210 11842 44222
rect 5954 44158 5966 44210
rect 6018 44158 6030 44210
rect 4174 44146 4226 44158
rect 11790 44146 11842 44158
rect 12350 44210 12402 44222
rect 17166 44210 17218 44222
rect 27806 44210 27858 44222
rect 37326 44210 37378 44222
rect 14578 44158 14590 44210
rect 14642 44158 14654 44210
rect 18834 44158 18846 44210
rect 18898 44158 18910 44210
rect 20626 44158 20638 44210
rect 20690 44158 20702 44210
rect 23986 44158 23998 44210
rect 24050 44158 24062 44210
rect 25890 44158 25902 44210
rect 25954 44158 25966 44210
rect 26226 44158 26238 44210
rect 26290 44158 26302 44210
rect 27682 44158 27694 44210
rect 27746 44158 27758 44210
rect 31042 44158 31054 44210
rect 31106 44158 31118 44210
rect 12350 44146 12402 44158
rect 17166 44146 17218 44158
rect 27806 44146 27858 44158
rect 37326 44146 37378 44158
rect 37438 44210 37490 44222
rect 37438 44146 37490 44158
rect 39118 44210 39170 44222
rect 42814 44210 42866 44222
rect 40450 44158 40462 44210
rect 40514 44158 40526 44210
rect 41570 44158 41582 44210
rect 41634 44158 41646 44210
rect 42130 44158 42142 44210
rect 42194 44158 42206 44210
rect 39118 44146 39170 44158
rect 42814 44146 42866 44158
rect 45390 44210 45442 44222
rect 50654 44210 50706 44222
rect 53118 44210 53170 44222
rect 49634 44158 49646 44210
rect 49698 44158 49710 44210
rect 51986 44158 51998 44210
rect 52050 44158 52062 44210
rect 56802 44158 56814 44210
rect 56866 44158 56878 44210
rect 61170 44158 61182 44210
rect 61234 44158 61246 44210
rect 61506 44158 61518 44210
rect 61570 44158 61582 44210
rect 45390 44146 45442 44158
rect 50654 44146 50706 44158
rect 53118 44146 53170 44158
rect 3166 44098 3218 44110
rect 3166 44034 3218 44046
rect 12910 44098 12962 44110
rect 12910 44034 12962 44046
rect 17054 44098 17106 44110
rect 17054 44034 17106 44046
rect 17502 44098 17554 44110
rect 17502 44034 17554 44046
rect 22094 44098 22146 44110
rect 27918 44098 27970 44110
rect 22530 44046 22542 44098
rect 22594 44046 22606 44098
rect 22094 44034 22146 44046
rect 27918 44034 27970 44046
rect 28142 44098 28194 44110
rect 28142 44034 28194 44046
rect 28702 44098 28754 44110
rect 28702 44034 28754 44046
rect 38334 44098 38386 44110
rect 53230 44098 53282 44110
rect 48738 44046 48750 44098
rect 48802 44046 48814 44098
rect 38334 44034 38386 44046
rect 53230 44034 53282 44046
rect 53454 44098 53506 44110
rect 58706 44046 58718 44098
rect 58770 44046 58782 44098
rect 53454 44034 53506 44046
rect 1344 43930 62608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 62608 43930
rect 1344 43844 62608 43878
rect 3950 43762 4002 43774
rect 14590 43762 14642 43774
rect 10210 43710 10222 43762
rect 10274 43710 10286 43762
rect 12002 43710 12014 43762
rect 12066 43710 12078 43762
rect 3950 43698 4002 43710
rect 14590 43698 14642 43710
rect 14814 43762 14866 43774
rect 27022 43762 27074 43774
rect 18946 43710 18958 43762
rect 19010 43710 19022 43762
rect 14814 43698 14866 43710
rect 27022 43698 27074 43710
rect 29598 43762 29650 43774
rect 29598 43698 29650 43710
rect 30382 43762 30434 43774
rect 30382 43698 30434 43710
rect 31502 43762 31554 43774
rect 31502 43698 31554 43710
rect 33406 43762 33458 43774
rect 33406 43698 33458 43710
rect 37998 43762 38050 43774
rect 42242 43710 42254 43762
rect 42306 43710 42318 43762
rect 54338 43710 54350 43762
rect 54402 43710 54414 43762
rect 37998 43698 38050 43710
rect 4286 43650 4338 43662
rect 2146 43598 2158 43650
rect 2210 43598 2222 43650
rect 4286 43586 4338 43598
rect 5182 43650 5234 43662
rect 8878 43650 8930 43662
rect 11230 43650 11282 43662
rect 6290 43598 6302 43650
rect 6354 43598 6366 43650
rect 8306 43598 8318 43650
rect 8370 43598 8382 43650
rect 9650 43598 9662 43650
rect 9714 43598 9726 43650
rect 10098 43598 10110 43650
rect 10162 43598 10174 43650
rect 5182 43586 5234 43598
rect 8878 43586 8930 43598
rect 11230 43586 11282 43598
rect 11342 43650 11394 43662
rect 11342 43586 11394 43598
rect 12910 43650 12962 43662
rect 12910 43586 12962 43598
rect 14702 43650 14754 43662
rect 14702 43586 14754 43598
rect 15374 43650 15426 43662
rect 15374 43586 15426 43598
rect 15598 43650 15650 43662
rect 15598 43586 15650 43598
rect 16158 43650 16210 43662
rect 23662 43650 23714 43662
rect 26462 43650 26514 43662
rect 16818 43598 16830 43650
rect 16882 43598 16894 43650
rect 21634 43598 21646 43650
rect 21698 43598 21710 43650
rect 25442 43598 25454 43650
rect 25506 43598 25518 43650
rect 16158 43586 16210 43598
rect 23662 43586 23714 43598
rect 26462 43586 26514 43598
rect 26910 43650 26962 43662
rect 31614 43650 31666 43662
rect 37774 43650 37826 43662
rect 27458 43598 27470 43650
rect 27522 43598 27534 43650
rect 28242 43598 28254 43650
rect 28306 43598 28318 43650
rect 32162 43598 32174 43650
rect 32226 43598 32238 43650
rect 33058 43598 33070 43650
rect 33122 43598 33134 43650
rect 34066 43598 34078 43650
rect 34130 43598 34142 43650
rect 36978 43598 36990 43650
rect 37042 43598 37054 43650
rect 26910 43586 26962 43598
rect 31614 43586 31666 43598
rect 37774 43586 37826 43598
rect 37886 43650 37938 43662
rect 37886 43586 37938 43598
rect 40910 43650 40962 43662
rect 40910 43586 40962 43598
rect 41358 43650 41410 43662
rect 43822 43650 43874 43662
rect 47966 43650 48018 43662
rect 41794 43598 41806 43650
rect 41858 43598 41870 43650
rect 45266 43598 45278 43650
rect 45330 43598 45342 43650
rect 41358 43586 41410 43598
rect 43822 43586 43874 43598
rect 47966 43586 48018 43598
rect 49310 43650 49362 43662
rect 55582 43650 55634 43662
rect 54226 43598 54238 43650
rect 54290 43598 54302 43650
rect 49310 43586 49362 43598
rect 55582 43586 55634 43598
rect 55806 43650 55858 43662
rect 55806 43586 55858 43598
rect 56702 43650 56754 43662
rect 57810 43598 57822 43650
rect 57874 43598 57886 43650
rect 56702 43586 56754 43598
rect 4174 43538 4226 43550
rect 4174 43474 4226 43486
rect 4510 43538 4562 43550
rect 4510 43474 4562 43486
rect 4734 43538 4786 43550
rect 4734 43474 4786 43486
rect 5518 43538 5570 43550
rect 8990 43538 9042 43550
rect 12462 43538 12514 43550
rect 14142 43538 14194 43550
rect 5954 43486 5966 43538
rect 6018 43486 6030 43538
rect 6962 43486 6974 43538
rect 7026 43486 7038 43538
rect 7970 43486 7982 43538
rect 8034 43486 8046 43538
rect 9538 43486 9550 43538
rect 9602 43486 9614 43538
rect 10994 43486 11006 43538
rect 11058 43486 11070 43538
rect 11666 43486 11678 43538
rect 11730 43486 11742 43538
rect 12226 43486 12238 43538
rect 12290 43486 12302 43538
rect 13682 43486 13694 43538
rect 13746 43486 13758 43538
rect 5518 43474 5570 43486
rect 8990 43474 9042 43486
rect 12462 43474 12514 43486
rect 14142 43474 14194 43486
rect 15262 43538 15314 43550
rect 18622 43538 18674 43550
rect 15922 43486 15934 43538
rect 15986 43486 15998 43538
rect 16594 43486 16606 43538
rect 16658 43486 16670 43538
rect 17714 43486 17726 43538
rect 17778 43486 17790 43538
rect 15262 43474 15314 43486
rect 18622 43474 18674 43486
rect 19518 43538 19570 43550
rect 23550 43538 23602 43550
rect 20626 43486 20638 43538
rect 20690 43486 20702 43538
rect 19518 43474 19570 43486
rect 23550 43474 23602 43486
rect 24110 43538 24162 43550
rect 26126 43538 26178 43550
rect 29374 43538 29426 43550
rect 25330 43486 25342 43538
rect 25394 43486 25406 43538
rect 27682 43486 27694 43538
rect 27746 43486 27758 43538
rect 28578 43486 28590 43538
rect 28642 43486 28654 43538
rect 24110 43474 24162 43486
rect 26126 43474 26178 43486
rect 29374 43474 29426 43486
rect 29710 43538 29762 43550
rect 29710 43474 29762 43486
rect 29934 43538 29986 43550
rect 29934 43474 29986 43486
rect 30270 43538 30322 43550
rect 30270 43474 30322 43486
rect 30606 43538 30658 43550
rect 36654 43538 36706 43550
rect 38110 43538 38162 43550
rect 31042 43486 31054 43538
rect 31106 43486 31118 43538
rect 32386 43486 32398 43538
rect 32450 43486 32462 43538
rect 34178 43486 34190 43538
rect 34242 43486 34254 43538
rect 34850 43486 34862 43538
rect 34914 43486 34926 43538
rect 35298 43486 35310 43538
rect 35362 43486 35374 43538
rect 37314 43486 37326 43538
rect 37378 43486 37390 43538
rect 30606 43474 30658 43486
rect 36654 43474 36706 43486
rect 38110 43474 38162 43486
rect 38558 43538 38610 43550
rect 44158 43538 44210 43550
rect 39554 43486 39566 43538
rect 39618 43486 39630 43538
rect 40226 43486 40238 43538
rect 40290 43486 40302 43538
rect 41122 43486 41134 43538
rect 41186 43486 41198 43538
rect 41682 43486 41694 43538
rect 41746 43486 41758 43538
rect 42914 43486 42926 43538
rect 42978 43486 42990 43538
rect 38558 43474 38610 43486
rect 44158 43474 44210 43486
rect 44270 43538 44322 43550
rect 47518 43538 47570 43550
rect 44370 43486 44382 43538
rect 44434 43486 44446 43538
rect 44270 43474 44322 43486
rect 47518 43474 47570 43486
rect 48190 43538 48242 43550
rect 52894 43538 52946 43550
rect 55918 43538 55970 43550
rect 49746 43486 49758 43538
rect 49810 43486 49822 43538
rect 50866 43486 50878 43538
rect 50930 43486 50942 43538
rect 52658 43486 52670 43538
rect 52722 43486 52734 43538
rect 53890 43486 53902 43538
rect 53954 43486 53966 43538
rect 55010 43486 55022 43538
rect 55074 43486 55086 43538
rect 55234 43486 55246 43538
rect 55298 43486 55310 43538
rect 48190 43474 48242 43486
rect 52894 43474 52946 43486
rect 55918 43474 55970 43486
rect 56478 43538 56530 43550
rect 56478 43474 56530 43486
rect 56814 43538 56866 43550
rect 59602 43486 59614 43538
rect 59666 43486 59678 43538
rect 56814 43474 56866 43486
rect 12798 43426 12850 43438
rect 18398 43426 18450 43438
rect 7410 43374 7422 43426
rect 7474 43374 7486 43426
rect 8082 43374 8094 43426
rect 8146 43374 8158 43426
rect 13458 43374 13470 43426
rect 13522 43374 13534 43426
rect 17938 43374 17950 43426
rect 18002 43374 18014 43426
rect 12798 43362 12850 43374
rect 18398 43362 18450 43374
rect 19294 43426 19346 43438
rect 19294 43362 19346 43374
rect 19854 43426 19906 43438
rect 40014 43426 40066 43438
rect 43934 43426 43986 43438
rect 20290 43374 20302 43426
rect 20354 43374 20366 43426
rect 24546 43374 24558 43426
rect 24610 43374 24622 43426
rect 28354 43374 28366 43426
rect 28418 43374 28430 43426
rect 42578 43374 42590 43426
rect 42642 43374 42654 43426
rect 19854 43362 19906 43374
rect 40014 43362 40066 43374
rect 43934 43362 43986 43374
rect 47182 43426 47234 43438
rect 47182 43362 47234 43374
rect 48078 43426 48130 43438
rect 48850 43374 48862 43426
rect 48914 43374 48926 43426
rect 50082 43374 50094 43426
rect 50146 43374 50158 43426
rect 48078 43362 48130 43374
rect 8878 43314 8930 43326
rect 8878 43250 8930 43262
rect 12014 43314 12066 43326
rect 12014 43250 12066 43262
rect 23102 43314 23154 43326
rect 23102 43250 23154 43262
rect 23662 43314 23714 43326
rect 31390 43314 31442 43326
rect 41470 43314 41522 43326
rect 30818 43262 30830 43314
rect 30882 43262 30894 43314
rect 39106 43262 39118 43314
rect 39170 43262 39182 43314
rect 23662 43250 23714 43262
rect 31390 43250 31442 43262
rect 41470 43250 41522 43262
rect 59166 43314 59218 43326
rect 59166 43250 59218 43262
rect 61966 43314 62018 43326
rect 61966 43250 62018 43262
rect 1344 43146 62608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 62608 43146
rect 1344 43060 62608 43094
rect 2494 42978 2546 42990
rect 2494 42914 2546 42926
rect 4174 42978 4226 42990
rect 4174 42914 4226 42926
rect 14702 42978 14754 42990
rect 14702 42914 14754 42926
rect 29262 42978 29314 42990
rect 29262 42914 29314 42926
rect 30046 42978 30098 42990
rect 30046 42914 30098 42926
rect 34750 42978 34802 42990
rect 44270 42978 44322 42990
rect 39890 42926 39902 42978
rect 39954 42926 39966 42978
rect 41010 42926 41022 42978
rect 41074 42926 41086 42978
rect 34750 42914 34802 42926
rect 44270 42914 44322 42926
rect 46062 42978 46114 42990
rect 46062 42914 46114 42926
rect 50878 42978 50930 42990
rect 50878 42914 50930 42926
rect 51214 42978 51266 42990
rect 56366 42978 56418 42990
rect 52770 42926 52782 42978
rect 52834 42926 52846 42978
rect 51214 42914 51266 42926
rect 56366 42914 56418 42926
rect 60622 42978 60674 42990
rect 60622 42914 60674 42926
rect 3278 42866 3330 42878
rect 12462 42866 12514 42878
rect 28142 42866 28194 42878
rect 4610 42814 4622 42866
rect 4674 42814 4686 42866
rect 8642 42814 8654 42866
rect 8706 42814 8718 42866
rect 21522 42814 21534 42866
rect 21586 42814 21598 42866
rect 22642 42814 22654 42866
rect 22706 42814 22718 42866
rect 23874 42814 23886 42866
rect 23938 42814 23950 42866
rect 3278 42802 3330 42814
rect 12462 42802 12514 42814
rect 28142 42802 28194 42814
rect 29822 42866 29874 42878
rect 29822 42802 29874 42814
rect 31726 42866 31778 42878
rect 31726 42802 31778 42814
rect 32510 42866 32562 42878
rect 32510 42802 32562 42814
rect 44158 42866 44210 42878
rect 44158 42802 44210 42814
rect 56478 42866 56530 42878
rect 56478 42802 56530 42814
rect 1822 42754 1874 42766
rect 1822 42690 1874 42702
rect 3726 42754 3778 42766
rect 3726 42690 3778 42702
rect 5630 42754 5682 42766
rect 5630 42690 5682 42702
rect 5966 42754 6018 42766
rect 12798 42754 12850 42766
rect 6626 42702 6638 42754
rect 6690 42702 6702 42754
rect 7074 42702 7086 42754
rect 7138 42702 7150 42754
rect 7634 42702 7646 42754
rect 7698 42702 7710 42754
rect 8306 42702 8318 42754
rect 8370 42702 8382 42754
rect 10546 42702 10558 42754
rect 10610 42702 10622 42754
rect 5966 42690 6018 42702
rect 12798 42690 12850 42702
rect 14254 42754 14306 42766
rect 14254 42690 14306 42702
rect 14590 42754 14642 42766
rect 14590 42690 14642 42702
rect 14814 42754 14866 42766
rect 14814 42690 14866 42702
rect 15150 42754 15202 42766
rect 15150 42690 15202 42702
rect 15374 42754 15426 42766
rect 15374 42690 15426 42702
rect 23102 42754 23154 42766
rect 29486 42754 29538 42766
rect 24098 42702 24110 42754
rect 24162 42702 24174 42754
rect 24882 42702 24894 42754
rect 24946 42702 24958 42754
rect 25218 42702 25230 42754
rect 25282 42702 25294 42754
rect 25666 42702 25678 42754
rect 25730 42702 25742 42754
rect 23102 42690 23154 42702
rect 29486 42690 29538 42702
rect 30494 42754 30546 42766
rect 30942 42754 30994 42766
rect 31502 42754 31554 42766
rect 30706 42702 30718 42754
rect 30770 42702 30782 42754
rect 31154 42702 31166 42754
rect 31218 42702 31230 42754
rect 30494 42690 30546 42702
rect 30942 42690 30994 42702
rect 31502 42690 31554 42702
rect 31838 42754 31890 42766
rect 31838 42690 31890 42702
rect 32062 42754 32114 42766
rect 35086 42754 35138 42766
rect 42814 42754 42866 42766
rect 45726 42754 45778 42766
rect 60958 42754 61010 42766
rect 33170 42702 33182 42754
rect 33234 42702 33246 42754
rect 34290 42702 34302 42754
rect 34354 42702 34366 42754
rect 37650 42702 37662 42754
rect 37714 42702 37726 42754
rect 38882 42702 38894 42754
rect 38946 42702 38958 42754
rect 40226 42702 40238 42754
rect 40290 42702 40302 42754
rect 40786 42702 40798 42754
rect 40850 42702 40862 42754
rect 41346 42702 41358 42754
rect 41410 42702 41422 42754
rect 41682 42702 41694 42754
rect 41746 42702 41758 42754
rect 43586 42702 43598 42754
rect 43650 42702 43662 42754
rect 45266 42702 45278 42754
rect 45330 42702 45342 42754
rect 46722 42702 46734 42754
rect 46786 42702 46798 42754
rect 47842 42702 47854 42754
rect 47906 42702 47918 42754
rect 51762 42702 51774 42754
rect 51826 42702 51838 42754
rect 52882 42702 52894 42754
rect 52946 42702 52958 42754
rect 54562 42702 54574 42754
rect 54626 42702 54638 42754
rect 55906 42702 55918 42754
rect 55970 42702 55982 42754
rect 57250 42702 57262 42754
rect 57314 42702 57326 42754
rect 58146 42702 58158 42754
rect 58210 42702 58222 42754
rect 58930 42702 58942 42754
rect 58994 42702 59006 42754
rect 59714 42702 59726 42754
rect 59778 42702 59790 42754
rect 61394 42702 61406 42754
rect 61458 42702 61470 42754
rect 32062 42690 32114 42702
rect 35086 42690 35138 42702
rect 42814 42690 42866 42702
rect 45726 42690 45778 42702
rect 60958 42690 61010 42702
rect 2830 42642 2882 42654
rect 2146 42590 2158 42642
rect 2210 42590 2222 42642
rect 2830 42578 2882 42590
rect 3166 42642 3218 42654
rect 3166 42578 3218 42590
rect 3502 42642 3554 42654
rect 3502 42578 3554 42590
rect 4062 42642 4114 42654
rect 4062 42578 4114 42590
rect 5742 42642 5794 42654
rect 10334 42642 10386 42654
rect 6290 42590 6302 42642
rect 6354 42590 6366 42642
rect 5742 42578 5794 42590
rect 10334 42578 10386 42590
rect 12350 42642 12402 42654
rect 12350 42578 12402 42590
rect 12686 42642 12738 42654
rect 12686 42578 12738 42590
rect 13694 42642 13746 42654
rect 27246 42642 27298 42654
rect 32622 42642 32674 42654
rect 16258 42590 16270 42642
rect 16322 42590 16334 42642
rect 19058 42590 19070 42642
rect 19122 42590 19134 42642
rect 23426 42590 23438 42642
rect 23490 42590 23502 42642
rect 26226 42590 26238 42642
rect 26290 42590 26302 42642
rect 27346 42590 27358 42642
rect 27410 42590 27422 42642
rect 35298 42590 35310 42642
rect 35362 42590 35374 42642
rect 35634 42590 35646 42642
rect 35698 42590 35710 42642
rect 37762 42590 37774 42642
rect 37826 42590 37838 42642
rect 43474 42590 43486 42642
rect 43538 42590 43550 42642
rect 45042 42590 45054 42642
rect 45106 42590 45118 42642
rect 51986 42590 51998 42642
rect 52050 42590 52062 42642
rect 53218 42590 53230 42642
rect 53282 42590 53294 42642
rect 61618 42590 61630 42642
rect 61682 42590 61694 42642
rect 13694 42578 13746 42590
rect 27246 42578 27298 42590
rect 32622 42578 32674 42590
rect 2606 42530 2658 42542
rect 2606 42466 2658 42478
rect 5070 42530 5122 42542
rect 12126 42530 12178 42542
rect 7186 42478 7198 42530
rect 7250 42478 7262 42530
rect 5070 42466 5122 42478
rect 12126 42466 12178 42478
rect 17950 42530 18002 42542
rect 17950 42466 18002 42478
rect 20302 42530 20354 42542
rect 20302 42466 20354 42478
rect 21982 42530 22034 42542
rect 26910 42530 26962 42542
rect 25218 42478 25230 42530
rect 25282 42478 25294 42530
rect 21982 42466 22034 42478
rect 26910 42466 26962 42478
rect 27022 42530 27074 42542
rect 27022 42466 27074 42478
rect 27134 42530 27186 42542
rect 27134 42466 27186 42478
rect 28030 42530 28082 42542
rect 28030 42466 28082 42478
rect 28254 42530 28306 42542
rect 28254 42466 28306 42478
rect 28478 42530 28530 42542
rect 28478 42466 28530 42478
rect 30158 42530 30210 42542
rect 30158 42466 30210 42478
rect 31278 42530 31330 42542
rect 31278 42466 31330 42478
rect 33406 42530 33458 42542
rect 36542 42530 36594 42542
rect 33730 42478 33742 42530
rect 33794 42478 33806 42530
rect 33406 42466 33458 42478
rect 36542 42466 36594 42478
rect 42478 42530 42530 42542
rect 42478 42466 42530 42478
rect 46510 42530 46562 42542
rect 49410 42478 49422 42530
rect 49474 42478 49486 42530
rect 58594 42478 58606 42530
rect 58658 42478 58670 42530
rect 59490 42478 59502 42530
rect 59554 42478 59566 42530
rect 46510 42466 46562 42478
rect 1344 42362 62608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 62608 42362
rect 1344 42276 62608 42310
rect 3390 42194 3442 42206
rect 12014 42194 12066 42206
rect 14702 42194 14754 42206
rect 5170 42142 5182 42194
rect 5234 42142 5246 42194
rect 12786 42142 12798 42194
rect 12850 42142 12862 42194
rect 3390 42130 3442 42142
rect 12014 42130 12066 42142
rect 14702 42130 14754 42142
rect 15486 42194 15538 42206
rect 15486 42130 15538 42142
rect 16606 42194 16658 42206
rect 16606 42130 16658 42142
rect 18398 42194 18450 42206
rect 18398 42130 18450 42142
rect 26126 42194 26178 42206
rect 26126 42130 26178 42142
rect 35198 42194 35250 42206
rect 42590 42194 42642 42206
rect 41906 42142 41918 42194
rect 41970 42142 41982 42194
rect 35198 42130 35250 42142
rect 42590 42130 42642 42142
rect 44382 42194 44434 42206
rect 53454 42194 53506 42206
rect 45154 42142 45166 42194
rect 45218 42142 45230 42194
rect 46386 42142 46398 42194
rect 46450 42142 46462 42194
rect 48178 42142 48190 42194
rect 48242 42142 48254 42194
rect 54898 42142 54910 42194
rect 54962 42142 54974 42194
rect 57810 42142 57822 42194
rect 57874 42142 57886 42194
rect 44382 42130 44434 42142
rect 53454 42130 53506 42142
rect 3278 42082 3330 42094
rect 3278 42018 3330 42030
rect 3950 42082 4002 42094
rect 3950 42018 4002 42030
rect 6638 42082 6690 42094
rect 6638 42018 6690 42030
rect 6750 42082 6802 42094
rect 6750 42018 6802 42030
rect 6974 42082 7026 42094
rect 7982 42082 8034 42094
rect 7858 42030 7870 42082
rect 7922 42030 7934 42082
rect 6974 42018 7026 42030
rect 7982 42018 8034 42030
rect 8094 42082 8146 42094
rect 14926 42082 14978 42094
rect 10770 42030 10782 42082
rect 10834 42030 10846 42082
rect 12674 42030 12686 42082
rect 12738 42030 12750 42082
rect 13234 42030 13246 42082
rect 13298 42030 13310 42082
rect 8094 42018 8146 42030
rect 14926 42018 14978 42030
rect 15038 42082 15090 42094
rect 15038 42018 15090 42030
rect 18286 42082 18338 42094
rect 26350 42082 26402 42094
rect 19170 42030 19182 42082
rect 19234 42030 19246 42082
rect 20514 42030 20526 42082
rect 20578 42030 20590 42082
rect 21410 42030 21422 42082
rect 21474 42030 21486 42082
rect 18286 42018 18338 42030
rect 26350 42018 26402 42030
rect 26910 42082 26962 42094
rect 26910 42018 26962 42030
rect 27806 42082 27858 42094
rect 27806 42018 27858 42030
rect 27918 42082 27970 42094
rect 42926 42082 42978 42094
rect 31266 42030 31278 42082
rect 31330 42030 31342 42082
rect 33394 42030 33406 42082
rect 33458 42030 33470 42082
rect 36754 42030 36766 42082
rect 36818 42030 36830 42082
rect 41122 42030 41134 42082
rect 41186 42030 41198 42082
rect 49410 42030 49422 42082
rect 49474 42030 49486 42082
rect 51986 42030 51998 42082
rect 52050 42030 52062 42082
rect 54002 42030 54014 42082
rect 54066 42030 54078 42082
rect 58034 42030 58046 42082
rect 58098 42030 58110 42082
rect 27918 42018 27970 42030
rect 42926 42018 42978 42030
rect 2942 41970 2994 41982
rect 2942 41906 2994 41918
rect 3614 41970 3666 41982
rect 3614 41906 3666 41918
rect 3838 41970 3890 41982
rect 3838 41906 3890 41918
rect 6302 41970 6354 41982
rect 6302 41906 6354 41918
rect 7310 41970 7362 41982
rect 7310 41906 7362 41918
rect 8318 41970 8370 41982
rect 12574 41970 12626 41982
rect 8642 41918 8654 41970
rect 8706 41918 8718 41970
rect 8318 41906 8370 41918
rect 12574 41906 12626 41918
rect 13918 41970 13970 41982
rect 13918 41906 13970 41918
rect 14142 41970 14194 41982
rect 14142 41906 14194 41918
rect 14478 41970 14530 41982
rect 14478 41906 14530 41918
rect 15374 41970 15426 41982
rect 17278 41970 17330 41982
rect 15586 41918 15598 41970
rect 15650 41918 15662 41970
rect 16146 41918 16158 41970
rect 16210 41918 16222 41970
rect 16818 41918 16830 41970
rect 16882 41918 16894 41970
rect 15374 41906 15426 41918
rect 17278 41906 17330 41918
rect 17502 41970 17554 41982
rect 17502 41906 17554 41918
rect 17614 41970 17666 41982
rect 17614 41906 17666 41918
rect 17950 41970 18002 41982
rect 20078 41970 20130 41982
rect 22430 41970 22482 41982
rect 19282 41918 19294 41970
rect 19346 41918 19358 41970
rect 20738 41918 20750 41970
rect 20802 41918 20814 41970
rect 21634 41918 21646 41970
rect 21698 41918 21710 41970
rect 17950 41906 18002 41918
rect 20078 41906 20130 41918
rect 22430 41906 22482 41918
rect 22766 41970 22818 41982
rect 22766 41906 22818 41918
rect 23214 41970 23266 41982
rect 23214 41906 23266 41918
rect 23438 41970 23490 41982
rect 23438 41906 23490 41918
rect 24670 41970 24722 41982
rect 24670 41906 24722 41918
rect 25790 41970 25842 41982
rect 25790 41906 25842 41918
rect 26014 41970 26066 41982
rect 29038 41970 29090 41982
rect 26562 41918 26574 41970
rect 26626 41918 26638 41970
rect 27122 41918 27134 41970
rect 27186 41918 27198 41970
rect 28130 41918 28142 41970
rect 28194 41918 28206 41970
rect 26014 41906 26066 41918
rect 29038 41906 29090 41918
rect 30046 41970 30098 41982
rect 30046 41906 30098 41918
rect 30270 41970 30322 41982
rect 30270 41906 30322 41918
rect 30606 41970 30658 41982
rect 37774 41970 37826 41982
rect 42254 41970 42306 41982
rect 31042 41918 31054 41970
rect 31106 41918 31118 41970
rect 39666 41918 39678 41970
rect 39730 41918 39742 41970
rect 40450 41918 40462 41970
rect 40514 41918 40526 41970
rect 40898 41918 40910 41970
rect 40962 41918 40974 41970
rect 42018 41918 42030 41970
rect 42082 41918 42094 41970
rect 30606 41906 30658 41918
rect 37774 41906 37826 41918
rect 42254 41906 42306 41918
rect 42702 41970 42754 41982
rect 42702 41906 42754 41918
rect 43262 41970 43314 41982
rect 44158 41970 44210 41982
rect 45838 41970 45890 41982
rect 43698 41918 43710 41970
rect 43762 41918 43774 41970
rect 45378 41918 45390 41970
rect 45442 41918 45454 41970
rect 43262 41906 43314 41918
rect 44158 41906 44210 41918
rect 45838 41906 45890 41918
rect 46734 41970 46786 41982
rect 46734 41906 46786 41918
rect 47854 41970 47906 41982
rect 55358 41970 55410 41982
rect 53890 41918 53902 41970
rect 53954 41918 53966 41970
rect 54786 41918 54798 41970
rect 54850 41918 54862 41970
rect 47854 41906 47906 41918
rect 55358 41906 55410 41918
rect 55918 41970 55970 41982
rect 62078 41970 62130 41982
rect 57026 41918 57038 41970
rect 57090 41918 57102 41970
rect 58146 41918 58158 41970
rect 58210 41918 58222 41970
rect 58818 41918 58830 41970
rect 58882 41918 58894 41970
rect 55918 41906 55970 41918
rect 62078 41906 62130 41918
rect 2158 41858 2210 41870
rect 2158 41794 2210 41806
rect 2606 41858 2658 41870
rect 9774 41858 9826 41870
rect 7522 41806 7534 41858
rect 7586 41806 7598 41858
rect 2606 41794 2658 41806
rect 9774 41794 9826 41806
rect 14366 41858 14418 41870
rect 30158 41858 30210 41870
rect 24322 41806 24334 41858
rect 24386 41806 24398 41858
rect 25330 41806 25342 41858
rect 25394 41806 25406 41858
rect 29474 41806 29486 41858
rect 29538 41806 29550 41858
rect 14366 41794 14418 41806
rect 30158 41794 30210 41806
rect 31838 41858 31890 41870
rect 31838 41794 31890 41806
rect 35646 41858 35698 41870
rect 35646 41794 35698 41806
rect 38334 41858 38386 41870
rect 46062 41858 46114 41870
rect 39778 41806 39790 41858
rect 39842 41806 39854 41858
rect 44482 41806 44494 41858
rect 44546 41806 44558 41858
rect 38334 41794 38386 41806
rect 46062 41794 46114 41806
rect 47630 41858 47682 41870
rect 47630 41794 47682 41806
rect 50542 41858 50594 41870
rect 50542 41794 50594 41806
rect 51102 41858 51154 41870
rect 51102 41794 51154 41806
rect 57374 41858 57426 41870
rect 59490 41806 59502 41858
rect 59554 41806 59566 41858
rect 61618 41806 61630 41858
rect 61682 41806 61694 41858
rect 57374 41794 57426 41806
rect 3950 41746 4002 41758
rect 3950 41682 4002 41694
rect 8766 41746 8818 41758
rect 8766 41682 8818 41694
rect 9662 41746 9714 41758
rect 16494 41746 16546 41758
rect 15922 41694 15934 41746
rect 15986 41694 15998 41746
rect 9662 41682 9714 41694
rect 16494 41682 16546 41694
rect 18398 41746 18450 41758
rect 18398 41682 18450 41694
rect 19742 41746 19794 41758
rect 19742 41682 19794 41694
rect 22094 41746 22146 41758
rect 22094 41682 22146 41694
rect 32174 41746 32226 41758
rect 46958 41746 47010 41758
rect 39554 41694 39566 41746
rect 39618 41694 39630 41746
rect 47282 41694 47294 41746
rect 47346 41694 47358 41746
rect 32174 41682 32226 41694
rect 46958 41682 47010 41694
rect 1344 41578 62608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 62608 41578
rect 1344 41492 62608 41526
rect 8654 41410 8706 41422
rect 8654 41346 8706 41358
rect 12014 41410 12066 41422
rect 34078 41410 34130 41422
rect 22978 41358 22990 41410
rect 23042 41358 23054 41410
rect 12014 41346 12066 41358
rect 34078 41346 34130 41358
rect 35534 41410 35586 41422
rect 35534 41346 35586 41358
rect 38110 41410 38162 41422
rect 38110 41346 38162 41358
rect 38782 41410 38834 41422
rect 38782 41346 38834 41358
rect 39118 41410 39170 41422
rect 39118 41346 39170 41358
rect 40798 41410 40850 41422
rect 40798 41346 40850 41358
rect 44382 41410 44434 41422
rect 44382 41346 44434 41358
rect 53678 41410 53730 41422
rect 53678 41346 53730 41358
rect 54238 41410 54290 41422
rect 54238 41346 54290 41358
rect 54462 41410 54514 41422
rect 54462 41346 54514 41358
rect 56478 41410 56530 41422
rect 56478 41346 56530 41358
rect 6526 41298 6578 41310
rect 2930 41246 2942 41298
rect 2994 41246 3006 41298
rect 5058 41246 5070 41298
rect 5122 41246 5134 41298
rect 5730 41246 5742 41298
rect 5794 41246 5806 41298
rect 6526 41234 6578 41246
rect 18286 41298 18338 41310
rect 18286 41234 18338 41246
rect 20750 41298 20802 41310
rect 32846 41298 32898 41310
rect 21746 41246 21758 41298
rect 21810 41246 21822 41298
rect 24210 41246 24222 41298
rect 24274 41246 24286 41298
rect 30930 41246 30942 41298
rect 30994 41246 31006 41298
rect 20750 41234 20802 41246
rect 32846 41234 32898 41246
rect 39342 41298 39394 41310
rect 39342 41234 39394 41246
rect 51998 41298 52050 41310
rect 51998 41234 52050 41246
rect 54798 41298 54850 41310
rect 54798 41234 54850 41246
rect 60734 41298 60786 41310
rect 60734 41234 60786 41246
rect 61070 41298 61122 41310
rect 61070 41234 61122 41246
rect 6190 41186 6242 41198
rect 2258 41134 2270 41186
rect 2322 41134 2334 41186
rect 6190 41122 6242 41134
rect 7086 41186 7138 41198
rect 8318 41186 8370 41198
rect 7522 41134 7534 41186
rect 7586 41134 7598 41186
rect 7086 41122 7138 41134
rect 8318 41122 8370 41134
rect 9326 41186 9378 41198
rect 9326 41122 9378 41134
rect 9886 41186 9938 41198
rect 9886 41122 9938 41134
rect 15262 41186 15314 41198
rect 15262 41122 15314 41134
rect 15486 41186 15538 41198
rect 15486 41122 15538 41134
rect 15822 41186 15874 41198
rect 15822 41122 15874 41134
rect 15934 41186 15986 41198
rect 16718 41186 16770 41198
rect 16034 41134 16046 41186
rect 16098 41134 16110 41186
rect 15934 41122 15986 41134
rect 16718 41122 16770 41134
rect 16942 41186 16994 41198
rect 16942 41122 16994 41134
rect 19182 41186 19234 41198
rect 19182 41122 19234 41134
rect 22094 41186 22146 41198
rect 28478 41186 28530 41198
rect 22642 41134 22654 41186
rect 22706 41134 22718 41186
rect 24322 41134 24334 41186
rect 24386 41134 24398 41186
rect 22094 41122 22146 41134
rect 28478 41122 28530 41134
rect 29374 41186 29426 41198
rect 34302 41186 34354 41198
rect 37886 41186 37938 41198
rect 29810 41134 29822 41186
rect 29874 41134 29886 41186
rect 30594 41134 30606 41186
rect 30658 41134 30670 41186
rect 31378 41134 31390 41186
rect 31442 41134 31454 41186
rect 32162 41134 32174 41186
rect 32226 41134 32238 41186
rect 32498 41134 32510 41186
rect 32562 41134 32574 41186
rect 34738 41134 34750 41186
rect 34802 41134 34814 41186
rect 29374 41122 29426 41134
rect 34302 41122 34354 41134
rect 37886 41122 37938 41134
rect 40126 41186 40178 41198
rect 40126 41122 40178 41134
rect 40350 41186 40402 41198
rect 41470 41186 41522 41198
rect 41122 41134 41134 41186
rect 41186 41134 41198 41186
rect 40350 41122 40402 41134
rect 41470 41122 41522 41134
rect 45726 41186 45778 41198
rect 51326 41186 51378 41198
rect 47170 41134 47182 41186
rect 47234 41134 47246 41186
rect 48626 41134 48638 41186
rect 48690 41134 48702 41186
rect 50082 41134 50094 41186
rect 50146 41134 50158 41186
rect 45726 41122 45778 41134
rect 51326 41122 51378 41134
rect 52670 41186 52722 41198
rect 52670 41122 52722 41134
rect 52894 41186 52946 41198
rect 52894 41122 52946 41134
rect 53790 41186 53842 41198
rect 60510 41186 60562 41198
rect 56018 41134 56030 41186
rect 56082 41134 56094 41186
rect 61730 41134 61742 41186
rect 61794 41134 61806 41186
rect 53790 41122 53842 41134
rect 60510 41122 60562 41134
rect 9550 41074 9602 41086
rect 12462 41074 12514 41086
rect 7746 41022 7758 41074
rect 7810 41022 7822 41074
rect 10770 41022 10782 41074
rect 10834 41022 10846 41074
rect 9550 41010 9602 41022
rect 12462 41010 12514 41022
rect 12910 41074 12962 41086
rect 12910 41010 12962 41022
rect 13806 41074 13858 41086
rect 13806 41010 13858 41022
rect 14142 41074 14194 41086
rect 14142 41010 14194 41022
rect 14366 41074 14418 41086
rect 14366 41010 14418 41022
rect 14926 41074 14978 41086
rect 14926 41010 14978 41022
rect 15038 41074 15090 41086
rect 15038 41010 15090 41022
rect 17166 41074 17218 41086
rect 21758 41074 21810 41086
rect 19394 41022 19406 41074
rect 19458 41022 19470 41074
rect 19730 41022 19742 41074
rect 19794 41022 19806 41074
rect 21634 41022 21646 41074
rect 21698 41022 21710 41074
rect 17166 41010 17218 41022
rect 21758 41010 21810 41022
rect 21870 41074 21922 41086
rect 32734 41074 32786 41086
rect 22978 41022 22990 41074
rect 23042 41022 23054 41074
rect 31042 41022 31054 41074
rect 31106 41022 31118 41074
rect 31714 41022 31726 41074
rect 31778 41022 31790 41074
rect 21870 41010 21922 41022
rect 32734 41010 32786 41022
rect 33406 41074 33458 41086
rect 37214 41074 37266 41086
rect 34962 41022 34974 41074
rect 35026 41022 35038 41074
rect 33406 41010 33458 41022
rect 37214 41010 37266 41022
rect 40574 41074 40626 41086
rect 56366 41074 56418 41086
rect 42578 41022 42590 41074
rect 42642 41022 42654 41074
rect 44930 41022 44942 41074
rect 44994 41022 45006 41074
rect 45378 41022 45390 41074
rect 45442 41022 45454 41074
rect 49858 41022 49870 41074
rect 49922 41022 49934 41074
rect 55346 41022 55358 41074
rect 55410 41022 55422 41074
rect 55906 41022 55918 41074
rect 55970 41022 55982 41074
rect 40574 41010 40626 41022
rect 56366 41010 56418 41022
rect 56478 41074 56530 41086
rect 56478 41010 56530 41022
rect 59726 41074 59778 41086
rect 59726 41010 59778 41022
rect 61182 41074 61234 41086
rect 61182 41010 61234 41022
rect 1934 40962 1986 40974
rect 1934 40898 1986 40910
rect 9774 40962 9826 40974
rect 9774 40898 9826 40910
rect 12350 40962 12402 40974
rect 12350 40898 12402 40910
rect 12686 40962 12738 40974
rect 12686 40898 12738 40910
rect 14030 40962 14082 40974
rect 14030 40898 14082 40910
rect 16270 40962 16322 40974
rect 16270 40898 16322 40910
rect 16942 40962 16994 40974
rect 16942 40898 16994 40910
rect 17950 40962 18002 40974
rect 17950 40898 18002 40910
rect 18174 40962 18226 40974
rect 18174 40898 18226 40910
rect 18398 40962 18450 40974
rect 18398 40898 18450 40910
rect 18846 40962 18898 40974
rect 18846 40898 18898 40910
rect 20638 40962 20690 40974
rect 32958 40962 33010 40974
rect 35870 40962 35922 40974
rect 27122 40910 27134 40962
rect 27186 40910 27198 40962
rect 33730 40910 33742 40962
rect 33794 40910 33806 40962
rect 20638 40898 20690 40910
rect 32958 40898 33010 40910
rect 35870 40898 35922 40910
rect 36542 40962 36594 40974
rect 36542 40898 36594 40910
rect 36990 40962 37042 40974
rect 36990 40898 37042 40910
rect 37102 40962 37154 40974
rect 37102 40898 37154 40910
rect 37438 40962 37490 40974
rect 40462 40962 40514 40974
rect 38434 40910 38446 40962
rect 38498 40910 38510 40962
rect 37438 40898 37490 40910
rect 40462 40898 40514 40910
rect 40910 40962 40962 40974
rect 40910 40898 40962 40910
rect 41806 40962 41858 40974
rect 41806 40898 41858 40910
rect 46062 40962 46114 40974
rect 50766 40962 50818 40974
rect 50082 40910 50094 40962
rect 50146 40910 50158 40962
rect 46062 40898 46114 40910
rect 50766 40898 50818 40910
rect 51886 40962 51938 40974
rect 51886 40898 51938 40910
rect 52782 40962 52834 40974
rect 52782 40898 52834 40910
rect 53118 40962 53170 40974
rect 53118 40898 53170 40910
rect 54574 40962 54626 40974
rect 60958 40962 61010 40974
rect 57810 40910 57822 40962
rect 57874 40910 57886 40962
rect 54574 40898 54626 40910
rect 60958 40898 61010 40910
rect 61742 40962 61794 40974
rect 61742 40898 61794 40910
rect 1344 40794 62608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 62608 40794
rect 1344 40708 62608 40742
rect 3726 40626 3778 40638
rect 10334 40626 10386 40638
rect 5170 40574 5182 40626
rect 5234 40574 5246 40626
rect 7746 40574 7758 40626
rect 7810 40574 7822 40626
rect 3726 40562 3778 40574
rect 10334 40562 10386 40574
rect 19518 40626 19570 40638
rect 19518 40562 19570 40574
rect 24446 40626 24498 40638
rect 24446 40562 24498 40574
rect 24670 40626 24722 40638
rect 24670 40562 24722 40574
rect 25342 40626 25394 40638
rect 25342 40562 25394 40574
rect 25902 40626 25954 40638
rect 25902 40562 25954 40574
rect 28702 40626 28754 40638
rect 28702 40562 28754 40574
rect 29486 40626 29538 40638
rect 29486 40562 29538 40574
rect 42814 40626 42866 40638
rect 42814 40562 42866 40574
rect 43038 40626 43090 40638
rect 45390 40626 45442 40638
rect 44258 40574 44270 40626
rect 44322 40574 44334 40626
rect 43038 40562 43090 40574
rect 45390 40562 45442 40574
rect 55470 40626 55522 40638
rect 55470 40562 55522 40574
rect 15598 40514 15650 40526
rect 21982 40514 22034 40526
rect 24334 40514 24386 40526
rect 2706 40462 2718 40514
rect 2770 40462 2782 40514
rect 7074 40462 7086 40514
rect 7138 40462 7150 40514
rect 7522 40462 7534 40514
rect 7586 40462 7598 40514
rect 17714 40462 17726 40514
rect 17778 40462 17790 40514
rect 24098 40462 24110 40514
rect 24162 40462 24174 40514
rect 15598 40450 15650 40462
rect 21982 40450 22034 40462
rect 24334 40450 24386 40462
rect 25678 40514 25730 40526
rect 25678 40450 25730 40462
rect 26014 40514 26066 40526
rect 26014 40450 26066 40462
rect 27694 40514 27746 40526
rect 27694 40450 27746 40462
rect 30270 40514 30322 40526
rect 37214 40514 37266 40526
rect 40238 40514 40290 40526
rect 42702 40514 42754 40526
rect 33618 40462 33630 40514
rect 33682 40462 33694 40514
rect 36082 40462 36094 40514
rect 36146 40462 36158 40514
rect 36530 40462 36542 40514
rect 36594 40462 36606 40514
rect 39218 40462 39230 40514
rect 39282 40462 39294 40514
rect 42466 40462 42478 40514
rect 42530 40462 42542 40514
rect 30270 40450 30322 40462
rect 37214 40450 37266 40462
rect 40238 40450 40290 40462
rect 42702 40450 42754 40462
rect 49310 40514 49362 40526
rect 55694 40514 55746 40526
rect 49970 40462 49982 40514
rect 50034 40462 50046 40514
rect 52434 40462 52446 40514
rect 52498 40462 52510 40514
rect 54226 40462 54238 40514
rect 54290 40462 54302 40514
rect 54562 40462 54574 40514
rect 54626 40462 54638 40514
rect 49310 40450 49362 40462
rect 55694 40450 55746 40462
rect 55806 40514 55858 40526
rect 57586 40462 57598 40514
rect 57650 40462 57662 40514
rect 60610 40462 60622 40514
rect 60674 40462 60686 40514
rect 55806 40450 55858 40462
rect 6302 40402 6354 40414
rect 2594 40350 2606 40402
rect 2658 40350 2670 40402
rect 6302 40338 6354 40350
rect 6750 40402 6802 40414
rect 15710 40402 15762 40414
rect 22094 40402 22146 40414
rect 26238 40402 26290 40414
rect 7410 40350 7422 40402
rect 7474 40350 7486 40402
rect 8530 40350 8542 40402
rect 8594 40350 8606 40402
rect 8978 40350 8990 40402
rect 9042 40350 9054 40402
rect 11330 40350 11342 40402
rect 11394 40350 11406 40402
rect 12114 40350 12126 40402
rect 12178 40350 12190 40402
rect 12786 40350 12798 40402
rect 12850 40350 12862 40402
rect 14578 40350 14590 40402
rect 14642 40350 14654 40402
rect 16818 40350 16830 40402
rect 16882 40350 16894 40402
rect 20178 40350 20190 40402
rect 20242 40350 20254 40402
rect 21410 40350 21422 40402
rect 21474 40350 21486 40402
rect 22530 40350 22542 40402
rect 22594 40350 22606 40402
rect 6750 40338 6802 40350
rect 15710 40338 15762 40350
rect 22094 40338 22146 40350
rect 26238 40338 26290 40350
rect 26798 40402 26850 40414
rect 26798 40338 26850 40350
rect 28926 40402 28978 40414
rect 28926 40338 28978 40350
rect 29150 40402 29202 40414
rect 34862 40402 34914 40414
rect 29474 40350 29486 40402
rect 29538 40350 29550 40402
rect 30034 40350 30046 40402
rect 30098 40350 30110 40402
rect 30482 40350 30494 40402
rect 30546 40350 30558 40402
rect 31266 40350 31278 40402
rect 31330 40350 31342 40402
rect 29150 40338 29202 40350
rect 34862 40338 34914 40350
rect 35646 40402 35698 40414
rect 35646 40338 35698 40350
rect 40126 40402 40178 40414
rect 40126 40338 40178 40350
rect 40462 40402 40514 40414
rect 40462 40338 40514 40350
rect 40798 40402 40850 40414
rect 40798 40338 40850 40350
rect 41134 40402 41186 40414
rect 41134 40338 41186 40350
rect 41358 40402 41410 40414
rect 49646 40402 49698 40414
rect 55134 40402 55186 40414
rect 58606 40402 58658 40414
rect 62078 40402 62130 40414
rect 46834 40350 46846 40402
rect 46898 40350 46910 40402
rect 47282 40350 47294 40402
rect 47346 40350 47358 40402
rect 47618 40350 47630 40402
rect 47682 40350 47694 40402
rect 53218 40350 53230 40402
rect 53282 40350 53294 40402
rect 57810 40350 57822 40402
rect 57874 40350 57886 40402
rect 58930 40350 58942 40402
rect 58994 40350 59006 40402
rect 60498 40350 60510 40402
rect 60562 40350 60574 40402
rect 61394 40350 61406 40402
rect 61458 40350 61470 40402
rect 41358 40338 41410 40350
rect 49646 40338 49698 40350
rect 55134 40338 55186 40350
rect 58606 40338 58658 40350
rect 62078 40338 62130 40350
rect 2270 40290 2322 40302
rect 2270 40226 2322 40238
rect 3390 40290 3442 40302
rect 16270 40290 16322 40302
rect 27358 40290 27410 40302
rect 9874 40238 9886 40290
rect 9938 40238 9950 40290
rect 11442 40238 11454 40290
rect 11506 40238 11518 40290
rect 14690 40238 14702 40290
rect 14754 40238 14766 40290
rect 23874 40238 23886 40290
rect 23938 40238 23950 40290
rect 3390 40226 3442 40238
rect 16270 40226 16322 40238
rect 27358 40226 27410 40238
rect 27918 40290 27970 40302
rect 27918 40226 27970 40238
rect 29038 40290 29090 40302
rect 32622 40290 32674 40302
rect 31154 40238 31166 40290
rect 31218 40238 31230 40290
rect 29038 40226 29090 40238
rect 32622 40226 32674 40238
rect 35422 40290 35474 40302
rect 35422 40226 35474 40238
rect 41022 40290 41074 40302
rect 41022 40226 41074 40238
rect 41918 40290 41970 40302
rect 42690 40238 42702 40290
rect 42754 40238 42766 40290
rect 46050 40238 46062 40290
rect 46114 40238 46126 40290
rect 50306 40238 50318 40290
rect 50370 40238 50382 40290
rect 61170 40238 61182 40290
rect 61234 40238 61246 40290
rect 41918 40226 41970 40238
rect 15598 40178 15650 40190
rect 10994 40126 11006 40178
rect 11058 40126 11070 40178
rect 14578 40126 14590 40178
rect 14642 40126 14654 40178
rect 15598 40114 15650 40126
rect 16494 40178 16546 40190
rect 16494 40114 16546 40126
rect 28254 40178 28306 40190
rect 28254 40114 28306 40126
rect 29822 40178 29874 40190
rect 48750 40178 48802 40190
rect 31602 40126 31614 40178
rect 31666 40126 31678 40178
rect 29822 40114 29874 40126
rect 48750 40114 48802 40126
rect 49086 40178 49138 40190
rect 49086 40114 49138 40126
rect 54798 40178 54850 40190
rect 54798 40114 54850 40126
rect 57262 40178 57314 40190
rect 57262 40114 57314 40126
rect 1344 40010 62608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 62608 40010
rect 1344 39924 62608 39958
rect 16830 39842 16882 39854
rect 8306 39790 8318 39842
rect 8370 39790 8382 39842
rect 12338 39790 12350 39842
rect 12402 39790 12414 39842
rect 16830 39778 16882 39790
rect 21422 39842 21474 39854
rect 44942 39842 44994 39854
rect 52110 39842 52162 39854
rect 28466 39790 28478 39842
rect 28530 39790 28542 39842
rect 30930 39790 30942 39842
rect 30994 39790 31006 39842
rect 49298 39790 49310 39842
rect 49362 39790 49374 39842
rect 21422 39778 21474 39790
rect 44942 39778 44994 39790
rect 52110 39778 52162 39790
rect 62078 39842 62130 39854
rect 62078 39778 62130 39790
rect 4174 39730 4226 39742
rect 4174 39666 4226 39678
rect 6078 39730 6130 39742
rect 13694 39730 13746 39742
rect 7746 39678 7758 39730
rect 7810 39678 7822 39730
rect 12450 39678 12462 39730
rect 12514 39678 12526 39730
rect 6078 39666 6130 39678
rect 13694 39666 13746 39678
rect 14814 39730 14866 39742
rect 26126 39730 26178 39742
rect 32958 39730 33010 39742
rect 41582 39730 41634 39742
rect 44270 39730 44322 39742
rect 24546 39678 24558 39730
rect 24610 39678 24622 39730
rect 28130 39678 28142 39730
rect 28194 39678 28206 39730
rect 31154 39678 31166 39730
rect 31218 39678 31230 39730
rect 40002 39678 40014 39730
rect 40066 39678 40078 39730
rect 43922 39678 43934 39730
rect 43986 39678 43998 39730
rect 14814 39666 14866 39678
rect 26126 39666 26178 39678
rect 32958 39666 33010 39678
rect 41582 39666 41634 39678
rect 44270 39666 44322 39678
rect 53230 39730 53282 39742
rect 53230 39666 53282 39678
rect 53566 39730 53618 39742
rect 59502 39730 59554 39742
rect 53778 39678 53790 39730
rect 53842 39678 53854 39730
rect 57922 39678 57934 39730
rect 57986 39678 57998 39730
rect 61058 39678 61070 39730
rect 61122 39678 61134 39730
rect 53566 39666 53618 39678
rect 59502 39666 59554 39678
rect 4398 39618 4450 39630
rect 4398 39554 4450 39566
rect 6414 39618 6466 39630
rect 9662 39618 9714 39630
rect 6850 39566 6862 39618
rect 6914 39566 6926 39618
rect 7858 39566 7870 39618
rect 7922 39566 7934 39618
rect 8866 39566 8878 39618
rect 8930 39566 8942 39618
rect 6414 39554 6466 39566
rect 9662 39554 9714 39566
rect 9998 39618 10050 39630
rect 11006 39618 11058 39630
rect 10322 39566 10334 39618
rect 10386 39566 10398 39618
rect 9998 39554 10050 39566
rect 11006 39554 11058 39566
rect 11454 39618 11506 39630
rect 23102 39618 23154 39630
rect 27470 39618 27522 39630
rect 14018 39566 14030 39618
rect 14082 39566 14094 39618
rect 15250 39566 15262 39618
rect 15314 39566 15326 39618
rect 18386 39566 18398 39618
rect 18450 39566 18462 39618
rect 19282 39566 19294 39618
rect 19346 39566 19358 39618
rect 20402 39566 20414 39618
rect 20466 39566 20478 39618
rect 21298 39566 21310 39618
rect 21362 39566 21374 39618
rect 23538 39566 23550 39618
rect 23602 39566 23614 39618
rect 24098 39566 24110 39618
rect 24162 39566 24174 39618
rect 26338 39566 26350 39618
rect 26402 39566 26414 39618
rect 11454 39554 11506 39566
rect 23102 39554 23154 39566
rect 27470 39554 27522 39566
rect 28254 39618 28306 39630
rect 28254 39554 28306 39566
rect 29598 39618 29650 39630
rect 29598 39554 29650 39566
rect 31054 39618 31106 39630
rect 32846 39618 32898 39630
rect 31490 39566 31502 39618
rect 31554 39566 31566 39618
rect 31054 39554 31106 39566
rect 32846 39554 32898 39566
rect 33518 39618 33570 39630
rect 47518 39618 47570 39630
rect 33842 39566 33854 39618
rect 33906 39566 33918 39618
rect 35074 39566 35086 39618
rect 35138 39566 35150 39618
rect 37202 39566 37214 39618
rect 37266 39566 37278 39618
rect 40786 39566 40798 39618
rect 40850 39566 40862 39618
rect 41906 39566 41918 39618
rect 41970 39566 41982 39618
rect 42914 39566 42926 39618
rect 42978 39566 42990 39618
rect 33518 39554 33570 39566
rect 47518 39554 47570 39566
rect 47966 39618 48018 39630
rect 49982 39618 50034 39630
rect 51998 39618 52050 39630
rect 58270 39618 58322 39630
rect 59278 39618 59330 39630
rect 49410 39566 49422 39618
rect 49474 39566 49486 39618
rect 50418 39566 50430 39618
rect 50482 39566 50494 39618
rect 56130 39566 56142 39618
rect 56194 39566 56206 39618
rect 59042 39566 59054 39618
rect 59106 39566 59118 39618
rect 47966 39554 48018 39566
rect 49982 39554 50034 39566
rect 51998 39554 52050 39566
rect 58270 39554 58322 39566
rect 59278 39554 59330 39566
rect 59614 39618 59666 39630
rect 59614 39554 59666 39566
rect 59838 39618 59890 39630
rect 60498 39566 60510 39618
rect 60562 39566 60574 39618
rect 61506 39566 61518 39618
rect 61570 39566 61582 39618
rect 59838 39554 59890 39566
rect 6302 39506 6354 39518
rect 2370 39454 2382 39506
rect 2434 39454 2446 39506
rect 6302 39442 6354 39454
rect 7310 39506 7362 39518
rect 7310 39442 7362 39454
rect 8654 39506 8706 39518
rect 17950 39506 18002 39518
rect 27358 39506 27410 39518
rect 47294 39506 47346 39518
rect 54798 39506 54850 39518
rect 12786 39454 12798 39506
rect 12850 39454 12862 39506
rect 14130 39454 14142 39506
rect 14194 39454 14206 39506
rect 14802 39454 14814 39506
rect 14866 39454 14878 39506
rect 16034 39454 16046 39506
rect 16098 39454 16110 39506
rect 16594 39454 16606 39506
rect 16658 39454 16670 39506
rect 17602 39454 17614 39506
rect 17666 39454 17678 39506
rect 22306 39454 22318 39506
rect 22370 39454 22382 39506
rect 22642 39454 22654 39506
rect 22706 39454 22718 39506
rect 29922 39454 29934 39506
rect 29986 39454 29998 39506
rect 30370 39454 30382 39506
rect 30434 39454 30446 39506
rect 33954 39454 33966 39506
rect 34018 39454 34030 39506
rect 35970 39454 35982 39506
rect 36034 39454 36046 39506
rect 37874 39454 37886 39506
rect 37938 39454 37950 39506
rect 41122 39454 41134 39506
rect 41186 39454 41198 39506
rect 41458 39454 41470 39506
rect 41522 39454 41534 39506
rect 42690 39454 42702 39506
rect 42754 39454 42766 39506
rect 46274 39454 46286 39506
rect 46338 39454 46350 39506
rect 48850 39454 48862 39506
rect 48914 39454 48926 39506
rect 54674 39454 54686 39506
rect 54738 39454 54750 39506
rect 8654 39442 8706 39454
rect 17950 39442 18002 39454
rect 27358 39442 27410 39454
rect 47294 39442 47346 39454
rect 54798 39442 54850 39454
rect 56366 39506 56418 39518
rect 62190 39506 62242 39518
rect 60610 39454 60622 39506
rect 60674 39454 60686 39506
rect 56366 39442 56418 39454
rect 62190 39442 62242 39454
rect 3726 39394 3778 39406
rect 9774 39394 9826 39406
rect 17166 39394 17218 39406
rect 4722 39342 4734 39394
rect 4786 39342 4798 39394
rect 10770 39342 10782 39394
rect 10834 39342 10846 39394
rect 3726 39330 3778 39342
rect 9774 39330 9826 39342
rect 17166 39330 17218 39342
rect 18510 39394 18562 39406
rect 29262 39394 29314 39406
rect 22866 39342 22878 39394
rect 22930 39342 22942 39394
rect 18510 39330 18562 39342
rect 29262 39330 29314 39342
rect 32510 39394 32562 39406
rect 32510 39330 32562 39342
rect 33070 39394 33122 39406
rect 33070 39330 33122 39342
rect 40462 39394 40514 39406
rect 40462 39330 40514 39342
rect 43598 39394 43650 39406
rect 43598 39330 43650 39342
rect 47406 39394 47458 39406
rect 47406 39330 47458 39342
rect 52670 39394 52722 39406
rect 52670 39330 52722 39342
rect 54910 39394 54962 39406
rect 54910 39330 54962 39342
rect 55022 39394 55074 39406
rect 55022 39330 55074 39342
rect 55134 39394 55186 39406
rect 55134 39330 55186 39342
rect 1344 39226 62608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 62608 39226
rect 1344 39140 62608 39174
rect 3838 39058 3890 39070
rect 10110 39058 10162 39070
rect 8866 39006 8878 39058
rect 8930 39006 8942 39058
rect 3838 38994 3890 39006
rect 10110 38994 10162 39006
rect 12014 39058 12066 39070
rect 17502 39058 17554 39070
rect 16818 39006 16830 39058
rect 16882 39006 16894 39058
rect 12014 38994 12066 39006
rect 17502 38994 17554 39006
rect 18510 39058 18562 39070
rect 18510 38994 18562 39006
rect 20414 39058 20466 39070
rect 20414 38994 20466 39006
rect 24558 39058 24610 39070
rect 24558 38994 24610 39006
rect 25566 39058 25618 39070
rect 25566 38994 25618 39006
rect 26126 39058 26178 39070
rect 41134 39058 41186 39070
rect 27234 39006 27246 39058
rect 27298 39006 27310 39058
rect 38658 39006 38670 39058
rect 38722 39006 38734 39058
rect 26126 38994 26178 39006
rect 41134 38994 41186 39006
rect 46510 39058 46562 39070
rect 46510 38994 46562 39006
rect 47854 39058 47906 39070
rect 47854 38994 47906 39006
rect 47966 39058 48018 39070
rect 47966 38994 48018 39006
rect 4734 38946 4786 38958
rect 16270 38946 16322 38958
rect 2146 38894 2158 38946
rect 2210 38894 2222 38946
rect 5058 38894 5070 38946
rect 5122 38894 5134 38946
rect 6962 38894 6974 38946
rect 7026 38894 7038 38946
rect 7298 38894 7310 38946
rect 7362 38894 7374 38946
rect 11106 38894 11118 38946
rect 11170 38894 11182 38946
rect 13010 38894 13022 38946
rect 13074 38894 13086 38946
rect 4734 38882 4786 38894
rect 16270 38882 16322 38894
rect 17614 38946 17666 38958
rect 17614 38882 17666 38894
rect 17726 38946 17778 38958
rect 30382 38946 30434 38958
rect 40238 38946 40290 38958
rect 17826 38894 17838 38946
rect 17890 38894 17902 38946
rect 21522 38894 21534 38946
rect 21586 38894 21598 38946
rect 23538 38894 23550 38946
rect 23602 38894 23614 38946
rect 23986 38894 23998 38946
rect 24050 38894 24062 38946
rect 30706 38894 30718 38946
rect 30770 38894 30782 38946
rect 36866 38894 36878 38946
rect 36930 38894 36942 38946
rect 17726 38882 17778 38894
rect 30382 38882 30434 38894
rect 40238 38882 40290 38894
rect 40350 38946 40402 38958
rect 40350 38882 40402 38894
rect 41358 38946 41410 38958
rect 41358 38882 41410 38894
rect 45502 38946 45554 38958
rect 47630 38946 47682 38958
rect 47506 38894 47518 38946
rect 47570 38894 47582 38946
rect 45502 38882 45554 38894
rect 47630 38882 47682 38894
rect 47742 38946 47794 38958
rect 47742 38882 47794 38894
rect 48750 38946 48802 38958
rect 52670 38946 52722 38958
rect 51762 38894 51774 38946
rect 51826 38894 51838 38946
rect 48750 38882 48802 38894
rect 52670 38882 52722 38894
rect 53006 38946 53058 38958
rect 53006 38882 53058 38894
rect 53454 38946 53506 38958
rect 60510 38946 60562 38958
rect 54786 38894 54798 38946
rect 54850 38894 54862 38946
rect 53454 38882 53506 38894
rect 60510 38882 60562 38894
rect 4062 38834 4114 38846
rect 4062 38770 4114 38782
rect 4510 38834 4562 38846
rect 4510 38770 4562 38782
rect 5406 38834 5458 38846
rect 5406 38770 5458 38782
rect 5630 38834 5682 38846
rect 7534 38834 7586 38846
rect 5954 38782 5966 38834
rect 6018 38782 6030 38834
rect 5630 38770 5682 38782
rect 7534 38770 7586 38782
rect 8542 38834 8594 38846
rect 8542 38770 8594 38782
rect 9550 38834 9602 38846
rect 9550 38770 9602 38782
rect 9998 38834 10050 38846
rect 9998 38770 10050 38782
rect 10222 38834 10274 38846
rect 16494 38834 16546 38846
rect 11218 38782 11230 38834
rect 11282 38782 11294 38834
rect 13346 38782 13358 38834
rect 13410 38782 13422 38834
rect 14354 38782 14366 38834
rect 14418 38782 14430 38834
rect 10222 38770 10274 38782
rect 16494 38770 16546 38782
rect 17390 38834 17442 38846
rect 17390 38770 17442 38782
rect 18734 38834 18786 38846
rect 18734 38770 18786 38782
rect 19182 38834 19234 38846
rect 19182 38770 19234 38782
rect 19406 38834 19458 38846
rect 24222 38834 24274 38846
rect 29038 38834 29090 38846
rect 19842 38782 19854 38834
rect 19906 38782 19918 38834
rect 28578 38782 28590 38834
rect 28642 38782 28654 38834
rect 19406 38770 19458 38782
rect 24222 38770 24274 38782
rect 29038 38770 29090 38782
rect 29262 38834 29314 38846
rect 32510 38834 32562 38846
rect 31042 38782 31054 38834
rect 31106 38782 31118 38834
rect 32162 38782 32174 38834
rect 32226 38782 32238 38834
rect 29262 38770 29314 38782
rect 32510 38770 32562 38782
rect 32958 38834 33010 38846
rect 32958 38770 33010 38782
rect 33406 38834 33458 38846
rect 33406 38770 33458 38782
rect 33518 38834 33570 38846
rect 35982 38834 36034 38846
rect 45838 38834 45890 38846
rect 35522 38782 35534 38834
rect 35586 38782 35598 38834
rect 36418 38782 36430 38834
rect 36482 38782 36494 38834
rect 42130 38782 42142 38834
rect 42194 38782 42206 38834
rect 33518 38770 33570 38782
rect 35982 38770 36034 38782
rect 45838 38770 45890 38782
rect 46062 38834 46114 38846
rect 46062 38770 46114 38782
rect 46734 38834 46786 38846
rect 52446 38834 52498 38846
rect 49074 38782 49086 38834
rect 49138 38782 49150 38834
rect 49858 38782 49870 38834
rect 49922 38782 49934 38834
rect 51986 38782 51998 38834
rect 52050 38782 52062 38834
rect 46734 38770 46786 38782
rect 52446 38770 52498 38782
rect 53342 38834 53394 38846
rect 53342 38770 53394 38782
rect 55918 38834 55970 38846
rect 59614 38834 59666 38846
rect 56802 38782 56814 38834
rect 56866 38782 56878 38834
rect 57698 38782 57710 38834
rect 57762 38782 57774 38834
rect 55918 38770 55970 38782
rect 59614 38770 59666 38782
rect 59726 38834 59778 38846
rect 61406 38834 61458 38846
rect 60722 38782 60734 38834
rect 60786 38782 60798 38834
rect 59726 38770 59778 38782
rect 61406 38770 61458 38782
rect 4286 38722 4338 38734
rect 8318 38722 8370 38734
rect 6290 38670 6302 38722
rect 6354 38670 6366 38722
rect 4286 38658 4338 38670
rect 8318 38658 8370 38670
rect 11678 38722 11730 38734
rect 18622 38722 18674 38734
rect 14690 38670 14702 38722
rect 14754 38670 14766 38722
rect 11678 38658 11730 38670
rect 18622 38658 18674 38670
rect 22542 38722 22594 38734
rect 22542 38658 22594 38670
rect 22654 38722 22706 38734
rect 22654 38658 22706 38670
rect 25678 38722 25730 38734
rect 33182 38722 33234 38734
rect 31266 38670 31278 38722
rect 31330 38670 31342 38722
rect 25678 38658 25730 38670
rect 33182 38658 33234 38670
rect 41246 38722 41298 38734
rect 41246 38658 41298 38670
rect 41582 38722 41634 38734
rect 46622 38722 46674 38734
rect 50878 38722 50930 38734
rect 42914 38670 42926 38722
rect 42978 38670 42990 38722
rect 45042 38670 45054 38722
rect 45106 38670 45118 38722
rect 49186 38670 49198 38722
rect 49250 38670 49262 38722
rect 50306 38670 50318 38722
rect 50370 38670 50382 38722
rect 41582 38658 41634 38670
rect 46622 38658 46674 38670
rect 50878 38658 50930 38670
rect 52894 38722 52946 38734
rect 57250 38670 57262 38722
rect 57314 38670 57326 38722
rect 61842 38670 61854 38722
rect 61906 38670 61918 38722
rect 52894 38658 52946 38670
rect 7870 38610 7922 38622
rect 7870 38546 7922 38558
rect 12686 38610 12738 38622
rect 12686 38546 12738 38558
rect 28702 38610 28754 38622
rect 28702 38546 28754 38558
rect 37438 38610 37490 38622
rect 37438 38546 37490 38558
rect 39790 38610 39842 38622
rect 39790 38546 39842 38558
rect 41806 38610 41858 38622
rect 41806 38546 41858 38558
rect 51214 38610 51266 38622
rect 51214 38546 51266 38558
rect 53454 38610 53506 38622
rect 53454 38546 53506 38558
rect 1344 38442 62608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 62608 38442
rect 1344 38356 62608 38390
rect 17278 38274 17330 38286
rect 58494 38274 58546 38286
rect 13570 38222 13582 38274
rect 13634 38222 13646 38274
rect 25218 38222 25230 38274
rect 25282 38222 25294 38274
rect 34178 38222 34190 38274
rect 34242 38222 34254 38274
rect 42690 38222 42702 38274
rect 42754 38222 42766 38274
rect 55794 38222 55806 38274
rect 55858 38222 55870 38274
rect 17278 38210 17330 38222
rect 58494 38210 58546 38222
rect 2046 38162 2098 38174
rect 2046 38098 2098 38110
rect 2382 38162 2434 38174
rect 20302 38162 20354 38174
rect 46398 38162 46450 38174
rect 3602 38110 3614 38162
rect 3666 38110 3678 38162
rect 4946 38110 4958 38162
rect 5010 38110 5022 38162
rect 11666 38110 11678 38162
rect 11730 38110 11742 38162
rect 12674 38110 12686 38162
rect 12738 38110 12750 38162
rect 22978 38110 22990 38162
rect 23042 38110 23054 38162
rect 28130 38110 28142 38162
rect 28194 38110 28206 38162
rect 32050 38110 32062 38162
rect 32114 38110 32126 38162
rect 34402 38110 34414 38162
rect 34466 38110 34478 38162
rect 43922 38110 43934 38162
rect 43986 38110 43998 38162
rect 44930 38110 44942 38162
rect 44994 38110 45006 38162
rect 2382 38098 2434 38110
rect 20302 38098 20354 38110
rect 46398 38098 46450 38110
rect 8094 38050 8146 38062
rect 3714 37998 3726 38050
rect 3778 37998 3790 38050
rect 4722 37998 4734 38050
rect 4786 37998 4798 38050
rect 8094 37986 8146 37998
rect 8318 38050 8370 38062
rect 8990 38050 9042 38062
rect 15150 38050 15202 38062
rect 19854 38050 19906 38062
rect 8642 37998 8654 38050
rect 8706 37998 8718 38050
rect 9538 37998 9550 38050
rect 9602 37998 9614 38050
rect 10434 37998 10446 38050
rect 10498 37998 10510 38050
rect 10994 37998 11006 38050
rect 11058 37998 11070 38050
rect 13682 37998 13694 38050
rect 13746 37998 13758 38050
rect 15586 37998 15598 38050
rect 15650 37998 15662 38050
rect 8318 37986 8370 37998
rect 8990 37986 9042 37998
rect 15150 37986 15202 37998
rect 19854 37986 19906 37998
rect 20414 38050 20466 38062
rect 20414 37986 20466 37998
rect 21198 38050 21250 38062
rect 21198 37986 21250 37998
rect 21534 38050 21586 38062
rect 25566 38050 25618 38062
rect 34862 38050 34914 38062
rect 37998 38050 38050 38062
rect 46062 38050 46114 38062
rect 22418 37998 22430 38050
rect 22482 37998 22494 38050
rect 23314 37998 23326 38050
rect 23378 37998 23390 38050
rect 24098 37998 24110 38050
rect 24162 37998 24174 38050
rect 25778 37998 25790 38050
rect 25842 37998 25854 38050
rect 28466 37998 28478 38050
rect 28530 37998 28542 38050
rect 29810 37998 29822 38050
rect 29874 37998 29886 38050
rect 30146 37998 30158 38050
rect 30210 37998 30222 38050
rect 31938 37998 31950 38050
rect 32002 37998 32014 38050
rect 34066 37998 34078 38050
rect 34130 37998 34142 38050
rect 35074 37998 35086 38050
rect 35138 37998 35150 38050
rect 36082 37998 36094 38050
rect 36146 37998 36158 38050
rect 41682 37998 41694 38050
rect 41746 37998 41758 38050
rect 42690 37998 42702 38050
rect 42754 37998 42766 38050
rect 43810 37998 43822 38050
rect 43874 37998 43886 38050
rect 45266 37998 45278 38050
rect 45330 37998 45342 38050
rect 21534 37986 21586 37998
rect 25566 37986 25618 37998
rect 34862 37986 34914 37998
rect 37998 37986 38050 37998
rect 46062 37986 46114 37998
rect 46622 38050 46674 38062
rect 46622 37986 46674 37998
rect 47182 38050 47234 38062
rect 47182 37986 47234 37998
rect 48414 38050 48466 38062
rect 58830 38050 58882 38062
rect 60510 38050 60562 38062
rect 48962 37998 48974 38050
rect 49026 37998 49038 38050
rect 50754 37998 50766 38050
rect 50818 37998 50830 38050
rect 52098 37998 52110 38050
rect 52162 37998 52174 38050
rect 52658 37998 52670 38050
rect 52722 37998 52734 38050
rect 53218 37998 53230 38050
rect 53282 37998 53294 38050
rect 53778 37998 53790 38050
rect 53842 37998 53854 38050
rect 54786 37998 54798 38050
rect 54850 37998 54862 38050
rect 55906 37998 55918 38050
rect 55970 37998 55982 38050
rect 57810 37998 57822 38050
rect 57874 37998 57886 38050
rect 59490 37998 59502 38050
rect 59554 37998 59566 38050
rect 61282 37998 61294 38050
rect 61346 37998 61358 38050
rect 61954 37998 61966 38050
rect 62018 37998 62030 38050
rect 48414 37986 48466 37998
rect 58830 37986 58882 37998
rect 60510 37986 60562 37998
rect 2606 37938 2658 37950
rect 3390 37938 3442 37950
rect 9102 37938 9154 37950
rect 19518 37938 19570 37950
rect 2706 37886 2718 37938
rect 2770 37886 2782 37938
rect 6066 37886 6078 37938
rect 6130 37886 6142 37938
rect 14354 37886 14366 37938
rect 14418 37886 14430 37938
rect 18498 37886 18510 37938
rect 18562 37886 18574 37938
rect 2606 37874 2658 37886
rect 3390 37874 3442 37886
rect 9102 37874 9154 37886
rect 19518 37874 19570 37886
rect 21422 37938 21474 37950
rect 21422 37874 21474 37886
rect 21870 37938 21922 37950
rect 21870 37874 21922 37886
rect 22878 37938 22930 37950
rect 29150 37938 29202 37950
rect 24546 37886 24558 37938
rect 24610 37886 24622 37938
rect 22878 37874 22930 37886
rect 29150 37874 29202 37886
rect 29486 37938 29538 37950
rect 37214 37938 37266 37950
rect 43262 37938 43314 37950
rect 32946 37886 32958 37938
rect 33010 37886 33022 37938
rect 38210 37886 38222 37938
rect 38274 37886 38286 37938
rect 38658 37886 38670 37938
rect 38722 37886 38734 37938
rect 40002 37886 40014 37938
rect 40066 37886 40078 37938
rect 43026 37886 43038 37938
rect 43090 37886 43102 37938
rect 29486 37874 29538 37886
rect 37214 37874 37266 37886
rect 43262 37874 43314 37886
rect 44158 37938 44210 37950
rect 44158 37874 44210 37886
rect 45726 37938 45778 37950
rect 45726 37874 45778 37886
rect 45838 37938 45890 37950
rect 45838 37874 45890 37886
rect 46286 37938 46338 37950
rect 46286 37874 46338 37886
rect 46846 37938 46898 37950
rect 46846 37874 46898 37886
rect 47294 37938 47346 37950
rect 48078 37938 48130 37950
rect 47842 37886 47854 37938
rect 47906 37886 47918 37938
rect 47294 37874 47346 37886
rect 48078 37874 48130 37886
rect 48190 37938 48242 37950
rect 50318 37938 50370 37950
rect 60846 37938 60898 37950
rect 49298 37886 49310 37938
rect 49362 37886 49374 37938
rect 53442 37886 53454 37938
rect 53506 37886 53518 37938
rect 53890 37886 53902 37938
rect 53954 37886 53966 37938
rect 57138 37886 57150 37938
rect 57202 37886 57214 37938
rect 59602 37886 59614 37938
rect 59666 37886 59678 37938
rect 48190 37874 48242 37886
rect 50318 37874 50370 37886
rect 60846 37874 60898 37886
rect 2270 37826 2322 37838
rect 2270 37762 2322 37774
rect 2494 37826 2546 37838
rect 2494 37762 2546 37774
rect 7758 37826 7810 37838
rect 7758 37762 7810 37774
rect 9326 37826 9378 37838
rect 9326 37762 9378 37774
rect 12238 37826 12290 37838
rect 12238 37762 12290 37774
rect 20190 37826 20242 37838
rect 20190 37762 20242 37774
rect 20638 37826 20690 37838
rect 20638 37762 20690 37774
rect 27806 37826 27858 37838
rect 36878 37826 36930 37838
rect 35858 37774 35870 37826
rect 35922 37774 35934 37826
rect 27806 37762 27858 37774
rect 36878 37762 36930 37774
rect 37102 37826 37154 37838
rect 37102 37762 37154 37774
rect 37662 37826 37714 37838
rect 37662 37762 37714 37774
rect 43150 37826 43202 37838
rect 43150 37762 43202 37774
rect 48302 37826 48354 37838
rect 48302 37762 48354 37774
rect 60622 37826 60674 37838
rect 60622 37762 60674 37774
rect 60734 37826 60786 37838
rect 61618 37774 61630 37826
rect 61682 37774 61694 37826
rect 60734 37762 60786 37774
rect 1344 37658 62608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 62608 37658
rect 1344 37572 62608 37606
rect 2046 37490 2098 37502
rect 2046 37426 2098 37438
rect 3054 37490 3106 37502
rect 8318 37490 8370 37502
rect 6402 37438 6414 37490
rect 6466 37438 6478 37490
rect 3054 37426 3106 37438
rect 8318 37426 8370 37438
rect 8654 37490 8706 37502
rect 8654 37426 8706 37438
rect 15710 37490 15762 37502
rect 15710 37426 15762 37438
rect 15822 37490 15874 37502
rect 15822 37426 15874 37438
rect 15934 37490 15986 37502
rect 15934 37426 15986 37438
rect 25342 37490 25394 37502
rect 25342 37426 25394 37438
rect 32510 37490 32562 37502
rect 32510 37426 32562 37438
rect 40910 37490 40962 37502
rect 40910 37426 40962 37438
rect 41134 37490 41186 37502
rect 47966 37490 48018 37502
rect 52670 37490 52722 37502
rect 43474 37438 43486 37490
rect 43538 37438 43550 37490
rect 48850 37438 48862 37490
rect 48914 37438 48926 37490
rect 51202 37438 51214 37490
rect 51266 37438 51278 37490
rect 41134 37426 41186 37438
rect 47966 37426 48018 37438
rect 52670 37426 52722 37438
rect 54014 37490 54066 37502
rect 61842 37438 61854 37490
rect 61906 37438 61918 37490
rect 54014 37426 54066 37438
rect 2718 37378 2770 37390
rect 2482 37326 2494 37378
rect 2546 37326 2558 37378
rect 2718 37314 2770 37326
rect 2830 37378 2882 37390
rect 8878 37378 8930 37390
rect 7410 37326 7422 37378
rect 7474 37326 7486 37378
rect 2830 37314 2882 37326
rect 8878 37314 8930 37326
rect 8990 37378 9042 37390
rect 14478 37378 14530 37390
rect 10210 37326 10222 37378
rect 10274 37326 10286 37378
rect 8990 37314 9042 37326
rect 14478 37314 14530 37326
rect 16046 37378 16098 37390
rect 25678 37378 25730 37390
rect 16146 37326 16158 37378
rect 16210 37326 16222 37378
rect 18610 37326 18622 37378
rect 18674 37326 18686 37378
rect 21634 37326 21646 37378
rect 21698 37326 21710 37378
rect 16046 37314 16098 37326
rect 25678 37314 25730 37326
rect 26574 37378 26626 37390
rect 41358 37378 41410 37390
rect 37426 37326 37438 37378
rect 37490 37326 37502 37378
rect 39666 37326 39678 37378
rect 39730 37326 39742 37378
rect 26574 37314 26626 37326
rect 41358 37314 41410 37326
rect 41918 37378 41970 37390
rect 41918 37314 41970 37326
rect 42142 37378 42194 37390
rect 46734 37378 46786 37390
rect 56590 37378 56642 37390
rect 43362 37326 43374 37378
rect 43426 37326 43438 37378
rect 45826 37326 45838 37378
rect 45890 37326 45902 37378
rect 46386 37326 46398 37378
rect 46450 37326 46462 37378
rect 49410 37326 49422 37378
rect 49474 37326 49486 37378
rect 50306 37326 50318 37378
rect 50370 37326 50382 37378
rect 55794 37326 55806 37378
rect 55858 37326 55870 37378
rect 42142 37314 42194 37326
rect 46734 37314 46786 37326
rect 56590 37314 56642 37326
rect 56702 37378 56754 37390
rect 60050 37326 60062 37378
rect 60114 37326 60126 37378
rect 56702 37314 56754 37326
rect 12574 37266 12626 37278
rect 17502 37266 17554 37278
rect 25902 37266 25954 37278
rect 3602 37214 3614 37266
rect 3666 37214 3678 37266
rect 5282 37214 5294 37266
rect 5346 37214 5358 37266
rect 6626 37214 6638 37266
rect 6690 37214 6702 37266
rect 7186 37214 7198 37266
rect 7250 37214 7262 37266
rect 12002 37214 12014 37266
rect 12066 37214 12078 37266
rect 14242 37214 14254 37266
rect 14306 37214 14318 37266
rect 14690 37214 14702 37266
rect 14754 37214 14766 37266
rect 17938 37214 17950 37266
rect 18002 37214 18014 37266
rect 12574 37202 12626 37214
rect 17502 37202 17554 37214
rect 25902 37202 25954 37214
rect 27022 37266 27074 37278
rect 29374 37266 29426 37278
rect 27682 37214 27694 37266
rect 27746 37214 27758 37266
rect 28578 37214 28590 37266
rect 28642 37214 28654 37266
rect 27022 37202 27074 37214
rect 29374 37202 29426 37214
rect 31166 37266 31218 37278
rect 31166 37202 31218 37214
rect 31502 37266 31554 37278
rect 41022 37266 41074 37278
rect 33394 37214 33406 37266
rect 33458 37214 33470 37266
rect 33618 37214 33630 37266
rect 33682 37214 33694 37266
rect 36418 37214 36430 37266
rect 36482 37214 36494 37266
rect 37986 37214 37998 37266
rect 38050 37214 38062 37266
rect 39330 37214 39342 37266
rect 39394 37214 39406 37266
rect 40338 37214 40350 37266
rect 40402 37214 40414 37266
rect 31502 37202 31554 37214
rect 41022 37202 41074 37214
rect 43150 37266 43202 37278
rect 43150 37202 43202 37214
rect 43598 37266 43650 37278
rect 46622 37266 46674 37278
rect 48190 37266 48242 37278
rect 51550 37266 51602 37278
rect 43698 37214 43710 37266
rect 43762 37214 43774 37266
rect 44258 37214 44270 37266
rect 44322 37214 44334 37266
rect 47506 37214 47518 37266
rect 47570 37214 47582 37266
rect 47730 37214 47742 37266
rect 47794 37214 47806 37266
rect 48738 37214 48750 37266
rect 48802 37214 48814 37266
rect 49298 37214 49310 37266
rect 49362 37214 49374 37266
rect 50194 37214 50206 37266
rect 50258 37214 50270 37266
rect 51090 37214 51102 37266
rect 51154 37214 51166 37266
rect 43598 37202 43650 37214
rect 46622 37202 46674 37214
rect 48190 37202 48242 37214
rect 51550 37202 51602 37214
rect 51886 37266 51938 37278
rect 51886 37202 51938 37214
rect 52222 37266 52274 37278
rect 53566 37266 53618 37278
rect 52546 37214 52558 37266
rect 52610 37214 52622 37266
rect 52222 37202 52274 37214
rect 53566 37202 53618 37214
rect 54238 37266 54290 37278
rect 56926 37266 56978 37278
rect 54898 37214 54910 37266
rect 54962 37214 54974 37266
rect 56018 37214 56030 37266
rect 56082 37214 56094 37266
rect 58482 37214 58494 37266
rect 58546 37214 58558 37266
rect 60386 37214 60398 37266
rect 60450 37214 60462 37266
rect 61058 37214 61070 37266
rect 61122 37214 61134 37266
rect 62066 37214 62078 37266
rect 62130 37214 62142 37266
rect 54238 37202 54290 37214
rect 56926 37202 56978 37214
rect 24670 37154 24722 37166
rect 2706 37102 2718 37154
rect 2770 37102 2782 37154
rect 3490 37102 3502 37154
rect 3554 37102 3566 37154
rect 5730 37102 5742 37154
rect 5794 37102 5806 37154
rect 20738 37102 20750 37154
rect 20802 37102 20814 37154
rect 24670 37090 24722 37102
rect 26238 37154 26290 37166
rect 38782 37154 38834 37166
rect 47182 37154 47234 37166
rect 27906 37102 27918 37154
rect 27970 37102 27982 37154
rect 28914 37102 28926 37154
rect 28978 37102 28990 37154
rect 33842 37102 33854 37154
rect 33906 37102 33918 37154
rect 36194 37102 36206 37154
rect 36258 37102 36270 37154
rect 39778 37102 39790 37154
rect 39842 37102 39854 37154
rect 44370 37102 44382 37154
rect 44434 37102 44446 37154
rect 26238 37090 26290 37102
rect 38782 37090 38834 37102
rect 47182 37090 47234 37102
rect 48078 37154 48130 37166
rect 48078 37090 48130 37102
rect 51774 37154 51826 37166
rect 51774 37090 51826 37102
rect 54126 37154 54178 37166
rect 61518 37154 61570 37166
rect 55346 37102 55358 37154
rect 55410 37102 55422 37154
rect 58370 37102 58382 37154
rect 58434 37102 58446 37154
rect 54126 37090 54178 37102
rect 61518 37090 61570 37102
rect 7982 37042 8034 37054
rect 7982 36978 8034 36990
rect 11342 37042 11394 37054
rect 11342 36978 11394 36990
rect 23662 37042 23714 37054
rect 23662 36978 23714 36990
rect 26686 37042 26738 37054
rect 26686 36978 26738 36990
rect 26910 37042 26962 37054
rect 42030 37042 42082 37054
rect 33170 36990 33182 37042
rect 33234 36990 33246 37042
rect 35970 36990 35982 37042
rect 36034 36990 36046 37042
rect 26910 36978 26962 36990
rect 42030 36978 42082 36990
rect 42478 37042 42530 37054
rect 42478 36978 42530 36990
rect 42702 37042 42754 37054
rect 57698 36990 57710 37042
rect 57762 36990 57774 37042
rect 42702 36978 42754 36990
rect 1344 36874 62608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 62608 36874
rect 1344 36788 62608 36822
rect 6526 36706 6578 36718
rect 48750 36706 48802 36718
rect 4162 36654 4174 36706
rect 4226 36654 4238 36706
rect 12786 36654 12798 36706
rect 12850 36654 12862 36706
rect 24658 36654 24670 36706
rect 24722 36654 24734 36706
rect 6526 36642 6578 36654
rect 48750 36642 48802 36654
rect 57374 36706 57426 36718
rect 57374 36642 57426 36654
rect 2494 36594 2546 36606
rect 5070 36594 5122 36606
rect 27918 36594 27970 36606
rect 37886 36594 37938 36606
rect 46846 36594 46898 36606
rect 3938 36542 3950 36594
rect 4002 36542 4014 36594
rect 8978 36542 8990 36594
rect 9042 36542 9054 36594
rect 13906 36542 13918 36594
rect 13970 36542 13982 36594
rect 17490 36542 17502 36594
rect 17554 36542 17566 36594
rect 18274 36542 18286 36594
rect 18338 36542 18350 36594
rect 20514 36542 20526 36594
rect 20578 36542 20590 36594
rect 23314 36542 23326 36594
rect 23378 36542 23390 36594
rect 32162 36542 32174 36594
rect 32226 36542 32238 36594
rect 46162 36542 46174 36594
rect 46226 36542 46238 36594
rect 2494 36530 2546 36542
rect 5070 36530 5122 36542
rect 27918 36530 27970 36542
rect 37886 36530 37938 36542
rect 46846 36530 46898 36542
rect 56030 36594 56082 36606
rect 56030 36530 56082 36542
rect 60622 36594 60674 36606
rect 60622 36530 60674 36542
rect 11230 36482 11282 36494
rect 19294 36482 19346 36494
rect 22318 36482 22370 36494
rect 25454 36482 25506 36494
rect 28254 36482 28306 36494
rect 35086 36482 35138 36494
rect 3266 36430 3278 36482
rect 3330 36430 3342 36482
rect 4386 36430 4398 36482
rect 4450 36430 4462 36482
rect 10994 36430 11006 36482
rect 11058 36430 11070 36482
rect 11778 36430 11790 36482
rect 11842 36430 11854 36482
rect 16818 36430 16830 36482
rect 16882 36430 16894 36482
rect 17602 36430 17614 36482
rect 17666 36430 17678 36482
rect 18386 36430 18398 36482
rect 18450 36430 18462 36482
rect 19730 36430 19742 36482
rect 19794 36430 19806 36482
rect 20738 36430 20750 36482
rect 20802 36430 20814 36482
rect 21634 36430 21646 36482
rect 21698 36430 21710 36482
rect 23986 36430 23998 36482
rect 24050 36430 24062 36482
rect 25666 36430 25678 36482
rect 25730 36430 25742 36482
rect 28018 36430 28030 36482
rect 28082 36430 28094 36482
rect 28354 36430 28366 36482
rect 28418 36430 28430 36482
rect 29362 36430 29374 36482
rect 29426 36430 29438 36482
rect 30370 36430 30382 36482
rect 30434 36430 30446 36482
rect 31602 36430 31614 36482
rect 31666 36430 31678 36482
rect 31938 36430 31950 36482
rect 32002 36430 32014 36482
rect 11230 36418 11282 36430
rect 19294 36418 19346 36430
rect 22318 36418 22370 36430
rect 25454 36418 25506 36430
rect 28254 36418 28306 36430
rect 35086 36418 35138 36430
rect 35870 36482 35922 36494
rect 35870 36418 35922 36430
rect 37438 36482 37490 36494
rect 37438 36418 37490 36430
rect 37774 36482 37826 36494
rect 41470 36482 41522 36494
rect 39890 36430 39902 36482
rect 39954 36430 39966 36482
rect 37774 36418 37826 36430
rect 41470 36418 41522 36430
rect 42030 36482 42082 36494
rect 42030 36418 42082 36430
rect 44830 36482 44882 36494
rect 44830 36418 44882 36430
rect 45054 36482 45106 36494
rect 47854 36482 47906 36494
rect 46386 36430 46398 36482
rect 46450 36430 46462 36482
rect 47170 36430 47182 36482
rect 47234 36430 47246 36482
rect 45054 36418 45106 36430
rect 47854 36418 47906 36430
rect 48190 36482 48242 36494
rect 50206 36482 50258 36494
rect 52782 36482 52834 36494
rect 48738 36430 48750 36482
rect 48802 36430 48814 36482
rect 50418 36430 50430 36482
rect 50482 36430 50494 36482
rect 48190 36418 48242 36430
rect 50206 36418 50258 36430
rect 52782 36418 52834 36430
rect 52894 36482 52946 36494
rect 52894 36418 52946 36430
rect 53118 36482 53170 36494
rect 53118 36418 53170 36430
rect 54014 36482 54066 36494
rect 61294 36482 61346 36494
rect 54450 36430 54462 36482
rect 54514 36430 54526 36482
rect 55794 36430 55806 36482
rect 55858 36430 55870 36482
rect 56690 36430 56702 36482
rect 56754 36430 56766 36482
rect 54014 36418 54066 36430
rect 61294 36418 61346 36430
rect 61630 36482 61682 36494
rect 61630 36418 61682 36430
rect 61966 36482 62018 36494
rect 61966 36418 62018 36430
rect 2158 36370 2210 36382
rect 2158 36306 2210 36318
rect 2942 36370 2994 36382
rect 9214 36370 9266 36382
rect 17950 36370 18002 36382
rect 5618 36318 5630 36370
rect 5682 36318 5694 36370
rect 12002 36318 12014 36370
rect 12066 36318 12078 36370
rect 16034 36318 16046 36370
rect 16098 36318 16110 36370
rect 2942 36306 2994 36318
rect 9214 36306 9266 36318
rect 17950 36306 18002 36318
rect 22542 36370 22594 36382
rect 27806 36370 27858 36382
rect 24322 36318 24334 36370
rect 24386 36318 24398 36370
rect 22542 36306 22594 36318
rect 27806 36306 27858 36318
rect 29150 36370 29202 36382
rect 36430 36370 36482 36382
rect 32946 36318 32958 36370
rect 33010 36318 33022 36370
rect 34514 36318 34526 36370
rect 34578 36318 34590 36370
rect 34850 36318 34862 36370
rect 34914 36318 34926 36370
rect 29150 36306 29202 36318
rect 36430 36306 36482 36318
rect 39678 36370 39730 36382
rect 39678 36306 39730 36318
rect 40910 36370 40962 36382
rect 48078 36370 48130 36382
rect 53230 36370 53282 36382
rect 60958 36370 61010 36382
rect 43922 36318 43934 36370
rect 43986 36318 43998 36370
rect 46274 36318 46286 36370
rect 46338 36318 46350 36370
rect 49074 36318 49086 36370
rect 49138 36318 49150 36370
rect 54786 36318 54798 36370
rect 54850 36318 54862 36370
rect 56018 36318 56030 36370
rect 56082 36318 56094 36370
rect 56466 36318 56478 36370
rect 56530 36318 56542 36370
rect 59266 36318 59278 36370
rect 59330 36318 59342 36370
rect 40910 36306 40962 36318
rect 48078 36306 48130 36318
rect 53230 36306 53282 36318
rect 60958 36306 61010 36318
rect 61518 36370 61570 36382
rect 61518 36306 61570 36318
rect 2382 36258 2434 36270
rect 2382 36194 2434 36206
rect 2606 36258 2658 36270
rect 2606 36194 2658 36206
rect 5966 36258 6018 36270
rect 13582 36258 13634 36270
rect 7858 36206 7870 36258
rect 7922 36206 7934 36258
rect 5966 36194 6018 36206
rect 13582 36194 13634 36206
rect 21534 36258 21586 36270
rect 22878 36258 22930 36270
rect 21970 36206 21982 36258
rect 22034 36206 22046 36258
rect 21534 36194 21586 36206
rect 22878 36194 22930 36206
rect 35422 36258 35474 36270
rect 53678 36258 53730 36270
rect 45378 36206 45390 36258
rect 45442 36206 45454 36258
rect 35422 36194 35474 36206
rect 53678 36194 53730 36206
rect 60510 36258 60562 36270
rect 60510 36194 60562 36206
rect 60734 36258 60786 36270
rect 60734 36194 60786 36206
rect 1344 36090 62608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 62608 36090
rect 1344 36004 62608 36038
rect 2046 35922 2098 35934
rect 2046 35858 2098 35870
rect 8878 35922 8930 35934
rect 11454 35922 11506 35934
rect 10994 35870 11006 35922
rect 11058 35870 11070 35922
rect 8878 35858 8930 35870
rect 11454 35858 11506 35870
rect 13022 35922 13074 35934
rect 13022 35858 13074 35870
rect 13134 35922 13186 35934
rect 13134 35858 13186 35870
rect 17502 35922 17554 35934
rect 17502 35858 17554 35870
rect 18286 35922 18338 35934
rect 18286 35858 18338 35870
rect 18398 35922 18450 35934
rect 18398 35858 18450 35870
rect 22430 35922 22482 35934
rect 32510 35922 32562 35934
rect 29138 35870 29150 35922
rect 29202 35870 29214 35922
rect 30594 35870 30606 35922
rect 30658 35870 30670 35922
rect 22430 35858 22482 35870
rect 32510 35858 32562 35870
rect 35198 35922 35250 35934
rect 35198 35858 35250 35870
rect 35422 35922 35474 35934
rect 35422 35858 35474 35870
rect 40126 35922 40178 35934
rect 40126 35858 40178 35870
rect 40238 35922 40290 35934
rect 56702 35922 56754 35934
rect 42914 35870 42926 35922
rect 42978 35870 42990 35922
rect 40238 35858 40290 35870
rect 56702 35858 56754 35870
rect 58382 35922 58434 35934
rect 58382 35858 58434 35870
rect 62190 35922 62242 35934
rect 62190 35858 62242 35870
rect 2382 35810 2434 35822
rect 10110 35810 10162 35822
rect 12798 35810 12850 35822
rect 3378 35758 3390 35810
rect 3442 35758 3454 35810
rect 7298 35758 7310 35810
rect 7362 35758 7374 35810
rect 7970 35758 7982 35810
rect 8034 35758 8046 35810
rect 12562 35758 12574 35810
rect 12626 35758 12638 35810
rect 2382 35746 2434 35758
rect 10110 35746 10162 35758
rect 12798 35746 12850 35758
rect 12910 35810 12962 35822
rect 22990 35810 23042 35822
rect 35086 35810 35138 35822
rect 40014 35810 40066 35822
rect 14130 35758 14142 35810
rect 14194 35758 14206 35810
rect 21074 35758 21086 35810
rect 21138 35758 21150 35810
rect 26002 35758 26014 35810
rect 26066 35758 26078 35810
rect 33842 35758 33854 35810
rect 33906 35758 33918 35810
rect 34178 35758 34190 35810
rect 34242 35758 34254 35810
rect 39778 35758 39790 35810
rect 39842 35758 39854 35810
rect 12910 35746 12962 35758
rect 22990 35746 23042 35758
rect 35086 35746 35138 35758
rect 40014 35746 40066 35758
rect 40350 35810 40402 35822
rect 47630 35810 47682 35822
rect 41122 35758 41134 35810
rect 41186 35758 41198 35810
rect 43698 35758 43710 35810
rect 43762 35758 43774 35810
rect 44258 35758 44270 35810
rect 44322 35758 44334 35810
rect 45042 35758 45054 35810
rect 45106 35758 45118 35810
rect 46834 35758 46846 35810
rect 46898 35758 46910 35810
rect 40350 35746 40402 35758
rect 47630 35746 47682 35758
rect 48750 35810 48802 35822
rect 48750 35746 48802 35758
rect 48862 35810 48914 35822
rect 53330 35758 53342 35810
rect 53394 35758 53406 35810
rect 57362 35758 57374 35810
rect 57426 35758 57438 35810
rect 59602 35758 59614 35810
rect 59666 35758 59678 35810
rect 48862 35746 48914 35758
rect 1934 35698 1986 35710
rect 1934 35634 1986 35646
rect 2158 35698 2210 35710
rect 8542 35698 8594 35710
rect 10670 35698 10722 35710
rect 3490 35646 3502 35698
rect 3554 35646 3566 35698
rect 4722 35646 4734 35698
rect 4786 35646 4798 35698
rect 5954 35646 5966 35698
rect 6018 35646 6030 35698
rect 7074 35646 7086 35698
rect 7138 35646 7150 35698
rect 7746 35646 7758 35698
rect 7810 35646 7822 35698
rect 9762 35646 9774 35698
rect 9826 35646 9838 35698
rect 2158 35634 2210 35646
rect 8542 35634 8594 35646
rect 10670 35634 10722 35646
rect 11342 35698 11394 35710
rect 11342 35634 11394 35646
rect 11566 35698 11618 35710
rect 11566 35634 11618 35646
rect 12014 35698 12066 35710
rect 15150 35698 15202 35710
rect 17390 35698 17442 35710
rect 14578 35646 14590 35698
rect 14642 35646 14654 35698
rect 15362 35646 15374 35698
rect 15426 35646 15438 35698
rect 12014 35634 12066 35646
rect 15150 35634 15202 35646
rect 17390 35634 17442 35646
rect 17614 35698 17666 35710
rect 17614 35634 17666 35646
rect 18062 35698 18114 35710
rect 18062 35634 18114 35646
rect 18510 35698 18562 35710
rect 36654 35698 36706 35710
rect 38782 35698 38834 35710
rect 47854 35698 47906 35710
rect 50094 35698 50146 35710
rect 18834 35646 18846 35698
rect 18898 35646 18910 35698
rect 19618 35646 19630 35698
rect 19682 35646 19694 35698
rect 23202 35646 23214 35698
rect 23266 35646 23278 35698
rect 24098 35646 24110 35698
rect 24162 35646 24174 35698
rect 25218 35646 25230 35698
rect 25282 35646 25294 35698
rect 33170 35646 33182 35698
rect 33234 35646 33246 35698
rect 33506 35646 33518 35698
rect 33570 35646 33582 35698
rect 34402 35646 34414 35698
rect 34466 35646 34478 35698
rect 36306 35646 36318 35698
rect 36370 35646 36382 35698
rect 38546 35646 38558 35698
rect 38610 35646 38622 35698
rect 40898 35646 40910 35698
rect 40962 35646 40974 35698
rect 42018 35646 42030 35698
rect 42082 35646 42094 35698
rect 42354 35646 42366 35698
rect 42418 35646 42430 35698
rect 42802 35646 42814 35698
rect 42866 35646 42878 35698
rect 43474 35646 43486 35698
rect 43538 35646 43550 35698
rect 44482 35646 44494 35698
rect 44546 35646 44558 35698
rect 45378 35646 45390 35698
rect 45442 35646 45454 35698
rect 47170 35646 47182 35698
rect 47234 35646 47246 35698
rect 48178 35646 48190 35698
rect 48242 35646 48254 35698
rect 49298 35646 49310 35698
rect 49362 35646 49374 35698
rect 18510 35634 18562 35646
rect 36654 35634 36706 35646
rect 38782 35634 38834 35646
rect 47854 35634 47906 35646
rect 50094 35634 50146 35646
rect 51886 35698 51938 35710
rect 51886 35634 51938 35646
rect 51998 35698 52050 35710
rect 52210 35646 52222 35698
rect 52274 35646 52286 35698
rect 53218 35646 53230 35698
rect 53282 35646 53294 35698
rect 54450 35646 54462 35698
rect 54514 35646 54526 35698
rect 57250 35646 57262 35698
rect 57314 35646 57326 35698
rect 58818 35646 58830 35698
rect 58882 35646 58894 35698
rect 51998 35634 52050 35646
rect 10446 35586 10498 35598
rect 31950 35586 32002 35598
rect 4274 35534 4286 35586
rect 4338 35534 4350 35586
rect 19954 35534 19966 35586
rect 20018 35534 20030 35586
rect 24434 35534 24446 35586
rect 24498 35534 24510 35586
rect 28130 35534 28142 35586
rect 28194 35534 28206 35586
rect 10446 35522 10498 35534
rect 31950 35522 32002 35534
rect 36542 35586 36594 35598
rect 47742 35586 47794 35598
rect 54014 35586 54066 35598
rect 41458 35534 41470 35586
rect 41522 35534 41534 35586
rect 53554 35534 53566 35586
rect 53618 35534 53630 35586
rect 36542 35522 36594 35534
rect 47742 35522 47794 35534
rect 54014 35522 54066 35534
rect 55470 35586 55522 35598
rect 61730 35534 61742 35586
rect 61794 35534 61806 35586
rect 55470 35522 55522 35534
rect 48862 35474 48914 35486
rect 14354 35422 14366 35474
rect 14418 35422 14430 35474
rect 23538 35422 23550 35474
rect 23602 35422 23614 35474
rect 48862 35410 48914 35422
rect 55694 35474 55746 35486
rect 58046 35474 58098 35486
rect 56018 35422 56030 35474
rect 56082 35422 56094 35474
rect 55694 35410 55746 35422
rect 58046 35410 58098 35422
rect 1344 35306 62608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 62608 35306
rect 1344 35220 62608 35254
rect 3054 35138 3106 35150
rect 3054 35074 3106 35086
rect 5854 35138 5906 35150
rect 5854 35074 5906 35086
rect 13582 35138 13634 35150
rect 13582 35074 13634 35086
rect 13918 35138 13970 35150
rect 13918 35074 13970 35086
rect 23326 35138 23378 35150
rect 44830 35138 44882 35150
rect 40562 35086 40574 35138
rect 40626 35086 40638 35138
rect 23326 35074 23378 35086
rect 44830 35074 44882 35086
rect 44942 35138 44994 35150
rect 44942 35074 44994 35086
rect 45166 35138 45218 35150
rect 45166 35074 45218 35086
rect 45278 35138 45330 35150
rect 50094 35138 50146 35150
rect 49074 35086 49086 35138
rect 49138 35086 49150 35138
rect 45278 35074 45330 35086
rect 50094 35074 50146 35086
rect 53006 35138 53058 35150
rect 53006 35074 53058 35086
rect 53566 35138 53618 35150
rect 53566 35074 53618 35086
rect 53790 35138 53842 35150
rect 53790 35074 53842 35086
rect 55470 35138 55522 35150
rect 55470 35074 55522 35086
rect 55582 35138 55634 35150
rect 55582 35074 55634 35086
rect 61070 35138 61122 35150
rect 61070 35074 61122 35086
rect 61742 35138 61794 35150
rect 61742 35074 61794 35086
rect 22542 35026 22594 35038
rect 4050 34974 4062 35026
rect 4114 34974 4126 35026
rect 22542 34962 22594 34974
rect 28478 35026 28530 35038
rect 37102 35026 37154 35038
rect 31378 34974 31390 35026
rect 31442 34974 31454 35026
rect 34402 34974 34414 35026
rect 34466 34974 34478 35026
rect 43698 34974 43710 35026
rect 43762 34974 43774 35026
rect 51762 34974 51774 35026
rect 51826 34974 51838 35026
rect 28478 34962 28530 34974
rect 37102 34962 37154 34974
rect 6190 34914 6242 34926
rect 7534 34914 7586 34926
rect 2594 34862 2606 34914
rect 2658 34862 2670 34914
rect 4162 34862 4174 34914
rect 4226 34862 4238 34914
rect 4498 34862 4510 34914
rect 4562 34862 4574 34914
rect 6850 34862 6862 34914
rect 6914 34862 6926 34914
rect 6190 34850 6242 34862
rect 7534 34850 7586 34862
rect 7870 34914 7922 34926
rect 7870 34850 7922 34862
rect 7982 34914 8034 34926
rect 8654 34914 8706 34926
rect 8082 34862 8094 34914
rect 8146 34862 8158 34914
rect 7982 34850 8034 34862
rect 8654 34850 8706 34862
rect 9102 34914 9154 34926
rect 9102 34850 9154 34862
rect 9326 34914 9378 34926
rect 15262 34914 15314 34926
rect 9650 34862 9662 34914
rect 9714 34862 9726 34914
rect 9986 34862 9998 34914
rect 10050 34862 10062 34914
rect 11106 34862 11118 34914
rect 11170 34862 11182 34914
rect 11778 34862 11790 34914
rect 11842 34862 11854 34914
rect 14578 34862 14590 34914
rect 14642 34862 14654 34914
rect 9326 34850 9378 34862
rect 15262 34850 15314 34862
rect 15598 34914 15650 34926
rect 15598 34850 15650 34862
rect 15822 34914 15874 34926
rect 15822 34850 15874 34862
rect 16046 34914 16098 34926
rect 16046 34850 16098 34862
rect 17390 34914 17442 34926
rect 22206 34914 22258 34926
rect 21522 34862 21534 34914
rect 21586 34862 21598 34914
rect 17390 34850 17442 34862
rect 22206 34850 22258 34862
rect 23102 34914 23154 34926
rect 28142 34914 28194 34926
rect 23650 34862 23662 34914
rect 23714 34862 23726 34914
rect 23986 34862 23998 34914
rect 24050 34862 24062 34914
rect 25106 34862 25118 34914
rect 25170 34862 25182 34914
rect 25666 34862 25678 34914
rect 25730 34862 25742 34914
rect 27122 34862 27134 34914
rect 27186 34862 27198 34914
rect 23102 34850 23154 34862
rect 28142 34850 28194 34862
rect 28366 34914 28418 34926
rect 28366 34850 28418 34862
rect 28590 34914 28642 34926
rect 33966 34914 34018 34926
rect 30146 34862 30158 34914
rect 30210 34862 30222 34914
rect 31826 34862 31838 34914
rect 31890 34862 31902 34914
rect 33058 34862 33070 34914
rect 33122 34862 33134 34914
rect 28590 34850 28642 34862
rect 33966 34850 34018 34862
rect 35086 34914 35138 34926
rect 42254 34914 42306 34926
rect 48190 34914 48242 34926
rect 50430 34914 50482 34926
rect 54238 34914 54290 34926
rect 37538 34862 37550 34914
rect 37602 34862 37614 34914
rect 38098 34862 38110 34914
rect 38162 34862 38174 34914
rect 39554 34862 39566 34914
rect 39618 34862 39630 34914
rect 41010 34862 41022 34914
rect 41074 34862 41086 34914
rect 42802 34862 42814 34914
rect 42866 34862 42878 34914
rect 43586 34862 43598 34914
rect 43650 34862 43662 34914
rect 46274 34862 46286 34914
rect 46338 34862 46350 34914
rect 47730 34862 47742 34914
rect 47794 34862 47806 34914
rect 49186 34862 49198 34914
rect 49250 34862 49262 34914
rect 51202 34862 51214 34914
rect 51266 34862 51278 34914
rect 51650 34862 51662 34914
rect 51714 34862 51726 34914
rect 35086 34850 35138 34862
rect 42254 34850 42306 34862
rect 48190 34850 48242 34862
rect 50430 34850 50482 34862
rect 54238 34850 54290 34862
rect 55806 34914 55858 34926
rect 60734 34914 60786 34926
rect 56914 34862 56926 34914
rect 56978 34862 56990 34914
rect 58034 34862 58046 34914
rect 58098 34862 58110 34914
rect 58258 34862 58270 34914
rect 58322 34862 58334 34914
rect 59826 34862 59838 34914
rect 59890 34862 59902 34914
rect 55806 34850 55858 34862
rect 60734 34850 60786 34862
rect 12798 34802 12850 34814
rect 15374 34802 15426 34814
rect 20750 34802 20802 34814
rect 27582 34802 27634 34814
rect 2370 34750 2382 34802
rect 2434 34750 2446 34802
rect 6738 34750 6750 34802
rect 6802 34750 6814 34802
rect 14466 34750 14478 34802
rect 14530 34750 14542 34802
rect 18274 34750 18286 34802
rect 18338 34750 18350 34802
rect 21410 34750 21422 34802
rect 21474 34750 21486 34802
rect 24882 34750 24894 34802
rect 24946 34750 24958 34802
rect 12798 34738 12850 34750
rect 15374 34738 15426 34750
rect 20750 34738 20802 34750
rect 27582 34738 27634 34750
rect 29150 34802 29202 34814
rect 53230 34802 53282 34814
rect 30258 34750 30270 34802
rect 30322 34750 30334 34802
rect 35522 34750 35534 34802
rect 35586 34750 35598 34802
rect 35858 34750 35870 34802
rect 35922 34750 35934 34802
rect 40562 34750 40574 34802
rect 40626 34750 40638 34802
rect 42914 34750 42926 34802
rect 42978 34750 42990 34802
rect 50978 34750 50990 34802
rect 51042 34750 51054 34802
rect 29150 34738 29202 34750
rect 53230 34738 53282 34750
rect 53342 34802 53394 34814
rect 53342 34738 53394 34750
rect 54574 34802 54626 34814
rect 55918 34802 55970 34814
rect 54674 34750 54686 34802
rect 54738 34750 54750 34802
rect 54574 34738 54626 34750
rect 55918 34738 55970 34750
rect 56590 34802 56642 34814
rect 60510 34802 60562 34814
rect 57138 34750 57150 34802
rect 57202 34750 57214 34802
rect 59602 34750 59614 34802
rect 59666 34750 59678 34802
rect 56590 34738 56642 34750
rect 60510 34738 60562 34750
rect 61966 34802 62018 34814
rect 61966 34738 62018 34750
rect 1934 34690 1986 34702
rect 1934 34626 1986 34638
rect 3390 34690 3442 34702
rect 8318 34690 8370 34702
rect 4722 34638 4734 34690
rect 4786 34638 4798 34690
rect 3390 34626 3442 34638
rect 8318 34626 8370 34638
rect 8766 34690 8818 34702
rect 8766 34626 8818 34638
rect 10110 34690 10162 34702
rect 10110 34626 10162 34638
rect 12686 34690 12738 34702
rect 16718 34690 16770 34702
rect 16370 34638 16382 34690
rect 16434 34638 16446 34690
rect 12686 34626 12738 34638
rect 16718 34626 16770 34638
rect 16830 34690 16882 34702
rect 16830 34626 16882 34638
rect 16942 34690 16994 34702
rect 16942 34626 16994 34638
rect 20078 34690 20130 34702
rect 20078 34626 20130 34638
rect 20414 34690 20466 34702
rect 20414 34626 20466 34638
rect 29262 34690 29314 34702
rect 29262 34626 29314 34638
rect 29374 34690 29426 34702
rect 41918 34690 41970 34702
rect 35074 34638 35086 34690
rect 35138 34638 35150 34690
rect 37762 34638 37774 34690
rect 37826 34638 37838 34690
rect 29374 34626 29426 34638
rect 41918 34626 41970 34638
rect 45838 34690 45890 34702
rect 45838 34626 45890 34638
rect 54350 34690 54402 34702
rect 54350 34626 54402 34638
rect 54462 34690 54514 34702
rect 54462 34626 54514 34638
rect 56254 34690 56306 34702
rect 61394 34638 61406 34690
rect 61458 34638 61470 34690
rect 56254 34626 56306 34638
rect 1344 34522 62608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 62608 34522
rect 1344 34436 62608 34470
rect 2494 34354 2546 34366
rect 2494 34290 2546 34302
rect 11790 34354 11842 34366
rect 11790 34290 11842 34302
rect 12910 34354 12962 34366
rect 17278 34354 17330 34366
rect 15474 34302 15486 34354
rect 15538 34302 15550 34354
rect 12910 34290 12962 34302
rect 17278 34290 17330 34302
rect 22654 34354 22706 34366
rect 27358 34354 27410 34366
rect 24658 34302 24670 34354
rect 24722 34302 24734 34354
rect 22654 34290 22706 34302
rect 27358 34290 27410 34302
rect 32398 34354 32450 34366
rect 32398 34290 32450 34302
rect 36206 34354 36258 34366
rect 36206 34290 36258 34302
rect 40350 34354 40402 34366
rect 40350 34290 40402 34302
rect 41470 34354 41522 34366
rect 41470 34290 41522 34302
rect 41694 34354 41746 34366
rect 41694 34290 41746 34302
rect 42702 34354 42754 34366
rect 42702 34290 42754 34302
rect 43598 34354 43650 34366
rect 55246 34354 55298 34366
rect 46834 34302 46846 34354
rect 46898 34302 46910 34354
rect 47730 34302 47742 34354
rect 47794 34302 47806 34354
rect 43598 34290 43650 34302
rect 55246 34290 55298 34302
rect 59166 34354 59218 34366
rect 59166 34290 59218 34302
rect 12126 34242 12178 34254
rect 17502 34242 17554 34254
rect 18398 34242 18450 34254
rect 3378 34190 3390 34242
rect 3442 34190 3454 34242
rect 10770 34190 10782 34242
rect 10834 34190 10846 34242
rect 13458 34190 13470 34242
rect 13522 34190 13534 34242
rect 14018 34190 14030 34242
rect 14082 34190 14094 34242
rect 15026 34190 15038 34242
rect 15090 34190 15102 34242
rect 15362 34190 15374 34242
rect 15426 34190 15438 34242
rect 18162 34190 18174 34242
rect 18226 34190 18238 34242
rect 12126 34178 12178 34190
rect 17502 34178 17554 34190
rect 18398 34178 18450 34190
rect 18510 34242 18562 34254
rect 28254 34242 28306 34254
rect 32174 34242 32226 34254
rect 19842 34190 19854 34242
rect 19906 34190 19918 34242
rect 29810 34190 29822 34242
rect 29874 34190 29886 34242
rect 30370 34190 30382 34242
rect 30434 34190 30446 34242
rect 18510 34178 18562 34190
rect 28254 34178 28306 34190
rect 32174 34178 32226 34190
rect 32286 34242 32338 34254
rect 35982 34242 36034 34254
rect 33394 34190 33406 34242
rect 33458 34190 33470 34242
rect 32286 34178 32338 34190
rect 35982 34178 36034 34190
rect 36094 34242 36146 34254
rect 36094 34178 36146 34190
rect 36654 34242 36706 34254
rect 41022 34242 41074 34254
rect 38882 34190 38894 34242
rect 38946 34190 38958 34242
rect 36654 34178 36706 34190
rect 41022 34178 41074 34190
rect 42590 34242 42642 34254
rect 42590 34178 42642 34190
rect 43150 34242 43202 34254
rect 48750 34242 48802 34254
rect 45378 34190 45390 34242
rect 45442 34190 45454 34242
rect 43150 34178 43202 34190
rect 48750 34178 48802 34190
rect 49086 34242 49138 34254
rect 49086 34178 49138 34190
rect 52110 34242 52162 34254
rect 52110 34178 52162 34190
rect 55918 34242 55970 34254
rect 61742 34242 61794 34254
rect 57026 34190 57038 34242
rect 57090 34190 57102 34242
rect 60722 34190 60734 34242
rect 60786 34190 60798 34242
rect 55918 34178 55970 34190
rect 61742 34178 61794 34190
rect 2158 34130 2210 34142
rect 2158 34066 2210 34078
rect 2382 34130 2434 34142
rect 2382 34066 2434 34078
rect 2718 34130 2770 34142
rect 15822 34130 15874 34142
rect 3154 34078 3166 34130
rect 3218 34078 3230 34130
rect 4722 34078 4734 34130
rect 4786 34078 4798 34130
rect 6066 34078 6078 34130
rect 6130 34078 6142 34130
rect 6850 34078 6862 34130
rect 6914 34078 6926 34130
rect 7634 34078 7646 34130
rect 7698 34078 7710 34130
rect 2718 34066 2770 34078
rect 15822 34066 15874 34078
rect 16270 34130 16322 34142
rect 16270 34066 16322 34078
rect 17614 34130 17666 34142
rect 17614 34066 17666 34078
rect 18734 34130 18786 34142
rect 18734 34066 18786 34078
rect 22990 34130 23042 34142
rect 22990 34066 23042 34078
rect 23438 34130 23490 34142
rect 23438 34066 23490 34078
rect 26126 34130 26178 34142
rect 26126 34066 26178 34078
rect 27694 34130 27746 34142
rect 27694 34066 27746 34078
rect 29598 34130 29650 34142
rect 29598 34066 29650 34078
rect 31054 34130 31106 34142
rect 32510 34130 32562 34142
rect 36318 34130 36370 34142
rect 39678 34130 39730 34142
rect 31714 34078 31726 34130
rect 31778 34078 31790 34130
rect 35634 34078 35646 34130
rect 35698 34078 35710 34130
rect 36866 34078 36878 34130
rect 36930 34078 36942 34130
rect 37762 34078 37774 34130
rect 37826 34078 37838 34130
rect 38994 34078 39006 34130
rect 39058 34078 39070 34130
rect 31054 34066 31106 34078
rect 32510 34066 32562 34078
rect 36318 34066 36370 34078
rect 39678 34066 39730 34078
rect 39902 34130 39954 34142
rect 39902 34066 39954 34078
rect 40798 34130 40850 34142
rect 40798 34066 40850 34078
rect 41134 34130 41186 34142
rect 42814 34130 42866 34142
rect 41906 34078 41918 34130
rect 41970 34078 41982 34130
rect 42130 34078 42142 34130
rect 42194 34078 42206 34130
rect 41134 34066 41186 34078
rect 42814 34066 42866 34078
rect 44158 34130 44210 34142
rect 44158 34066 44210 34078
rect 46510 34130 46562 34142
rect 49870 34130 49922 34142
rect 47170 34078 47182 34130
rect 47234 34078 47246 34130
rect 46510 34066 46562 34078
rect 49870 34066 49922 34078
rect 49982 34130 50034 34142
rect 53342 34130 53394 34142
rect 51874 34078 51886 34130
rect 51938 34078 51950 34130
rect 52322 34078 52334 34130
rect 52386 34078 52398 34130
rect 49982 34066 50034 34078
rect 53342 34066 53394 34078
rect 53790 34130 53842 34142
rect 53790 34066 53842 34078
rect 54014 34130 54066 34142
rect 54014 34066 54066 34078
rect 54462 34130 54514 34142
rect 54910 34130 54962 34142
rect 62078 34130 62130 34142
rect 54674 34078 54686 34130
rect 54738 34078 54750 34130
rect 55010 34078 55022 34130
rect 55074 34078 55086 34130
rect 55570 34078 55582 34130
rect 55634 34078 55646 34130
rect 54462 34066 54514 34078
rect 54910 34066 54962 34078
rect 62078 34066 62130 34078
rect 8990 34018 9042 34030
rect 4050 33966 4062 34018
rect 4114 33966 4126 34018
rect 7522 33966 7534 34018
rect 7586 33966 7598 34018
rect 8990 33954 9042 33966
rect 16830 34018 16882 34030
rect 24110 34018 24162 34030
rect 18386 33966 18398 34018
rect 18450 33966 18462 34018
rect 23202 33966 23214 34018
rect 23266 33966 23278 34018
rect 16830 33954 16882 33966
rect 24110 33954 24162 33966
rect 24334 34018 24386 34030
rect 26462 34018 26514 34030
rect 25666 33966 25678 34018
rect 25730 33966 25742 34018
rect 24334 33954 24386 33966
rect 26462 33954 26514 33966
rect 28142 34018 28194 34030
rect 28142 33954 28194 33966
rect 28814 34018 28866 34030
rect 28814 33954 28866 33966
rect 30830 34018 30882 34030
rect 30830 33954 30882 33966
rect 31390 34018 31442 34030
rect 31390 33954 31442 33966
rect 38222 34018 38274 34030
rect 38222 33954 38274 33966
rect 38334 34018 38386 34030
rect 46286 34018 46338 34030
rect 42242 33966 42254 34018
rect 42306 33966 42318 34018
rect 38334 33954 38386 33966
rect 46286 33954 46338 33966
rect 48078 34018 48130 34030
rect 48078 33954 48130 33966
rect 53566 34018 53618 34030
rect 53566 33954 53618 33966
rect 53902 34018 53954 34030
rect 53902 33954 53954 33966
rect 7086 33906 7138 33918
rect 7086 33842 7138 33854
rect 9662 33906 9714 33918
rect 9662 33842 9714 33854
rect 13246 33906 13298 33918
rect 22878 33906 22930 33918
rect 21410 33854 21422 33906
rect 21474 33854 21486 33906
rect 13246 33842 13298 33854
rect 22878 33842 22930 33854
rect 23662 33906 23714 33918
rect 23662 33842 23714 33854
rect 26686 33906 26738 33918
rect 28030 33906 28082 33918
rect 27010 33854 27022 33906
rect 27074 33854 27086 33906
rect 26686 33842 26738 33854
rect 28030 33842 28082 33854
rect 29262 33906 29314 33918
rect 29262 33842 29314 33854
rect 35310 33906 35362 33918
rect 48190 33906 48242 33918
rect 39330 33854 39342 33906
rect 39394 33854 39406 33906
rect 35310 33842 35362 33854
rect 48190 33842 48242 33854
rect 55582 33906 55634 33918
rect 55582 33842 55634 33854
rect 58830 33906 58882 33918
rect 58830 33842 58882 33854
rect 59614 33906 59666 33918
rect 59614 33842 59666 33854
rect 1344 33738 62608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 62608 33738
rect 1344 33652 62608 33686
rect 1934 33570 1986 33582
rect 1934 33506 1986 33518
rect 17726 33570 17778 33582
rect 37102 33570 37154 33582
rect 25442 33518 25454 33570
rect 25506 33518 25518 33570
rect 30370 33518 30382 33570
rect 30434 33518 30446 33570
rect 17726 33506 17778 33518
rect 37102 33506 37154 33518
rect 37326 33570 37378 33582
rect 37326 33506 37378 33518
rect 37886 33570 37938 33582
rect 46062 33570 46114 33582
rect 40562 33518 40574 33570
rect 40626 33518 40638 33570
rect 37886 33506 37938 33518
rect 46062 33506 46114 33518
rect 50766 33570 50818 33582
rect 53118 33570 53170 33582
rect 51314 33518 51326 33570
rect 51378 33518 51390 33570
rect 50766 33506 50818 33518
rect 53118 33506 53170 33518
rect 54462 33570 54514 33582
rect 54462 33506 54514 33518
rect 10558 33458 10610 33470
rect 14142 33458 14194 33470
rect 7074 33406 7086 33458
rect 7138 33406 7150 33458
rect 12786 33406 12798 33458
rect 12850 33406 12862 33458
rect 10558 33394 10610 33406
rect 14142 33394 14194 33406
rect 19070 33458 19122 33470
rect 19070 33394 19122 33406
rect 21646 33458 21698 33470
rect 21646 33394 21698 33406
rect 21982 33458 22034 33470
rect 21982 33394 22034 33406
rect 28254 33458 28306 33470
rect 32734 33458 32786 33470
rect 53454 33458 53506 33470
rect 30034 33406 30046 33458
rect 30098 33406 30110 33458
rect 36194 33406 36206 33458
rect 36258 33406 36270 33458
rect 47394 33406 47406 33458
rect 47458 33406 47470 33458
rect 55458 33406 55470 33458
rect 55522 33406 55534 33458
rect 28254 33394 28306 33406
rect 32734 33394 32786 33406
rect 53454 33394 53506 33406
rect 11006 33346 11058 33358
rect 14030 33346 14082 33358
rect 20526 33346 20578 33358
rect 4050 33294 4062 33346
rect 4114 33294 4126 33346
rect 5618 33294 5630 33346
rect 5682 33294 5694 33346
rect 6178 33294 6190 33346
rect 6242 33294 6254 33346
rect 7186 33294 7198 33346
rect 7250 33294 7262 33346
rect 10210 33294 10222 33346
rect 10274 33294 10286 33346
rect 12002 33294 12014 33346
rect 12066 33294 12078 33346
rect 12338 33294 12350 33346
rect 12402 33294 12414 33346
rect 14578 33294 14590 33346
rect 14642 33294 14654 33346
rect 16034 33294 16046 33346
rect 16098 33294 16110 33346
rect 16818 33294 16830 33346
rect 16882 33294 16894 33346
rect 18610 33294 18622 33346
rect 18674 33294 18686 33346
rect 19282 33294 19294 33346
rect 19346 33294 19358 33346
rect 11006 33282 11058 33294
rect 14030 33282 14082 33294
rect 20526 33282 20578 33294
rect 20750 33346 20802 33358
rect 20750 33282 20802 33294
rect 22542 33346 22594 33358
rect 29262 33346 29314 33358
rect 33070 33346 33122 33358
rect 35086 33346 35138 33358
rect 25218 33294 25230 33346
rect 25282 33294 25294 33346
rect 29922 33294 29934 33346
rect 29986 33294 29998 33346
rect 31714 33294 31726 33346
rect 31778 33294 31790 33346
rect 34402 33294 34414 33346
rect 34466 33294 34478 33346
rect 22542 33282 22594 33294
rect 29262 33282 29314 33294
rect 33070 33282 33122 33294
rect 35086 33282 35138 33294
rect 35422 33346 35474 33358
rect 40126 33346 40178 33358
rect 44158 33346 44210 33358
rect 45726 33346 45778 33358
rect 53902 33346 53954 33358
rect 38210 33294 38222 33346
rect 38274 33294 38286 33346
rect 39666 33294 39678 33346
rect 39730 33294 39742 33346
rect 41346 33294 41358 33346
rect 41410 33294 41422 33346
rect 45042 33294 45054 33346
rect 45106 33294 45118 33346
rect 51538 33294 51550 33346
rect 51602 33294 51614 33346
rect 52770 33294 52782 33346
rect 52834 33294 52846 33346
rect 53330 33294 53342 33346
rect 53394 33294 53406 33346
rect 35422 33282 35474 33294
rect 40126 33282 40178 33294
rect 44158 33282 44210 33294
rect 45726 33282 45778 33294
rect 53902 33282 53954 33294
rect 54126 33346 54178 33358
rect 58158 33346 58210 33358
rect 61742 33346 61794 33358
rect 55010 33294 55022 33346
rect 55074 33294 55086 33346
rect 56466 33294 56478 33346
rect 56530 33294 56542 33346
rect 56802 33294 56814 33346
rect 56866 33294 56878 33346
rect 60722 33294 60734 33346
rect 60786 33294 60798 33346
rect 54126 33282 54178 33294
rect 58158 33282 58210 33294
rect 61742 33282 61794 33294
rect 11342 33234 11394 33246
rect 21870 33234 21922 33246
rect 26014 33234 26066 33246
rect 33294 33234 33346 33246
rect 6850 33182 6862 33234
rect 6914 33182 6926 33234
rect 9538 33182 9550 33234
rect 9602 33182 9614 33234
rect 10770 33182 10782 33234
rect 10834 33182 10846 33234
rect 12674 33182 12686 33234
rect 12738 33182 12750 33234
rect 17378 33182 17390 33234
rect 17442 33182 17454 33234
rect 18498 33182 18510 33234
rect 18562 33182 18574 33234
rect 19058 33182 19070 33234
rect 19122 33182 19134 33234
rect 23202 33182 23214 33234
rect 23266 33182 23278 33234
rect 25778 33182 25790 33234
rect 25842 33182 25854 33234
rect 27122 33182 27134 33234
rect 27186 33182 27198 33234
rect 11342 33170 11394 33182
rect 21870 33170 21922 33182
rect 26014 33170 26066 33182
rect 33294 33170 33346 33182
rect 33742 33234 33794 33246
rect 35870 33234 35922 33246
rect 34290 33182 34302 33234
rect 34354 33182 34366 33234
rect 33742 33170 33794 33182
rect 35870 33170 35922 33182
rect 37662 33234 37714 33246
rect 53566 33234 53618 33246
rect 61966 33234 62018 33246
rect 42242 33182 42254 33234
rect 42306 33182 42318 33234
rect 45154 33182 45166 33234
rect 45218 33182 45230 33234
rect 46834 33182 46846 33234
rect 46898 33182 46910 33234
rect 48738 33182 48750 33234
rect 48802 33182 48814 33234
rect 59378 33182 59390 33234
rect 59442 33182 59454 33234
rect 60498 33182 60510 33234
rect 60562 33182 60574 33234
rect 37662 33170 37714 33182
rect 53566 33170 53618 33182
rect 61966 33170 62018 33182
rect 5182 33122 5234 33134
rect 5182 33058 5234 33070
rect 7758 33122 7810 33134
rect 7758 33058 7810 33070
rect 10222 33122 10274 33134
rect 10222 33058 10274 33070
rect 11454 33122 11506 33134
rect 11454 33058 11506 33070
rect 13806 33122 13858 33134
rect 13806 33058 13858 33070
rect 14254 33122 14306 33134
rect 22094 33122 22146 33134
rect 20178 33070 20190 33122
rect 20242 33070 20254 33122
rect 14254 33058 14306 33070
rect 22094 33058 22146 33070
rect 25006 33122 25058 33134
rect 33854 33122 33906 33134
rect 25554 33070 25566 33122
rect 25618 33070 25630 33122
rect 25006 33058 25058 33070
rect 33854 33058 33906 33070
rect 36094 33122 36146 33134
rect 36094 33058 36146 33070
rect 36990 33122 37042 33134
rect 36990 33058 37042 33070
rect 46510 33122 46562 33134
rect 46510 33058 46562 33070
rect 47854 33122 47906 33134
rect 61394 33070 61406 33122
rect 61458 33070 61470 33122
rect 47854 33058 47906 33070
rect 1344 32954 62608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 62608 32954
rect 1344 32868 62608 32902
rect 8990 32786 9042 32798
rect 8990 32722 9042 32734
rect 9886 32786 9938 32798
rect 22766 32786 22818 32798
rect 11218 32734 11230 32786
rect 11282 32734 11294 32786
rect 9886 32722 9938 32734
rect 22766 32722 22818 32734
rect 23438 32786 23490 32798
rect 23438 32722 23490 32734
rect 28254 32786 28306 32798
rect 28254 32722 28306 32734
rect 28814 32786 28866 32798
rect 34526 32786 34578 32798
rect 30482 32734 30494 32786
rect 30546 32734 30558 32786
rect 31490 32734 31502 32786
rect 31554 32734 31566 32786
rect 33506 32734 33518 32786
rect 33570 32734 33582 32786
rect 28814 32722 28866 32734
rect 34526 32722 34578 32734
rect 38334 32786 38386 32798
rect 38334 32722 38386 32734
rect 38446 32786 38498 32798
rect 38446 32722 38498 32734
rect 38782 32786 38834 32798
rect 40238 32786 40290 32798
rect 39778 32734 39790 32786
rect 39842 32734 39854 32786
rect 38782 32722 38834 32734
rect 40238 32722 40290 32734
rect 40462 32786 40514 32798
rect 48974 32786 49026 32798
rect 43586 32734 43598 32786
rect 43650 32734 43662 32786
rect 40462 32722 40514 32734
rect 48974 32722 49026 32734
rect 49198 32786 49250 32798
rect 57486 32786 57538 32798
rect 54450 32734 54462 32786
rect 54514 32734 54526 32786
rect 56018 32734 56030 32786
rect 56082 32734 56094 32786
rect 49198 32722 49250 32734
rect 57486 32722 57538 32734
rect 58382 32786 58434 32798
rect 58382 32722 58434 32734
rect 16270 32674 16322 32686
rect 22878 32674 22930 32686
rect 27918 32674 27970 32686
rect 38558 32674 38610 32686
rect 44158 32674 44210 32686
rect 48862 32674 48914 32686
rect 57934 32674 57986 32686
rect 3042 32622 3054 32674
rect 3106 32622 3118 32674
rect 4834 32622 4846 32674
rect 4898 32622 4910 32674
rect 15586 32622 15598 32674
rect 15650 32622 15662 32674
rect 16594 32622 16606 32674
rect 16658 32622 16670 32674
rect 17938 32622 17950 32674
rect 18002 32622 18014 32674
rect 22194 32622 22206 32674
rect 22258 32622 22270 32674
rect 24546 32622 24558 32674
rect 24610 32622 24622 32674
rect 36194 32622 36206 32674
rect 36258 32622 36270 32674
rect 42354 32622 42366 32674
rect 42418 32622 42430 32674
rect 44482 32622 44494 32674
rect 44546 32622 44558 32674
rect 46050 32622 46062 32674
rect 46114 32622 46126 32674
rect 51986 32622 51998 32674
rect 52050 32622 52062 32674
rect 61618 32622 61630 32674
rect 61682 32622 61694 32674
rect 16270 32610 16322 32622
rect 22878 32610 22930 32622
rect 27918 32610 27970 32622
rect 38558 32610 38610 32622
rect 44158 32610 44210 32622
rect 48862 32610 48914 32622
rect 57934 32610 57986 32622
rect 4062 32562 4114 32574
rect 9550 32562 9602 32574
rect 2034 32510 2046 32562
rect 2098 32510 2110 32562
rect 2370 32510 2382 32562
rect 2434 32510 2446 32562
rect 3602 32510 3614 32562
rect 3666 32510 3678 32562
rect 5842 32510 5854 32562
rect 5906 32510 5918 32562
rect 6178 32510 6190 32562
rect 6242 32510 6254 32562
rect 7522 32510 7534 32562
rect 7586 32510 7598 32562
rect 4062 32498 4114 32510
rect 9550 32498 9602 32510
rect 9886 32562 9938 32574
rect 9886 32498 9938 32510
rect 10222 32562 10274 32574
rect 14814 32562 14866 32574
rect 16046 32562 16098 32574
rect 19070 32562 19122 32574
rect 21534 32562 21586 32574
rect 29374 32562 29426 32574
rect 13346 32510 13358 32562
rect 13410 32510 13422 32562
rect 15474 32510 15486 32562
rect 15538 32510 15550 32562
rect 16482 32510 16494 32562
rect 16546 32510 16558 32562
rect 17602 32510 17614 32562
rect 17666 32510 17678 32562
rect 19282 32510 19294 32562
rect 19346 32510 19358 32562
rect 22306 32510 22318 32562
rect 22370 32510 22382 32562
rect 24434 32510 24446 32562
rect 24498 32510 24510 32562
rect 26226 32510 26238 32562
rect 26290 32510 26302 32562
rect 26450 32510 26462 32562
rect 26514 32510 26526 32562
rect 27010 32510 27022 32562
rect 27074 32510 27086 32562
rect 28914 32510 28926 32562
rect 28978 32510 28990 32562
rect 10222 32498 10274 32510
rect 14814 32498 14866 32510
rect 16046 32498 16098 32510
rect 19070 32498 19122 32510
rect 21534 32498 21586 32510
rect 29374 32498 29426 32510
rect 31838 32562 31890 32574
rect 31838 32498 31890 32510
rect 32062 32562 32114 32574
rect 32062 32498 32114 32510
rect 33070 32562 33122 32574
rect 37774 32562 37826 32574
rect 33282 32510 33294 32562
rect 33346 32510 33358 32562
rect 33842 32510 33854 32562
rect 33906 32510 33918 32562
rect 33070 32498 33122 32510
rect 37774 32498 37826 32510
rect 37998 32562 38050 32574
rect 37998 32498 38050 32510
rect 39454 32562 39506 32574
rect 39454 32498 39506 32510
rect 40126 32562 40178 32574
rect 58494 32562 58546 32574
rect 60510 32562 60562 32574
rect 41682 32510 41694 32562
rect 41746 32510 41758 32562
rect 42242 32510 42254 32562
rect 42306 32510 42318 32562
rect 42690 32510 42702 32562
rect 42754 32510 42766 32562
rect 44706 32510 44718 32562
rect 44770 32510 44782 32562
rect 45378 32510 45390 32562
rect 45442 32510 45454 32562
rect 50530 32510 50542 32562
rect 50594 32510 50606 32562
rect 51202 32510 51214 32562
rect 51266 32510 51278 32562
rect 54674 32510 54686 32562
rect 54738 32510 54750 32562
rect 57026 32510 57038 32562
rect 57090 32510 57102 32562
rect 57698 32510 57710 32562
rect 57762 32510 57774 32562
rect 60162 32510 60174 32562
rect 60226 32510 60238 32562
rect 61058 32510 61070 32562
rect 61122 32510 61134 32562
rect 40126 32498 40178 32510
rect 58494 32498 58546 32510
rect 60510 32498 60562 32510
rect 12574 32450 12626 32462
rect 14030 32450 14082 32462
rect 2258 32398 2270 32450
rect 2322 32398 2334 32450
rect 4498 32398 4510 32450
rect 4562 32398 4574 32450
rect 8530 32398 8542 32450
rect 8594 32398 8606 32450
rect 13122 32398 13134 32450
rect 13186 32398 13198 32450
rect 12574 32386 12626 32398
rect 14030 32386 14082 32398
rect 16158 32450 16210 32462
rect 32510 32450 32562 32462
rect 26674 32398 26686 32450
rect 26738 32398 26750 32450
rect 16158 32386 16210 32398
rect 32510 32386 32562 32398
rect 37102 32450 37154 32462
rect 37102 32386 37154 32398
rect 39230 32450 39282 32462
rect 49534 32450 49586 32462
rect 55470 32450 55522 32462
rect 48178 32398 48190 32450
rect 48242 32398 48254 32450
rect 50418 32398 50430 32450
rect 50482 32398 50494 32450
rect 54114 32398 54126 32450
rect 54178 32398 54190 32450
rect 56914 32398 56926 32450
rect 56978 32398 56990 32450
rect 39230 32386 39282 32398
rect 49534 32386 49586 32398
rect 55470 32386 55522 32398
rect 14478 32338 14530 32350
rect 21198 32338 21250 32350
rect 17490 32286 17502 32338
rect 17554 32286 17566 32338
rect 14478 32274 14530 32286
rect 21198 32274 21250 32286
rect 23774 32338 23826 32350
rect 43934 32338 43986 32350
rect 50206 32338 50258 32350
rect 33618 32286 33630 32338
rect 33682 32286 33694 32338
rect 37426 32286 37438 32338
rect 37490 32286 37502 32338
rect 49522 32286 49534 32338
rect 49586 32335 49598 32338
rect 49970 32335 49982 32338
rect 49586 32289 49982 32335
rect 49586 32286 49598 32289
rect 49970 32286 49982 32289
rect 50034 32286 50046 32338
rect 23774 32274 23826 32286
rect 43934 32274 43986 32286
rect 50206 32274 50258 32286
rect 55694 32338 55746 32350
rect 55694 32274 55746 32286
rect 57374 32338 57426 32350
rect 57374 32274 57426 32286
rect 58382 32338 58434 32350
rect 61282 32286 61294 32338
rect 61346 32286 61358 32338
rect 58382 32274 58434 32286
rect 1344 32170 62608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 62608 32170
rect 1344 32084 62608 32118
rect 10222 32002 10274 32014
rect 2706 31950 2718 32002
rect 2770 31950 2782 32002
rect 3490 31950 3502 32002
rect 3554 31950 3566 32002
rect 6178 31950 6190 32002
rect 6242 31950 6254 32002
rect 10222 31938 10274 31950
rect 17502 32002 17554 32014
rect 17502 31938 17554 31950
rect 22318 32002 22370 32014
rect 34190 32002 34242 32014
rect 33282 31950 33294 32002
rect 33346 31950 33358 32002
rect 22318 31938 22370 31950
rect 34190 31938 34242 31950
rect 51326 32002 51378 32014
rect 51326 31938 51378 31950
rect 52110 32002 52162 32014
rect 52110 31938 52162 31950
rect 57150 32002 57202 32014
rect 61058 31950 61070 32002
rect 61122 31950 61134 32002
rect 57150 31938 57202 31950
rect 1934 31890 1986 31902
rect 4734 31890 4786 31902
rect 3714 31838 3726 31890
rect 3778 31838 3790 31890
rect 1934 31826 1986 31838
rect 4734 31826 4786 31838
rect 8542 31890 8594 31902
rect 8542 31826 8594 31838
rect 9214 31890 9266 31902
rect 9214 31826 9266 31838
rect 9886 31890 9938 31902
rect 28366 31890 28418 31902
rect 19506 31838 19518 31890
rect 19570 31838 19582 31890
rect 28018 31838 28030 31890
rect 28082 31838 28094 31890
rect 9886 31826 9938 31838
rect 28366 31826 28418 31838
rect 34974 31890 35026 31902
rect 34974 31826 35026 31838
rect 36430 31890 36482 31902
rect 36430 31826 36482 31838
rect 43598 31890 43650 31902
rect 43598 31826 43650 31838
rect 45726 31890 45778 31902
rect 51998 31890 52050 31902
rect 47170 31838 47182 31890
rect 47234 31838 47246 31890
rect 45726 31826 45778 31838
rect 51998 31826 52050 31838
rect 57486 31890 57538 31902
rect 57486 31826 57538 31838
rect 2158 31778 2210 31790
rect 4846 31778 4898 31790
rect 2370 31726 2382 31778
rect 2434 31726 2446 31778
rect 2706 31726 2718 31778
rect 2770 31726 2782 31778
rect 2158 31714 2210 31726
rect 4846 31714 4898 31726
rect 5630 31778 5682 31790
rect 5630 31714 5682 31726
rect 5966 31778 6018 31790
rect 7086 31778 7138 31790
rect 6178 31726 6190 31778
rect 6242 31726 6254 31778
rect 5966 31714 6018 31726
rect 7086 31714 7138 31726
rect 7982 31778 8034 31790
rect 7982 31714 8034 31726
rect 8318 31778 8370 31790
rect 9438 31778 9490 31790
rect 14366 31778 14418 31790
rect 8978 31726 8990 31778
rect 9042 31726 9054 31778
rect 11554 31726 11566 31778
rect 11618 31726 11630 31778
rect 13458 31726 13470 31778
rect 13522 31726 13534 31778
rect 8318 31714 8370 31726
rect 9438 31714 9490 31726
rect 14366 31714 14418 31726
rect 14478 31778 14530 31790
rect 14478 31714 14530 31726
rect 16494 31778 16546 31790
rect 17838 31778 17890 31790
rect 16818 31726 16830 31778
rect 16882 31726 16894 31778
rect 16494 31714 16546 31726
rect 17838 31714 17890 31726
rect 18062 31778 18114 31790
rect 22542 31778 22594 31790
rect 18498 31726 18510 31778
rect 18562 31726 18574 31778
rect 20178 31726 20190 31778
rect 20242 31726 20254 31778
rect 21522 31726 21534 31778
rect 21586 31726 21598 31778
rect 18062 31714 18114 31726
rect 22542 31714 22594 31726
rect 22766 31778 22818 31790
rect 22766 31714 22818 31726
rect 22878 31778 22930 31790
rect 22878 31714 22930 31726
rect 23998 31778 24050 31790
rect 28478 31778 28530 31790
rect 34302 31778 34354 31790
rect 24322 31726 24334 31778
rect 24386 31726 24398 31778
rect 25218 31726 25230 31778
rect 25282 31726 25294 31778
rect 33394 31726 33406 31778
rect 33458 31726 33470 31778
rect 23998 31714 24050 31726
rect 28478 31714 28530 31726
rect 34302 31714 34354 31726
rect 34750 31778 34802 31790
rect 34750 31714 34802 31726
rect 35534 31778 35586 31790
rect 35534 31714 35586 31726
rect 35758 31778 35810 31790
rect 37998 31778 38050 31790
rect 35970 31726 35982 31778
rect 36034 31726 36046 31778
rect 35758 31714 35810 31726
rect 37998 31714 38050 31726
rect 38222 31778 38274 31790
rect 46622 31778 46674 31790
rect 53678 31778 53730 31790
rect 61406 31778 61458 31790
rect 38546 31726 38558 31778
rect 38610 31726 38622 31778
rect 39666 31726 39678 31778
rect 39730 31726 39742 31778
rect 40674 31726 40686 31778
rect 40738 31726 40750 31778
rect 45266 31726 45278 31778
rect 45330 31726 45342 31778
rect 47506 31726 47518 31778
rect 47570 31726 47582 31778
rect 54562 31726 54574 31778
rect 54626 31726 54638 31778
rect 60498 31726 60510 31778
rect 60562 31726 60574 31778
rect 38222 31714 38274 31726
rect 46622 31714 46674 31726
rect 53678 31714 53730 31726
rect 61406 31714 61458 31726
rect 61630 31778 61682 31790
rect 61630 31714 61682 31726
rect 3278 31666 3330 31678
rect 3278 31602 3330 31614
rect 6862 31666 6914 31678
rect 6862 31602 6914 31614
rect 7422 31666 7474 31678
rect 7422 31602 7474 31614
rect 7758 31666 7810 31678
rect 7758 31602 7810 31614
rect 8094 31666 8146 31678
rect 8094 31602 8146 31614
rect 11118 31666 11170 31678
rect 12686 31666 12738 31678
rect 23102 31666 23154 31678
rect 11778 31614 11790 31666
rect 11842 31614 11854 31666
rect 18722 31614 18734 31666
rect 18786 31614 18798 31666
rect 21298 31614 21310 31666
rect 21362 31614 21374 31666
rect 11118 31602 11170 31614
rect 12686 31602 12738 31614
rect 23102 31602 23154 31614
rect 23550 31666 23602 31678
rect 23550 31602 23602 31614
rect 23662 31666 23714 31678
rect 23662 31602 23714 31614
rect 24446 31666 24498 31678
rect 24446 31602 24498 31614
rect 24558 31666 24610 31678
rect 29710 31666 29762 31678
rect 32734 31666 32786 31678
rect 34526 31666 34578 31678
rect 25890 31614 25902 31666
rect 25954 31614 25966 31666
rect 31154 31614 31166 31666
rect 31218 31614 31230 31666
rect 32946 31614 32958 31666
rect 33010 31614 33022 31666
rect 24558 31602 24610 31614
rect 29710 31602 29762 31614
rect 32734 31602 32786 31614
rect 34526 31602 34578 31614
rect 36318 31666 36370 31678
rect 36318 31602 36370 31614
rect 37326 31666 37378 31678
rect 37326 31602 37378 31614
rect 37662 31666 37714 31678
rect 44158 31666 44210 31678
rect 61854 31666 61906 31678
rect 38882 31614 38894 31666
rect 38946 31614 38958 31666
rect 41122 31614 41134 31666
rect 41186 31614 41198 31666
rect 42242 31614 42254 31666
rect 42306 31614 42318 31666
rect 49298 31614 49310 31666
rect 49362 31614 49374 31666
rect 52994 31614 53006 31666
rect 53058 31614 53070 31666
rect 53330 31614 53342 31666
rect 53394 31614 53406 31666
rect 55346 31614 55358 31666
rect 55410 31614 55422 31666
rect 58818 31614 58830 31666
rect 58882 31614 58894 31666
rect 37662 31602 37714 31614
rect 44158 31602 44210 31614
rect 61854 31602 61906 31614
rect 2942 31554 2994 31566
rect 2942 31490 2994 31502
rect 6414 31554 6466 31566
rect 6414 31490 6466 31502
rect 6974 31554 7026 31566
rect 6974 31490 7026 31502
rect 9102 31554 9154 31566
rect 9102 31490 9154 31502
rect 10110 31554 10162 31566
rect 10110 31490 10162 31502
rect 11006 31554 11058 31566
rect 11006 31490 11058 31502
rect 12126 31554 12178 31566
rect 12126 31490 12178 31502
rect 23326 31554 23378 31566
rect 23326 31490 23378 31502
rect 24670 31554 24722 31566
rect 24670 31490 24722 31502
rect 29150 31554 29202 31566
rect 29150 31490 29202 31502
rect 30270 31554 30322 31566
rect 30270 31490 30322 31502
rect 32286 31554 32338 31566
rect 32286 31490 32338 31502
rect 33518 31554 33570 31566
rect 33518 31490 33570 31502
rect 35870 31554 35922 31566
rect 35870 31490 35922 31502
rect 46062 31554 46114 31566
rect 46062 31490 46114 31502
rect 48190 31554 48242 31566
rect 48190 31490 48242 31502
rect 52670 31554 52722 31566
rect 52670 31490 52722 31502
rect 54462 31554 54514 31566
rect 54462 31490 54514 31502
rect 59950 31554 60002 31566
rect 59950 31490 60002 31502
rect 61518 31554 61570 31566
rect 61518 31490 61570 31502
rect 1344 31386 62608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 62608 31386
rect 1344 31300 62608 31334
rect 2270 31218 2322 31230
rect 2270 31154 2322 31166
rect 2494 31218 2546 31230
rect 2494 31154 2546 31166
rect 6974 31218 7026 31230
rect 6974 31154 7026 31166
rect 7646 31218 7698 31230
rect 7646 31154 7698 31166
rect 8542 31218 8594 31230
rect 8542 31154 8594 31166
rect 8766 31218 8818 31230
rect 11678 31218 11730 31230
rect 10546 31166 10558 31218
rect 10610 31166 10622 31218
rect 8766 31154 8818 31166
rect 11678 31154 11730 31166
rect 12574 31218 12626 31230
rect 12574 31154 12626 31166
rect 12798 31218 12850 31230
rect 12798 31154 12850 31166
rect 15150 31218 15202 31230
rect 16270 31218 16322 31230
rect 15150 31154 15202 31166
rect 15374 31162 15426 31174
rect 2046 31106 2098 31118
rect 2046 31042 2098 31054
rect 2158 31106 2210 31118
rect 2158 31042 2210 31054
rect 5630 31106 5682 31118
rect 5630 31042 5682 31054
rect 13358 31106 13410 31118
rect 13358 31042 13410 31054
rect 14814 31106 14866 31118
rect 16270 31154 16322 31166
rect 16382 31218 16434 31230
rect 16382 31154 16434 31166
rect 17502 31218 17554 31230
rect 20190 31218 20242 31230
rect 18834 31166 18846 31218
rect 18898 31166 18910 31218
rect 17502 31154 17554 31166
rect 20190 31154 20242 31166
rect 20862 31218 20914 31230
rect 20862 31154 20914 31166
rect 24558 31218 24610 31230
rect 24558 31154 24610 31166
rect 27694 31218 27746 31230
rect 27694 31154 27746 31166
rect 30382 31218 30434 31230
rect 31166 31218 31218 31230
rect 30706 31166 30718 31218
rect 30770 31166 30782 31218
rect 30382 31154 30434 31166
rect 31166 31154 31218 31166
rect 33070 31218 33122 31230
rect 33854 31218 33906 31230
rect 33394 31166 33406 31218
rect 33458 31166 33470 31218
rect 33070 31154 33122 31166
rect 33854 31154 33906 31166
rect 37550 31218 37602 31230
rect 37550 31154 37602 31166
rect 39678 31218 39730 31230
rect 39678 31154 39730 31166
rect 41470 31218 41522 31230
rect 44830 31218 44882 31230
rect 43698 31166 43710 31218
rect 43762 31166 43774 31218
rect 41470 31154 41522 31166
rect 44830 31154 44882 31166
rect 46510 31218 46562 31230
rect 46510 31154 46562 31166
rect 47070 31218 47122 31230
rect 47070 31154 47122 31166
rect 47630 31218 47682 31230
rect 47630 31154 47682 31166
rect 50542 31218 50594 31230
rect 50542 31154 50594 31166
rect 51102 31218 51154 31230
rect 51102 31154 51154 31166
rect 57598 31218 57650 31230
rect 57598 31154 57650 31166
rect 15374 31098 15426 31110
rect 15486 31106 15538 31118
rect 24110 31106 24162 31118
rect 47742 31106 47794 31118
rect 53902 31106 53954 31118
rect 56030 31106 56082 31118
rect 14814 31042 14866 31054
rect 15698 31054 15710 31106
rect 15762 31054 15774 31106
rect 17826 31054 17838 31106
rect 17890 31054 17902 31106
rect 22530 31054 22542 31106
rect 22594 31054 22606 31106
rect 23090 31054 23102 31106
rect 23154 31054 23166 31106
rect 29922 31054 29934 31106
rect 29986 31054 29998 31106
rect 32162 31054 32174 31106
rect 32226 31054 32238 31106
rect 38770 31054 38782 31106
rect 38834 31054 38846 31106
rect 45602 31054 45614 31106
rect 45666 31054 45678 31106
rect 45938 31054 45950 31106
rect 46002 31054 46014 31106
rect 49298 31054 49310 31106
rect 49362 31054 49374 31106
rect 51762 31054 51774 31106
rect 51826 31054 51838 31106
rect 52434 31054 52446 31106
rect 52498 31054 52510 31106
rect 53554 31054 53566 31106
rect 53618 31054 53630 31106
rect 54226 31054 54238 31106
rect 54290 31054 54302 31106
rect 15486 31042 15538 31054
rect 24110 31042 24162 31054
rect 47742 31042 47794 31054
rect 53902 31042 53954 31054
rect 56030 31042 56082 31054
rect 56590 31106 56642 31118
rect 58146 31054 58158 31106
rect 58210 31054 58222 31106
rect 58706 31054 58718 31106
rect 58770 31054 58782 31106
rect 56590 31042 56642 31054
rect 3726 30994 3778 31006
rect 7870 30994 7922 31006
rect 3154 30942 3166 30994
rect 3218 30942 3230 30994
rect 5954 30942 5966 30994
rect 6018 30942 6030 30994
rect 3726 30930 3778 30942
rect 7870 30930 7922 30942
rect 8094 30994 8146 31006
rect 8094 30930 8146 30942
rect 8318 30994 8370 31006
rect 8318 30930 8370 30942
rect 8878 30994 8930 31006
rect 8878 30930 8930 30942
rect 12462 30994 12514 31006
rect 12462 30930 12514 30942
rect 12910 30994 12962 31006
rect 12910 30930 12962 30942
rect 13694 30994 13746 31006
rect 13694 30930 13746 30942
rect 16494 30994 16546 31006
rect 16494 30930 16546 30942
rect 16942 30994 16994 31006
rect 16942 30930 16994 30942
rect 20750 30994 20802 31006
rect 20750 30930 20802 30942
rect 21086 30994 21138 31006
rect 21086 30930 21138 30942
rect 21310 30994 21362 31006
rect 23550 30994 23602 31006
rect 22082 30942 22094 30994
rect 22146 30942 22158 30994
rect 23202 30942 23214 30994
rect 23266 30942 23278 30994
rect 21310 30930 21362 30942
rect 23550 30930 23602 30942
rect 23886 30994 23938 31006
rect 23886 30930 23938 30942
rect 24334 30994 24386 31006
rect 24334 30930 24386 30942
rect 24670 30994 24722 31006
rect 24670 30930 24722 30942
rect 25790 30994 25842 31006
rect 25790 30930 25842 30942
rect 27358 30994 27410 31006
rect 31502 30994 31554 31006
rect 41806 30994 41858 31006
rect 46174 30994 46226 31006
rect 28914 30942 28926 30994
rect 28978 30942 28990 30994
rect 29586 30942 29598 30994
rect 29650 30942 29662 30994
rect 32274 30942 32286 30994
rect 32338 30942 32350 30994
rect 27358 30930 27410 30942
rect 31502 30930 31554 30942
rect 34178 30930 34190 30982
rect 34242 30930 34254 30982
rect 42242 30942 42254 30994
rect 42306 30942 42318 30994
rect 41806 30930 41858 30942
rect 46174 30930 46226 30942
rect 47406 30994 47458 31006
rect 51438 30994 51490 31006
rect 48178 30942 48190 30994
rect 48242 30942 48254 30994
rect 47406 30930 47458 30942
rect 51438 30930 51490 30942
rect 52110 30994 52162 31006
rect 52110 30930 52162 30942
rect 54574 30994 54626 31006
rect 54574 30930 54626 30942
rect 55806 30994 55858 31006
rect 55806 30930 55858 30942
rect 56814 30994 56866 31006
rect 56814 30930 56866 30942
rect 57262 30994 57314 31006
rect 57262 30930 57314 30942
rect 57934 30994 57986 31006
rect 59602 30942 59614 30994
rect 59666 30942 59678 30994
rect 57934 30930 57986 30942
rect 3838 30882 3890 30894
rect 3838 30818 3890 30830
rect 6862 30882 6914 30894
rect 6862 30818 6914 30830
rect 7758 30882 7810 30894
rect 22430 30882 22482 30894
rect 15922 30830 15934 30882
rect 15986 30830 15998 30882
rect 7758 30818 7810 30830
rect 22430 30818 22482 30830
rect 23662 30882 23714 30894
rect 23662 30818 23714 30830
rect 26126 30882 26178 30894
rect 27806 30882 27858 30894
rect 40910 30882 40962 30894
rect 53230 30882 53282 30894
rect 27010 30830 27022 30882
rect 27074 30830 27086 30882
rect 28690 30830 28702 30882
rect 28754 30830 28766 30882
rect 34962 30830 34974 30882
rect 35026 30830 35038 30882
rect 37090 30830 37102 30882
rect 37154 30830 37166 30882
rect 40114 30830 40126 30882
rect 40178 30830 40190 30882
rect 47730 30830 47742 30882
rect 47794 30830 47806 30882
rect 52994 30830 53006 30882
rect 53058 30830 53070 30882
rect 26126 30818 26178 30830
rect 27806 30818 27858 30830
rect 40910 30818 40962 30830
rect 53230 30818 53282 30830
rect 55022 30882 55074 30894
rect 55022 30818 55074 30830
rect 57038 30882 57090 30894
rect 57038 30818 57090 30830
rect 59278 30882 59330 30894
rect 59278 30818 59330 30830
rect 61966 30882 62018 30894
rect 61966 30818 62018 30830
rect 25678 30770 25730 30782
rect 55470 30770 55522 30782
rect 14578 30718 14590 30770
rect 14642 30718 14654 30770
rect 29474 30718 29486 30770
rect 29538 30718 29550 30770
rect 25678 30706 25730 30718
rect 55470 30706 55522 30718
rect 1344 30602 62608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 62608 30602
rect 1344 30516 62608 30550
rect 15150 30434 15202 30446
rect 4946 30382 4958 30434
rect 5010 30382 5022 30434
rect 15150 30370 15202 30382
rect 19518 30434 19570 30446
rect 43934 30434 43986 30446
rect 24658 30382 24670 30434
rect 24722 30382 24734 30434
rect 32050 30382 32062 30434
rect 32114 30382 32126 30434
rect 43250 30382 43262 30434
rect 43314 30382 43326 30434
rect 19518 30370 19570 30382
rect 43934 30370 43986 30382
rect 50878 30434 50930 30446
rect 56690 30382 56702 30434
rect 56754 30382 56766 30434
rect 50878 30370 50930 30382
rect 34302 30322 34354 30334
rect 4610 30270 4622 30322
rect 4674 30270 4686 30322
rect 10658 30270 10670 30322
rect 10722 30270 10734 30322
rect 16706 30270 16718 30322
rect 16770 30270 16782 30322
rect 25218 30270 25230 30322
rect 25282 30270 25294 30322
rect 30930 30270 30942 30322
rect 30994 30270 31006 30322
rect 39330 30270 39342 30322
rect 39394 30270 39406 30322
rect 34302 30258 34354 30270
rect 4734 30210 4786 30222
rect 4734 30146 4786 30158
rect 5742 30210 5794 30222
rect 5742 30146 5794 30158
rect 6078 30210 6130 30222
rect 6078 30146 6130 30158
rect 7310 30210 7362 30222
rect 11230 30210 11282 30222
rect 7746 30158 7758 30210
rect 7810 30158 7822 30210
rect 7310 30146 7362 30158
rect 11230 30146 11282 30158
rect 11566 30210 11618 30222
rect 11566 30146 11618 30158
rect 12798 30210 12850 30222
rect 12798 30146 12850 30158
rect 13806 30210 13858 30222
rect 19854 30210 19906 30222
rect 26014 30210 26066 30222
rect 14242 30158 14254 30210
rect 14306 30158 14318 30210
rect 15026 30158 15038 30210
rect 15090 30158 15102 30210
rect 16594 30158 16606 30210
rect 16658 30158 16670 30210
rect 20290 30158 20302 30210
rect 20354 30158 20366 30210
rect 21410 30158 21422 30210
rect 21474 30158 21486 30210
rect 22642 30158 22654 30210
rect 22706 30158 22718 30210
rect 24546 30158 24558 30210
rect 24610 30158 24622 30210
rect 13806 30146 13858 30158
rect 19854 30146 19906 30158
rect 26014 30146 26066 30158
rect 28478 30210 28530 30222
rect 34190 30210 34242 30222
rect 29698 30158 29710 30210
rect 29762 30158 29774 30210
rect 31154 30158 31166 30210
rect 31218 30158 31230 30210
rect 28478 30146 28530 30158
rect 34190 30146 34242 30158
rect 34414 30210 34466 30222
rect 34974 30210 35026 30222
rect 34738 30158 34750 30210
rect 34802 30158 34814 30210
rect 34414 30146 34466 30158
rect 34974 30146 35026 30158
rect 35646 30210 35698 30222
rect 35646 30146 35698 30158
rect 36094 30210 36146 30222
rect 37662 30210 37714 30222
rect 37202 30158 37214 30210
rect 37266 30158 37278 30210
rect 36094 30146 36146 30158
rect 37662 30146 37714 30158
rect 38558 30210 38610 30222
rect 44158 30210 44210 30222
rect 51214 30210 51266 30222
rect 54462 30210 54514 30222
rect 41458 30158 41470 30210
rect 41522 30158 41534 30210
rect 43026 30158 43038 30210
rect 43090 30158 43102 30210
rect 48626 30158 48638 30210
rect 48690 30158 48702 30210
rect 49410 30158 49422 30210
rect 49474 30158 49486 30210
rect 51874 30158 51886 30210
rect 51938 30158 51950 30210
rect 38558 30146 38610 30158
rect 44158 30146 44210 30158
rect 51214 30146 51266 30158
rect 54462 30146 54514 30158
rect 55358 30210 55410 30222
rect 55358 30146 55410 30158
rect 56030 30210 56082 30222
rect 61518 30210 61570 30222
rect 56466 30158 56478 30210
rect 56530 30158 56542 30210
rect 56914 30158 56926 30210
rect 56978 30158 56990 30210
rect 57362 30158 57374 30210
rect 57426 30158 57438 30210
rect 56030 30146 56082 30158
rect 61518 30146 61570 30158
rect 7422 30098 7474 30110
rect 11342 30098 11394 30110
rect 13022 30098 13074 30110
rect 20750 30098 20802 30110
rect 41918 30098 41970 30110
rect 55582 30098 55634 30110
rect 2258 30046 2270 30098
rect 2322 30046 2334 30098
rect 6290 30046 6302 30098
rect 6354 30046 6366 30098
rect 6626 30046 6638 30098
rect 6690 30046 6702 30098
rect 8530 30046 8542 30098
rect 8594 30046 8606 30098
rect 12114 30046 12126 30098
rect 12178 30046 12190 30098
rect 12338 30046 12350 30098
rect 12402 30046 12414 30098
rect 15586 30046 15598 30098
rect 15650 30046 15662 30098
rect 18946 30046 18958 30098
rect 19010 30046 19022 30098
rect 19282 30046 19294 30098
rect 19346 30046 19358 30098
rect 23874 30046 23886 30098
rect 23938 30046 23950 30098
rect 29922 30046 29934 30098
rect 29986 30046 29998 30098
rect 47618 30046 47630 30098
rect 47682 30046 47694 30098
rect 49746 30046 49758 30098
rect 49810 30046 49822 30098
rect 51986 30046 51998 30098
rect 52050 30046 52062 30098
rect 53330 30046 53342 30098
rect 53394 30046 53406 30098
rect 7422 30034 7474 30046
rect 11342 30034 11394 30046
rect 13022 30034 13074 30046
rect 20750 30034 20802 30046
rect 41918 30034 41970 30046
rect 55582 30034 55634 30046
rect 61854 30098 61906 30110
rect 61854 30034 61906 30046
rect 62190 30098 62242 30110
rect 62190 30034 62242 30046
rect 3502 29986 3554 29998
rect 3502 29922 3554 29934
rect 20526 29986 20578 29998
rect 20526 29922 20578 29934
rect 20862 29986 20914 29998
rect 20862 29922 20914 29934
rect 25678 29986 25730 29998
rect 25678 29922 25730 29934
rect 26126 29986 26178 29998
rect 26126 29922 26178 29934
rect 26350 29986 26402 29998
rect 33182 29986 33234 29998
rect 27346 29934 27358 29986
rect 27410 29934 27422 29986
rect 26350 29922 26402 29934
rect 33182 29922 33234 29934
rect 33406 29986 33458 29998
rect 33406 29922 33458 29934
rect 33630 29986 33682 29998
rect 33630 29922 33682 29934
rect 35086 29986 35138 29998
rect 35086 29922 35138 29934
rect 35310 29986 35362 29998
rect 35310 29922 35362 29934
rect 35758 29986 35810 29998
rect 35758 29922 35810 29934
rect 35982 29986 36034 29998
rect 35982 29922 36034 29934
rect 37998 29986 38050 29998
rect 37998 29922 38050 29934
rect 38894 29986 38946 29998
rect 40126 29986 40178 29998
rect 39778 29934 39790 29986
rect 39842 29934 39854 29986
rect 38894 29922 38946 29934
rect 40126 29922 40178 29934
rect 40462 29986 40514 29998
rect 42478 29986 42530 29998
rect 45054 29986 45106 29998
rect 47182 29986 47234 29998
rect 40786 29934 40798 29986
rect 40850 29934 40862 29986
rect 43586 29934 43598 29986
rect 43650 29934 43662 29986
rect 46050 29934 46062 29986
rect 46114 29934 46126 29986
rect 40462 29922 40514 29934
rect 42478 29922 42530 29934
rect 45054 29922 45106 29934
rect 47182 29922 47234 29934
rect 50542 29986 50594 29998
rect 50542 29922 50594 29934
rect 55022 29986 55074 29998
rect 55022 29922 55074 29934
rect 55806 29986 55858 29998
rect 59838 29986 59890 29998
rect 58706 29934 58718 29986
rect 58770 29934 58782 29986
rect 55806 29922 55858 29934
rect 59838 29922 59890 29934
rect 60510 29986 60562 29998
rect 60510 29922 60562 29934
rect 60622 29986 60674 29998
rect 60622 29922 60674 29934
rect 60734 29986 60786 29998
rect 60734 29922 60786 29934
rect 60958 29986 61010 29998
rect 60958 29922 61010 29934
rect 1344 29818 62608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 62608 29818
rect 1344 29732 62608 29766
rect 9886 29650 9938 29662
rect 14142 29650 14194 29662
rect 7970 29598 7982 29650
rect 8034 29598 8046 29650
rect 12338 29598 12350 29650
rect 12402 29598 12414 29650
rect 9886 29586 9938 29598
rect 14142 29586 14194 29598
rect 15822 29650 15874 29662
rect 15822 29586 15874 29598
rect 16382 29650 16434 29662
rect 16382 29586 16434 29598
rect 25566 29650 25618 29662
rect 25566 29586 25618 29598
rect 25790 29650 25842 29662
rect 25790 29586 25842 29598
rect 31950 29650 32002 29662
rect 31950 29586 32002 29598
rect 32398 29650 32450 29662
rect 36654 29650 36706 29662
rect 33394 29598 33406 29650
rect 33458 29598 33470 29650
rect 32398 29586 32450 29598
rect 36654 29586 36706 29598
rect 38446 29650 38498 29662
rect 38446 29586 38498 29598
rect 41470 29650 41522 29662
rect 43822 29650 43874 29662
rect 42354 29598 42366 29650
rect 42418 29598 42430 29650
rect 41470 29586 41522 29598
rect 43822 29586 43874 29598
rect 46958 29650 47010 29662
rect 49298 29598 49310 29650
rect 49362 29598 49374 29650
rect 46958 29586 47010 29598
rect 15710 29538 15762 29550
rect 3826 29486 3838 29538
rect 3890 29486 3902 29538
rect 5506 29486 5518 29538
rect 5570 29486 5582 29538
rect 7858 29486 7870 29538
rect 7922 29486 7934 29538
rect 10770 29486 10782 29538
rect 10834 29486 10846 29538
rect 15026 29486 15038 29538
rect 15090 29486 15102 29538
rect 15710 29474 15762 29486
rect 16494 29538 16546 29550
rect 16494 29474 16546 29486
rect 17950 29538 18002 29550
rect 17950 29474 18002 29486
rect 25454 29538 25506 29550
rect 25454 29474 25506 29486
rect 28814 29538 28866 29550
rect 34526 29538 34578 29550
rect 31266 29486 31278 29538
rect 31330 29486 31342 29538
rect 33282 29486 33294 29538
rect 33346 29486 33358 29538
rect 33842 29486 33854 29538
rect 33906 29486 33918 29538
rect 28814 29474 28866 29486
rect 34526 29474 34578 29486
rect 36542 29538 36594 29550
rect 36542 29474 36594 29486
rect 38110 29538 38162 29550
rect 38110 29474 38162 29486
rect 39006 29538 39058 29550
rect 55918 29538 55970 29550
rect 48066 29486 48078 29538
rect 48130 29486 48142 29538
rect 50194 29486 50206 29538
rect 50258 29486 50270 29538
rect 52322 29486 52334 29538
rect 52386 29486 52398 29538
rect 39006 29474 39058 29486
rect 55918 29474 55970 29486
rect 56702 29538 56754 29550
rect 58370 29486 58382 29538
rect 58434 29486 58446 29538
rect 61282 29486 61294 29538
rect 61346 29486 61358 29538
rect 56702 29474 56754 29486
rect 9550 29426 9602 29438
rect 16046 29426 16098 29438
rect 4498 29374 4510 29426
rect 4562 29374 4574 29426
rect 7746 29374 7758 29426
rect 7810 29374 7822 29426
rect 8418 29374 8430 29426
rect 8482 29374 8494 29426
rect 8978 29374 8990 29426
rect 9042 29374 9054 29426
rect 15250 29374 15262 29426
rect 15314 29374 15326 29426
rect 9550 29362 9602 29374
rect 16046 29362 16098 29374
rect 16270 29426 16322 29438
rect 16270 29362 16322 29374
rect 16942 29426 16994 29438
rect 18174 29426 18226 29438
rect 20526 29426 20578 29438
rect 23998 29426 24050 29438
rect 28702 29426 28754 29438
rect 30494 29426 30546 29438
rect 32510 29426 32562 29438
rect 17378 29374 17390 29426
rect 17442 29374 17454 29426
rect 17714 29374 17726 29426
rect 17778 29374 17790 29426
rect 18722 29374 18734 29426
rect 18786 29374 18798 29426
rect 19842 29374 19854 29426
rect 19906 29374 19918 29426
rect 20738 29374 20750 29426
rect 20802 29374 20814 29426
rect 22194 29374 22206 29426
rect 22258 29374 22270 29426
rect 23090 29374 23102 29426
rect 23154 29374 23166 29426
rect 24210 29374 24222 29426
rect 24274 29374 24286 29426
rect 26226 29374 26238 29426
rect 26290 29374 26302 29426
rect 26786 29374 26798 29426
rect 26850 29374 26862 29426
rect 29026 29374 29038 29426
rect 29090 29374 29102 29426
rect 31154 29374 31166 29426
rect 31218 29374 31230 29426
rect 16942 29362 16994 29374
rect 18174 29362 18226 29374
rect 20526 29362 20578 29374
rect 23998 29362 24050 29374
rect 28702 29362 28754 29374
rect 30494 29362 30546 29374
rect 32510 29362 32562 29374
rect 33182 29426 33234 29438
rect 35534 29426 35586 29438
rect 34738 29374 34750 29426
rect 34802 29374 34814 29426
rect 33182 29362 33234 29374
rect 35534 29362 35586 29374
rect 35982 29426 36034 29438
rect 35982 29362 36034 29374
rect 36206 29426 36258 29438
rect 37214 29426 37266 29438
rect 36866 29374 36878 29426
rect 36930 29374 36942 29426
rect 36206 29362 36258 29374
rect 37214 29362 37266 29374
rect 39678 29426 39730 29438
rect 39678 29362 39730 29374
rect 40126 29426 40178 29438
rect 40126 29362 40178 29374
rect 40350 29426 40402 29438
rect 40350 29362 40402 29374
rect 41918 29426 41970 29438
rect 41918 29362 41970 29374
rect 42702 29426 42754 29438
rect 42702 29362 42754 29374
rect 42926 29426 42978 29438
rect 42926 29362 42978 29374
rect 44158 29426 44210 29438
rect 44158 29362 44210 29374
rect 46286 29426 46338 29438
rect 46286 29362 46338 29374
rect 47294 29426 47346 29438
rect 55134 29426 55186 29438
rect 55806 29426 55858 29438
rect 47842 29374 47854 29426
rect 47906 29374 47918 29426
rect 53218 29374 53230 29426
rect 53282 29374 53294 29426
rect 54562 29374 54574 29426
rect 54626 29374 54638 29426
rect 55458 29374 55470 29426
rect 55522 29374 55534 29426
rect 47294 29362 47346 29374
rect 55134 29362 55186 29374
rect 55806 29362 55858 29374
rect 56590 29426 56642 29438
rect 56590 29362 56642 29374
rect 57598 29426 57650 29438
rect 58034 29374 58046 29426
rect 58098 29374 58110 29426
rect 58818 29374 58830 29426
rect 58882 29374 58894 29426
rect 60274 29374 60286 29426
rect 60338 29374 60350 29426
rect 61394 29374 61406 29426
rect 61458 29374 61470 29426
rect 57598 29362 57650 29374
rect 6974 29314 7026 29326
rect 1698 29262 1710 29314
rect 1762 29262 1774 29314
rect 6974 29250 7026 29262
rect 13358 29314 13410 29326
rect 23438 29314 23490 29326
rect 13682 29262 13694 29314
rect 13746 29262 13758 29314
rect 17938 29262 17950 29314
rect 18002 29262 18014 29314
rect 13358 29250 13410 29262
rect 23438 29250 23490 29262
rect 30158 29314 30210 29326
rect 30158 29250 30210 29262
rect 35198 29314 35250 29326
rect 35198 29250 35250 29262
rect 35310 29314 35362 29326
rect 35310 29250 35362 29262
rect 40238 29314 40290 29326
rect 43262 29314 43314 29326
rect 41010 29262 41022 29314
rect 41074 29262 41086 29314
rect 40238 29250 40290 29262
rect 43262 29250 43314 29262
rect 44718 29314 44770 29326
rect 44718 29250 44770 29262
rect 45054 29314 45106 29326
rect 45054 29250 45106 29262
rect 46510 29314 46562 29326
rect 46510 29250 46562 29262
rect 48750 29314 48802 29326
rect 48750 29250 48802 29262
rect 51998 29314 52050 29326
rect 54910 29314 54962 29326
rect 53666 29262 53678 29314
rect 53730 29262 53742 29314
rect 51998 29250 52050 29262
rect 54910 29250 54962 29262
rect 14478 29202 14530 29214
rect 14478 29138 14530 29150
rect 21758 29202 21810 29214
rect 21758 29138 21810 29150
rect 22766 29202 22818 29214
rect 22766 29138 22818 29150
rect 38782 29202 38834 29214
rect 38782 29138 38834 29150
rect 42030 29202 42082 29214
rect 42030 29138 42082 29150
rect 45278 29202 45330 29214
rect 45950 29202 46002 29214
rect 45602 29150 45614 29202
rect 45666 29150 45678 29202
rect 45278 29138 45330 29150
rect 45950 29138 46002 29150
rect 48974 29202 49026 29214
rect 48974 29138 49026 29150
rect 55918 29202 55970 29214
rect 55918 29138 55970 29150
rect 56702 29202 56754 29214
rect 56702 29138 56754 29150
rect 57262 29202 57314 29214
rect 57262 29138 57314 29150
rect 61966 29202 62018 29214
rect 61966 29138 62018 29150
rect 1344 29034 62608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 62608 29034
rect 1344 28948 62608 28982
rect 2382 28866 2434 28878
rect 2382 28802 2434 28814
rect 15598 28866 15650 28878
rect 15598 28802 15650 28814
rect 20302 28866 20354 28878
rect 20302 28802 20354 28814
rect 25006 28866 25058 28878
rect 36430 28866 36482 28878
rect 31042 28814 31054 28866
rect 31106 28814 31118 28866
rect 25006 28802 25058 28814
rect 36430 28802 36482 28814
rect 37326 28866 37378 28878
rect 49870 28866 49922 28878
rect 40674 28814 40686 28866
rect 40738 28814 40750 28866
rect 47058 28814 47070 28866
rect 47122 28814 47134 28866
rect 37326 28802 37378 28814
rect 49870 28802 49922 28814
rect 51326 28866 51378 28878
rect 51326 28802 51378 28814
rect 52782 28866 52834 28878
rect 52782 28802 52834 28814
rect 55358 28866 55410 28878
rect 55358 28802 55410 28814
rect 58158 28866 58210 28878
rect 58158 28802 58210 28814
rect 1710 28754 1762 28766
rect 10558 28754 10610 28766
rect 6962 28702 6974 28754
rect 7026 28702 7038 28754
rect 9090 28702 9102 28754
rect 9154 28702 9166 28754
rect 1710 28690 1762 28702
rect 10558 28690 10610 28702
rect 13806 28754 13858 28766
rect 13806 28690 13858 28702
rect 14702 28754 14754 28766
rect 14702 28690 14754 28702
rect 18958 28754 19010 28766
rect 18958 28690 19010 28702
rect 19742 28754 19794 28766
rect 29150 28754 29202 28766
rect 35198 28754 35250 28766
rect 24546 28702 24558 28754
rect 24610 28702 24622 28754
rect 30482 28702 30494 28754
rect 30546 28702 30558 28754
rect 33058 28702 33070 28754
rect 33122 28702 33134 28754
rect 19742 28690 19794 28702
rect 29150 28690 29202 28702
rect 35198 28690 35250 28702
rect 37214 28754 37266 28766
rect 37214 28690 37266 28702
rect 37774 28754 37826 28766
rect 37774 28690 37826 28702
rect 40126 28754 40178 28766
rect 56254 28754 56306 28766
rect 45714 28702 45726 28754
rect 45778 28702 45790 28754
rect 57138 28702 57150 28754
rect 57202 28702 57214 28754
rect 60722 28702 60734 28754
rect 60786 28702 60798 28754
rect 40126 28690 40178 28702
rect 56254 28690 56306 28702
rect 1822 28642 1874 28654
rect 1822 28578 1874 28590
rect 5966 28642 6018 28654
rect 9774 28642 9826 28654
rect 6178 28590 6190 28642
rect 6242 28590 6254 28642
rect 5966 28578 6018 28590
rect 9774 28578 9826 28590
rect 12798 28642 12850 28654
rect 16942 28642 16994 28654
rect 19070 28642 19122 28654
rect 14130 28590 14142 28642
rect 14194 28590 14206 28642
rect 14354 28590 14366 28642
rect 14418 28590 14430 28642
rect 16370 28590 16382 28642
rect 16434 28590 16446 28642
rect 17266 28590 17278 28642
rect 17330 28590 17342 28642
rect 12798 28578 12850 28590
rect 16942 28578 16994 28590
rect 19070 28578 19122 28590
rect 19518 28642 19570 28654
rect 19518 28578 19570 28590
rect 19966 28642 20018 28654
rect 19966 28578 20018 28590
rect 20862 28642 20914 28654
rect 28478 28642 28530 28654
rect 21746 28590 21758 28642
rect 21810 28590 21822 28642
rect 20862 28578 20914 28590
rect 28478 28578 28530 28590
rect 29710 28642 29762 28654
rect 34974 28642 35026 28654
rect 30370 28590 30382 28642
rect 30434 28590 30446 28642
rect 31154 28590 31166 28642
rect 31218 28590 31230 28642
rect 32946 28590 32958 28642
rect 33010 28590 33022 28642
rect 29710 28578 29762 28590
rect 34974 28578 35026 28590
rect 35534 28642 35586 28654
rect 35534 28578 35586 28590
rect 35758 28642 35810 28654
rect 35758 28578 35810 28590
rect 35982 28642 36034 28654
rect 39790 28642 39842 28654
rect 36978 28590 36990 28642
rect 37042 28590 37054 28642
rect 38210 28590 38222 28642
rect 38274 28590 38286 28642
rect 39218 28590 39230 28642
rect 39282 28590 39294 28642
rect 35982 28578 36034 28590
rect 39790 28578 39842 28590
rect 39902 28642 39954 28654
rect 39902 28578 39954 28590
rect 40350 28642 40402 28654
rect 45166 28642 45218 28654
rect 41458 28590 41470 28642
rect 41522 28590 41534 28642
rect 42690 28590 42702 28642
rect 42754 28590 42766 28642
rect 43922 28590 43934 28642
rect 43986 28590 43998 28642
rect 40350 28578 40402 28590
rect 45166 28578 45218 28590
rect 45390 28642 45442 28654
rect 50990 28642 51042 28654
rect 46722 28590 46734 28642
rect 46786 28590 46798 28642
rect 47058 28590 47070 28642
rect 47122 28590 47134 28642
rect 50530 28590 50542 28642
rect 50594 28590 50606 28642
rect 45390 28578 45442 28590
rect 50990 28578 51042 28590
rect 51774 28642 51826 28654
rect 51774 28578 51826 28590
rect 53118 28642 53170 28654
rect 60510 28642 60562 28654
rect 61630 28642 61682 28654
rect 55010 28590 55022 28642
rect 55074 28590 55086 28642
rect 55570 28590 55582 28642
rect 55634 28590 55646 28642
rect 56578 28590 56590 28642
rect 56642 28590 56654 28642
rect 57362 28590 57374 28642
rect 57426 28590 57438 28642
rect 61170 28590 61182 28642
rect 61234 28590 61246 28642
rect 53118 28578 53170 28590
rect 60510 28578 60562 28590
rect 61630 28578 61682 28590
rect 62190 28642 62242 28654
rect 62190 28578 62242 28590
rect 5630 28530 5682 28542
rect 4386 28478 4398 28530
rect 4450 28478 4462 28530
rect 5630 28466 5682 28478
rect 5742 28530 5794 28542
rect 14814 28530 14866 28542
rect 46062 28530 46114 28542
rect 9426 28478 9438 28530
rect 9490 28478 9502 28530
rect 11330 28478 11342 28530
rect 11394 28478 11406 28530
rect 15810 28478 15822 28530
rect 15874 28478 15886 28530
rect 22418 28478 22430 28530
rect 22482 28478 22494 28530
rect 26226 28478 26238 28530
rect 26290 28478 26302 28530
rect 27794 28478 27806 28530
rect 27858 28478 27870 28530
rect 28354 28478 28366 28530
rect 28418 28478 28430 28530
rect 31714 28478 31726 28530
rect 31778 28478 31790 28530
rect 38322 28478 38334 28530
rect 38386 28478 38398 28530
rect 41346 28478 41358 28530
rect 41410 28478 41422 28530
rect 5742 28466 5794 28478
rect 14814 28466 14866 28478
rect 46062 28466 46114 28478
rect 46510 28530 46562 28542
rect 54350 28530 54402 28542
rect 47954 28478 47966 28530
rect 48018 28478 48030 28530
rect 50194 28478 50206 28530
rect 50258 28478 50270 28530
rect 52098 28478 52110 28530
rect 52162 28478 52174 28530
rect 53330 28478 53342 28530
rect 53394 28478 53406 28530
rect 53890 28478 53902 28530
rect 53954 28478 53966 28530
rect 46510 28466 46562 28478
rect 54350 28466 54402 28478
rect 54686 28530 54738 28542
rect 54686 28466 54738 28478
rect 55806 28530 55858 28542
rect 60846 28530 60898 28542
rect 57698 28478 57710 28530
rect 57762 28478 57774 28530
rect 59266 28478 59278 28530
rect 59330 28478 59342 28530
rect 55806 28466 55858 28478
rect 60846 28466 60898 28478
rect 14590 28418 14642 28430
rect 14590 28354 14642 28366
rect 18846 28418 18898 28430
rect 45838 28418 45890 28430
rect 28018 28366 28030 28418
rect 28082 28366 28094 28418
rect 34626 28366 34638 28418
rect 34690 28366 34702 28418
rect 39106 28366 39118 28418
rect 39170 28366 39182 28418
rect 44818 28366 44830 28418
rect 44882 28366 44894 28418
rect 18846 28354 18898 28366
rect 45838 28354 45890 28366
rect 47294 28418 47346 28430
rect 47294 28354 47346 28366
rect 55022 28418 55074 28430
rect 55022 28354 55074 28366
rect 60734 28418 60786 28430
rect 60734 28354 60786 28366
rect 1344 28250 62608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 62608 28250
rect 1344 28164 62608 28198
rect 3166 28082 3218 28094
rect 2258 28030 2270 28082
rect 2322 28030 2334 28082
rect 3166 28018 3218 28030
rect 4286 28082 4338 28094
rect 4286 28018 4338 28030
rect 6302 28082 6354 28094
rect 21422 28082 21474 28094
rect 7634 28030 7646 28082
rect 7698 28030 7710 28082
rect 10546 28030 10558 28082
rect 10610 28030 10622 28082
rect 6302 28018 6354 28030
rect 21422 28018 21474 28030
rect 21646 28082 21698 28094
rect 21646 28018 21698 28030
rect 22654 28082 22706 28094
rect 22654 28018 22706 28030
rect 24558 28082 24610 28094
rect 24558 28018 24610 28030
rect 25230 28082 25282 28094
rect 25230 28018 25282 28030
rect 27582 28082 27634 28094
rect 27582 28018 27634 28030
rect 31166 28082 31218 28094
rect 31166 28018 31218 28030
rect 31390 28082 31442 28094
rect 31390 28018 31442 28030
rect 32510 28082 32562 28094
rect 32510 28018 32562 28030
rect 33070 28082 33122 28094
rect 33070 28018 33122 28030
rect 33182 28082 33234 28094
rect 33182 28018 33234 28030
rect 33854 28082 33906 28094
rect 33854 28018 33906 28030
rect 34078 28082 34130 28094
rect 34078 28018 34130 28030
rect 36654 28082 36706 28094
rect 36654 28018 36706 28030
rect 37774 28082 37826 28094
rect 37774 28018 37826 28030
rect 38446 28082 38498 28094
rect 38446 28018 38498 28030
rect 38558 28082 38610 28094
rect 38558 28018 38610 28030
rect 38670 28082 38722 28094
rect 48862 28082 48914 28094
rect 43138 28030 43150 28082
rect 43202 28030 43214 28082
rect 38670 28018 38722 28030
rect 48862 28018 48914 28030
rect 54126 28082 54178 28094
rect 54126 28018 54178 28030
rect 56814 28082 56866 28094
rect 56814 28018 56866 28030
rect 56926 28082 56978 28094
rect 61506 28030 61518 28082
rect 61570 28030 61582 28082
rect 56926 28018 56978 28030
rect 4510 27970 4562 27982
rect 3490 27918 3502 27970
rect 3554 27918 3566 27970
rect 4510 27906 4562 27918
rect 4622 27970 4674 27982
rect 4622 27906 4674 27918
rect 5406 27970 5458 27982
rect 5406 27906 5458 27918
rect 11678 27970 11730 27982
rect 13358 27970 13410 27982
rect 12450 27918 12462 27970
rect 12514 27918 12526 27970
rect 11678 27906 11730 27918
rect 13358 27906 13410 27918
rect 14702 27970 14754 27982
rect 23438 27970 23490 27982
rect 16258 27918 16270 27970
rect 16322 27918 16334 27970
rect 14702 27906 14754 27918
rect 23438 27906 23490 27918
rect 24670 27970 24722 27982
rect 24670 27906 24722 27918
rect 26014 27970 26066 27982
rect 26014 27906 26066 27918
rect 26350 27970 26402 27982
rect 32398 27970 32450 27982
rect 28578 27918 28590 27970
rect 28642 27918 28654 27970
rect 26350 27906 26402 27918
rect 32398 27906 32450 27918
rect 34750 27970 34802 27982
rect 34750 27906 34802 27918
rect 34862 27970 34914 27982
rect 52110 27970 52162 27982
rect 57038 27970 57090 27982
rect 40002 27918 40014 27970
rect 40066 27918 40078 27970
rect 41010 27918 41022 27970
rect 41074 27918 41086 27970
rect 44034 27918 44046 27970
rect 44098 27918 44110 27970
rect 47506 27918 47518 27970
rect 47570 27918 47582 27970
rect 50194 27918 50206 27970
rect 50258 27918 50270 27970
rect 52658 27918 52670 27970
rect 52722 27918 52734 27970
rect 55682 27918 55694 27970
rect 55746 27918 55758 27970
rect 34862 27906 34914 27918
rect 52110 27906 52162 27918
rect 57038 27906 57090 27918
rect 2606 27858 2658 27870
rect 22542 27858 22594 27870
rect 1922 27806 1934 27858
rect 1986 27806 1998 27858
rect 3714 27806 3726 27858
rect 3778 27806 3790 27858
rect 4946 27806 4958 27858
rect 5010 27806 5022 27858
rect 5618 27806 5630 27858
rect 5682 27806 5694 27858
rect 12226 27806 12238 27858
rect 12290 27806 12302 27858
rect 13794 27806 13806 27858
rect 13858 27806 13870 27858
rect 14914 27806 14926 27858
rect 14978 27806 14990 27858
rect 15922 27806 15934 27858
rect 15986 27806 15998 27858
rect 17490 27806 17502 27858
rect 17554 27806 17566 27858
rect 18610 27806 18622 27858
rect 18674 27806 18686 27858
rect 19618 27806 19630 27858
rect 19682 27806 19694 27858
rect 20962 27806 20974 27858
rect 21026 27806 21038 27858
rect 21858 27806 21870 27858
rect 21922 27806 21934 27858
rect 22194 27806 22206 27858
rect 22258 27806 22270 27858
rect 2606 27794 2658 27806
rect 22542 27794 22594 27806
rect 22766 27858 22818 27870
rect 22766 27794 22818 27806
rect 23214 27858 23266 27870
rect 24222 27858 24274 27870
rect 23650 27806 23662 27858
rect 23714 27806 23726 27858
rect 23214 27794 23266 27806
rect 24222 27794 24274 27806
rect 24334 27858 24386 27870
rect 25678 27858 25730 27870
rect 33294 27858 33346 27870
rect 34190 27858 34242 27870
rect 25330 27806 25342 27858
rect 25394 27806 25406 27858
rect 26562 27806 26574 27858
rect 26626 27806 26638 27858
rect 26786 27806 26798 27858
rect 26850 27806 26862 27858
rect 27682 27806 27694 27858
rect 27746 27806 27758 27858
rect 30370 27806 30382 27858
rect 30434 27806 30446 27858
rect 31602 27806 31614 27858
rect 31666 27806 31678 27858
rect 31938 27806 31950 27858
rect 32002 27806 32014 27858
rect 33618 27806 33630 27858
rect 33682 27806 33694 27858
rect 24334 27794 24386 27806
rect 25678 27794 25730 27806
rect 33294 27794 33346 27806
rect 34190 27794 34242 27806
rect 35534 27858 35586 27870
rect 35534 27794 35586 27806
rect 35758 27858 35810 27870
rect 35758 27794 35810 27806
rect 35982 27858 36034 27870
rect 37998 27858 38050 27870
rect 42814 27858 42866 27870
rect 46734 27858 46786 27870
rect 51550 27858 51602 27870
rect 36418 27806 36430 27858
rect 36482 27806 36494 27858
rect 37314 27806 37326 27858
rect 37378 27806 37390 27858
rect 37538 27806 37550 27858
rect 37602 27806 37614 27858
rect 40114 27806 40126 27858
rect 40178 27806 40190 27858
rect 41122 27806 41134 27858
rect 41186 27806 41198 27858
rect 42018 27806 42030 27858
rect 42082 27806 42094 27858
rect 44146 27806 44158 27858
rect 44210 27806 44222 27858
rect 45602 27806 45614 27858
rect 45666 27806 45678 27858
rect 47282 27806 47294 27858
rect 47346 27806 47358 27858
rect 35982 27794 36034 27806
rect 37998 27794 38050 27806
rect 42814 27794 42866 27806
rect 46734 27794 46786 27806
rect 51550 27794 51602 27806
rect 51998 27858 52050 27870
rect 51998 27794 52050 27806
rect 52446 27858 52498 27870
rect 53566 27858 53618 27870
rect 58158 27858 58210 27870
rect 59726 27858 59778 27870
rect 52994 27806 53006 27858
rect 53058 27806 53070 27858
rect 54786 27806 54798 27858
rect 54850 27806 54862 27858
rect 55794 27806 55806 27858
rect 55858 27806 55870 27858
rect 57250 27806 57262 27858
rect 57314 27806 57326 27858
rect 57586 27806 57598 27858
rect 57650 27806 57662 27858
rect 58706 27806 58718 27858
rect 58770 27806 58782 27858
rect 52446 27794 52498 27806
rect 53566 27794 53618 27806
rect 58158 27794 58210 27806
rect 59726 27794 59778 27806
rect 9102 27746 9154 27758
rect 16718 27746 16770 27758
rect 31278 27746 31330 27758
rect 4610 27694 4622 27746
rect 4674 27694 4686 27746
rect 14242 27694 14254 27746
rect 14306 27694 14318 27746
rect 16034 27694 16046 27746
rect 16098 27694 16110 27746
rect 18274 27694 18286 27746
rect 18338 27694 18350 27746
rect 20626 27694 20638 27746
rect 20690 27694 20702 27746
rect 21746 27694 21758 27746
rect 21810 27694 21822 27746
rect 9102 27682 9154 27694
rect 16718 27682 16770 27694
rect 31278 27682 31330 27694
rect 37886 27746 37938 27758
rect 37886 27682 37938 27694
rect 41582 27746 41634 27758
rect 41582 27682 41634 27694
rect 41694 27746 41746 27758
rect 48078 27746 48130 27758
rect 43922 27694 43934 27746
rect 43986 27694 43998 27746
rect 41694 27682 41746 27694
rect 48078 27682 48130 27694
rect 51326 27746 51378 27758
rect 51326 27682 51378 27694
rect 52558 27746 52610 27758
rect 52558 27682 52610 27694
rect 52894 27746 52946 27758
rect 52894 27682 52946 27694
rect 55246 27746 55298 27758
rect 55246 27682 55298 27694
rect 55358 27746 55410 27758
rect 55358 27682 55410 27694
rect 13022 27634 13074 27646
rect 13022 27570 13074 27582
rect 16830 27634 16882 27646
rect 26686 27634 26738 27646
rect 25442 27582 25454 27634
rect 25506 27582 25518 27634
rect 16830 27570 16882 27582
rect 26686 27570 26738 27582
rect 36766 27634 36818 27646
rect 36766 27570 36818 27582
rect 39118 27634 39170 27646
rect 39118 27570 39170 27582
rect 39454 27634 39506 27646
rect 39454 27570 39506 27582
rect 46398 27634 46450 27646
rect 46398 27570 46450 27582
rect 51998 27634 52050 27646
rect 51998 27570 52050 27582
rect 58046 27634 58098 27646
rect 60174 27634 60226 27646
rect 59378 27582 59390 27634
rect 59442 27582 59454 27634
rect 58046 27570 58098 27582
rect 60174 27570 60226 27582
rect 1344 27466 62608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 62608 27466
rect 1344 27380 62608 27414
rect 11342 27298 11394 27310
rect 11342 27234 11394 27246
rect 11678 27298 11730 27310
rect 11678 27234 11730 27246
rect 27694 27298 27746 27310
rect 27694 27234 27746 27246
rect 44942 27298 44994 27310
rect 44942 27234 44994 27246
rect 45390 27298 45442 27310
rect 45390 27234 45442 27246
rect 45614 27298 45666 27310
rect 45614 27234 45666 27246
rect 49758 27298 49810 27310
rect 49758 27234 49810 27246
rect 50094 27298 50146 27310
rect 50094 27234 50146 27246
rect 52110 27298 52162 27310
rect 52110 27234 52162 27246
rect 53118 27298 53170 27310
rect 53118 27234 53170 27246
rect 58270 27298 58322 27310
rect 62078 27298 62130 27310
rect 59378 27246 59390 27298
rect 59442 27246 59454 27298
rect 58270 27234 58322 27246
rect 62078 27234 62130 27246
rect 6190 27186 6242 27198
rect 2594 27134 2606 27186
rect 2658 27134 2670 27186
rect 4386 27134 4398 27186
rect 4450 27134 4462 27186
rect 6190 27122 6242 27134
rect 7758 27186 7810 27198
rect 7758 27122 7810 27134
rect 9326 27186 9378 27198
rect 9326 27122 9378 27134
rect 9886 27186 9938 27198
rect 9886 27122 9938 27134
rect 10222 27186 10274 27198
rect 19070 27186 19122 27198
rect 18050 27134 18062 27186
rect 18114 27134 18126 27186
rect 10222 27122 10274 27134
rect 19070 27122 19122 27134
rect 25118 27186 25170 27198
rect 33406 27186 33458 27198
rect 26002 27134 26014 27186
rect 26066 27134 26078 27186
rect 31154 27134 31166 27186
rect 31218 27134 31230 27186
rect 25118 27122 25170 27134
rect 33406 27122 33458 27134
rect 36318 27186 36370 27198
rect 36318 27122 36370 27134
rect 37102 27186 37154 27198
rect 50542 27186 50594 27198
rect 37762 27134 37774 27186
rect 37826 27134 37838 27186
rect 41682 27134 41694 27186
rect 41746 27134 41758 27186
rect 43138 27134 43150 27186
rect 43202 27134 43214 27186
rect 37102 27122 37154 27134
rect 50542 27122 50594 27134
rect 53902 27186 53954 27198
rect 57822 27186 57874 27198
rect 60846 27186 60898 27198
rect 56802 27134 56814 27186
rect 56866 27134 56878 27186
rect 60610 27134 60622 27186
rect 60674 27134 60686 27186
rect 53902 27122 53954 27134
rect 57822 27122 57874 27134
rect 60846 27122 60898 27134
rect 62190 27186 62242 27198
rect 62190 27122 62242 27134
rect 3054 27074 3106 27086
rect 1922 27022 1934 27074
rect 1986 27022 1998 27074
rect 3054 27010 3106 27022
rect 3390 27074 3442 27086
rect 5630 27074 5682 27086
rect 3714 27022 3726 27074
rect 3778 27022 3790 27074
rect 4610 27022 4622 27074
rect 4674 27022 4686 27074
rect 3390 27010 3442 27022
rect 5630 27010 5682 27022
rect 6974 27074 7026 27086
rect 6974 27010 7026 27022
rect 7646 27074 7698 27086
rect 7646 27010 7698 27022
rect 7870 27074 7922 27086
rect 7870 27010 7922 27022
rect 10894 27074 10946 27086
rect 22430 27074 22482 27086
rect 16146 27022 16158 27074
rect 16210 27022 16222 27074
rect 16930 27022 16942 27074
rect 16994 27022 17006 27074
rect 17602 27022 17614 27074
rect 17666 27022 17678 27074
rect 20514 27022 20526 27074
rect 20578 27022 20590 27074
rect 10894 27010 10946 27022
rect 22430 27010 22482 27022
rect 22990 27074 23042 27086
rect 22990 27010 23042 27022
rect 23662 27074 23714 27086
rect 25006 27074 25058 27086
rect 24098 27022 24110 27074
rect 24162 27022 24174 27074
rect 23662 27010 23714 27022
rect 25006 27010 25058 27022
rect 25342 27074 25394 27086
rect 29934 27074 29986 27086
rect 32510 27074 32562 27086
rect 34862 27074 34914 27086
rect 39118 27074 39170 27086
rect 46174 27074 46226 27086
rect 50430 27074 50482 27086
rect 25890 27022 25902 27074
rect 25954 27022 25966 27074
rect 26674 27022 26686 27074
rect 26738 27022 26750 27074
rect 31378 27022 31390 27074
rect 31442 27022 31454 27074
rect 32162 27022 32174 27074
rect 32226 27022 32238 27074
rect 32946 27022 32958 27074
rect 33010 27022 33022 27074
rect 35746 27022 35758 27074
rect 35810 27022 35822 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 38658 27022 38670 27074
rect 38722 27022 38734 27074
rect 40674 27022 40686 27074
rect 40738 27022 40750 27074
rect 41458 27022 41470 27074
rect 41522 27022 41534 27074
rect 47058 27022 47070 27074
rect 47122 27022 47134 27074
rect 25342 27010 25394 27022
rect 29934 27010 29986 27022
rect 32510 27010 32562 27022
rect 34862 27010 34914 27022
rect 39118 27010 39170 27022
rect 46174 27010 46226 27022
rect 50430 27010 50482 27022
rect 50766 27074 50818 27086
rect 50766 27010 50818 27022
rect 50990 27074 51042 27086
rect 50990 27010 51042 27022
rect 51438 27074 51490 27086
rect 51438 27010 51490 27022
rect 51662 27074 51714 27086
rect 51662 27010 51714 27022
rect 51886 27074 51938 27086
rect 53790 27074 53842 27086
rect 52882 27022 52894 27074
rect 52946 27022 52958 27074
rect 53442 27022 53454 27074
rect 53506 27022 53518 27074
rect 51886 27010 51938 27022
rect 53790 27010 53842 27022
rect 54574 27074 54626 27086
rect 54574 27010 54626 27022
rect 54686 27074 54738 27086
rect 54686 27010 54738 27022
rect 55246 27074 55298 27086
rect 55246 27010 55298 27022
rect 55470 27074 55522 27086
rect 55470 27010 55522 27022
rect 55582 27074 55634 27086
rect 55582 27010 55634 27022
rect 55806 27074 55858 27086
rect 58046 27074 58098 27086
rect 56690 27022 56702 27074
rect 56754 27022 56766 27074
rect 57474 27022 57486 27074
rect 57538 27022 57550 27074
rect 55806 27010 55858 27022
rect 58046 27010 58098 27022
rect 58830 27074 58882 27086
rect 61394 27022 61406 27074
rect 61458 27022 61470 27074
rect 58830 27010 58882 27022
rect 6750 26962 6802 26974
rect 2146 26910 2158 26962
rect 2210 26910 2222 26962
rect 4722 26910 4734 26962
rect 4786 26910 4798 26962
rect 6750 26898 6802 26910
rect 7310 26962 7362 26974
rect 7310 26898 7362 26910
rect 8206 26962 8258 26974
rect 15486 26962 15538 26974
rect 11890 26910 11902 26962
rect 11954 26910 11966 26962
rect 12450 26910 12462 26962
rect 12514 26910 12526 26962
rect 14018 26910 14030 26962
rect 14082 26910 14094 26962
rect 8206 26898 8258 26910
rect 15486 26898 15538 26910
rect 18734 26962 18786 26974
rect 21646 26962 21698 26974
rect 19282 26910 19294 26962
rect 19346 26910 19358 26962
rect 19618 26910 19630 26962
rect 19682 26910 19694 26962
rect 20738 26910 20750 26962
rect 20802 26910 20814 26962
rect 18734 26898 18786 26910
rect 21646 26898 21698 26910
rect 21982 26962 22034 26974
rect 24670 26962 24722 26974
rect 29150 26962 29202 26974
rect 23314 26910 23326 26962
rect 23378 26910 23390 26962
rect 24322 26910 24334 26962
rect 24386 26910 24398 26962
rect 25666 26910 25678 26962
rect 25730 26910 25742 26962
rect 27906 26910 27918 26962
rect 27970 26910 27982 26962
rect 28466 26910 28478 26962
rect 28530 26910 28542 26962
rect 21982 26898 22034 26910
rect 24670 26898 24722 26910
rect 29150 26898 29202 26910
rect 29262 26962 29314 26974
rect 29262 26898 29314 26910
rect 30494 26962 30546 26974
rect 33966 26962 34018 26974
rect 31490 26910 31502 26962
rect 31554 26910 31566 26962
rect 30494 26898 30546 26910
rect 33966 26898 34018 26910
rect 34526 26962 34578 26974
rect 34526 26898 34578 26910
rect 35198 26962 35250 26974
rect 41022 26962 41074 26974
rect 43598 26962 43650 26974
rect 37538 26910 37550 26962
rect 37602 26910 37614 26962
rect 40226 26910 40238 26962
rect 40290 26910 40302 26962
rect 43474 26910 43486 26962
rect 43538 26910 43550 26962
rect 44830 26962 44882 26974
rect 35198 26898 35250 26910
rect 41022 26898 41074 26910
rect 43598 26898 43650 26910
rect 43710 26906 43762 26918
rect 6862 26850 6914 26862
rect 8878 26850 8930 26862
rect 27358 26850 27410 26862
rect 8530 26798 8542 26850
rect 8594 26798 8606 26850
rect 10546 26798 10558 26850
rect 10610 26798 10622 26850
rect 6862 26786 6914 26798
rect 8878 26786 8930 26798
rect 27358 26786 27410 26798
rect 29486 26850 29538 26862
rect 44830 26898 44882 26910
rect 45054 26962 45106 26974
rect 49870 26962 49922 26974
rect 48738 26910 48750 26962
rect 48802 26910 48814 26962
rect 45054 26898 45106 26910
rect 49870 26898 49922 26910
rect 51550 26962 51602 26974
rect 51550 26898 51602 26910
rect 52670 26962 52722 26974
rect 56578 26910 56590 26962
rect 56642 26910 56654 26962
rect 59826 26910 59838 26962
rect 59890 26910 59902 26962
rect 52670 26898 52722 26910
rect 35522 26798 35534 26850
rect 35586 26798 35598 26850
rect 43710 26842 43762 26854
rect 43934 26850 43986 26862
rect 29486 26786 29538 26798
rect 43934 26786 43986 26798
rect 52782 26850 52834 26862
rect 52782 26786 52834 26798
rect 54350 26850 54402 26862
rect 54350 26786 54402 26798
rect 54798 26850 54850 26862
rect 61170 26798 61182 26850
rect 61234 26798 61246 26850
rect 54798 26786 54850 26798
rect 1344 26682 62608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 62608 26682
rect 1344 26596 62608 26630
rect 2046 26514 2098 26526
rect 2046 26450 2098 26462
rect 11790 26514 11842 26526
rect 13134 26514 13186 26526
rect 12226 26462 12238 26514
rect 12290 26462 12302 26514
rect 11790 26450 11842 26462
rect 13134 26450 13186 26462
rect 14590 26514 14642 26526
rect 14590 26450 14642 26462
rect 14926 26514 14978 26526
rect 14926 26450 14978 26462
rect 15038 26514 15090 26526
rect 19630 26514 19682 26526
rect 16818 26462 16830 26514
rect 16882 26462 16894 26514
rect 15038 26450 15090 26462
rect 19630 26450 19682 26462
rect 26238 26514 26290 26526
rect 26238 26450 26290 26462
rect 26350 26514 26402 26526
rect 26350 26450 26402 26462
rect 26798 26514 26850 26526
rect 33182 26514 33234 26526
rect 31714 26462 31726 26514
rect 31778 26462 31790 26514
rect 26798 26450 26850 26462
rect 33182 26450 33234 26462
rect 39902 26514 39954 26526
rect 39902 26450 39954 26462
rect 40126 26514 40178 26526
rect 40126 26450 40178 26462
rect 42926 26514 42978 26526
rect 49758 26514 49810 26526
rect 48738 26462 48750 26514
rect 48802 26462 48814 26514
rect 42926 26450 42978 26462
rect 49758 26450 49810 26462
rect 57710 26514 57762 26526
rect 57710 26450 57762 26462
rect 61630 26514 61682 26526
rect 61630 26450 61682 26462
rect 61742 26514 61794 26526
rect 61742 26450 61794 26462
rect 61966 26514 62018 26526
rect 61966 26450 62018 26462
rect 1710 26402 1762 26414
rect 22318 26402 22370 26414
rect 26126 26402 26178 26414
rect 33070 26402 33122 26414
rect 50094 26402 50146 26414
rect 62190 26402 62242 26414
rect 2930 26350 2942 26402
rect 2994 26350 3006 26402
rect 5170 26350 5182 26402
rect 5234 26350 5246 26402
rect 5618 26350 5630 26402
rect 5682 26350 5694 26402
rect 9986 26350 9998 26402
rect 10050 26350 10062 26402
rect 17938 26350 17950 26402
rect 18002 26350 18014 26402
rect 21298 26350 21310 26402
rect 21362 26350 21374 26402
rect 23314 26350 23326 26402
rect 23378 26350 23390 26402
rect 25778 26350 25790 26402
rect 25842 26350 25854 26402
rect 28018 26350 28030 26402
rect 28082 26350 28094 26402
rect 36306 26350 36318 26402
rect 36370 26350 36382 26402
rect 41122 26350 41134 26402
rect 41186 26350 41198 26402
rect 44706 26350 44718 26402
rect 44770 26350 44782 26402
rect 46162 26350 46174 26402
rect 46226 26350 46238 26402
rect 46610 26350 46622 26402
rect 46674 26350 46686 26402
rect 51650 26350 51662 26402
rect 51714 26350 51726 26402
rect 55794 26350 55806 26402
rect 55858 26350 55870 26402
rect 58594 26350 58606 26402
rect 58658 26350 58670 26402
rect 1710 26338 1762 26350
rect 22318 26338 22370 26350
rect 26126 26338 26178 26350
rect 33070 26338 33122 26350
rect 50094 26338 50146 26350
rect 62190 26338 62242 26350
rect 6750 26290 6802 26302
rect 6750 26226 6802 26238
rect 6862 26290 6914 26302
rect 7982 26290 8034 26302
rect 7298 26238 7310 26290
rect 7362 26238 7374 26290
rect 7746 26238 7758 26290
rect 7810 26238 7822 26290
rect 6862 26226 6914 26238
rect 7982 26226 8034 26238
rect 8206 26290 8258 26302
rect 8206 26226 8258 26238
rect 8542 26290 8594 26302
rect 8542 26226 8594 26238
rect 8766 26290 8818 26302
rect 8766 26226 8818 26238
rect 12574 26290 12626 26302
rect 13918 26290 13970 26302
rect 13122 26238 13134 26290
rect 13186 26238 13198 26290
rect 13682 26238 13694 26290
rect 13746 26238 13758 26290
rect 12574 26226 12626 26238
rect 13918 26226 13970 26238
rect 14814 26290 14866 26302
rect 16270 26290 16322 26302
rect 15810 26238 15822 26290
rect 15874 26238 15886 26290
rect 14814 26226 14866 26238
rect 16270 26226 16322 26238
rect 22206 26290 22258 26302
rect 22206 26226 22258 26238
rect 22542 26290 22594 26302
rect 31166 26290 31218 26302
rect 34526 26290 34578 26302
rect 47294 26290 47346 26302
rect 25890 26238 25902 26290
rect 25954 26238 25966 26290
rect 27906 26238 27918 26290
rect 27970 26238 27982 26290
rect 29026 26238 29038 26290
rect 29090 26238 29102 26290
rect 30482 26238 30494 26290
rect 30546 26238 30558 26290
rect 32162 26238 32174 26290
rect 32226 26238 32238 26290
rect 38098 26238 38110 26290
rect 38162 26238 38174 26290
rect 39442 26238 39454 26290
rect 39506 26238 39518 26290
rect 39666 26238 39678 26290
rect 39730 26238 39742 26290
rect 41010 26238 41022 26290
rect 41074 26238 41086 26290
rect 42242 26238 42254 26290
rect 42306 26238 42318 26290
rect 42466 26238 42478 26290
rect 42530 26238 42542 26290
rect 22542 26226 22594 26238
rect 31166 26226 31218 26238
rect 34526 26226 34578 26238
rect 47294 26226 47346 26238
rect 47518 26290 47570 26302
rect 47518 26226 47570 26238
rect 47742 26290 47794 26302
rect 49646 26290 49698 26302
rect 48962 26238 48974 26290
rect 49026 26238 49038 26290
rect 47742 26226 47794 26238
rect 49646 26226 49698 26238
rect 49870 26290 49922 26302
rect 59726 26290 59778 26302
rect 50978 26238 50990 26290
rect 51042 26238 51054 26290
rect 54450 26238 54462 26290
rect 54514 26238 54526 26290
rect 54786 26238 54798 26290
rect 54850 26238 54862 26290
rect 56018 26238 56030 26290
rect 56082 26238 56094 26290
rect 57026 26238 57038 26290
rect 57090 26238 57102 26290
rect 59042 26238 59054 26290
rect 59106 26238 59118 26290
rect 60162 26238 60174 26290
rect 60226 26238 60238 26290
rect 49870 26226 49922 26238
rect 59726 26226 59778 26238
rect 5854 26178 5906 26190
rect 5854 26114 5906 26126
rect 7870 26178 7922 26190
rect 7870 26114 7922 26126
rect 8430 26178 8482 26190
rect 8430 26114 8482 26126
rect 12798 26178 12850 26190
rect 12798 26114 12850 26126
rect 15374 26178 15426 26190
rect 15374 26114 15426 26126
rect 31390 26178 31442 26190
rect 33630 26178 33682 26190
rect 32386 26126 32398 26178
rect 32450 26126 32462 26178
rect 31390 26114 31442 26126
rect 33630 26114 33682 26126
rect 34190 26178 34242 26190
rect 34190 26114 34242 26126
rect 34750 26178 34802 26190
rect 40014 26178 40066 26190
rect 38546 26126 38558 26178
rect 38610 26126 38622 26178
rect 34750 26114 34802 26126
rect 40014 26114 40066 26126
rect 41694 26178 41746 26190
rect 41694 26114 41746 26126
rect 47630 26178 47682 26190
rect 55358 26178 55410 26190
rect 53778 26126 53790 26178
rect 53842 26126 53854 26178
rect 56690 26126 56702 26178
rect 56754 26126 56766 26178
rect 47630 26114 47682 26126
rect 55358 26114 55410 26126
rect 4734 26066 4786 26078
rect 4734 26002 4786 26014
rect 6190 26066 6242 26078
rect 16494 26066 16546 26078
rect 7410 26014 7422 26066
rect 7474 26014 7486 26066
rect 13346 26014 13358 26066
rect 13410 26014 13422 26066
rect 6190 26002 6242 26014
rect 16494 26002 16546 26014
rect 20078 26066 20130 26078
rect 20078 26002 20130 26014
rect 24558 26066 24610 26078
rect 37438 26066 37490 26078
rect 29138 26014 29150 26066
rect 29202 26014 29214 26066
rect 35074 26014 35086 26066
rect 35138 26014 35150 26066
rect 24558 26002 24610 26014
rect 37438 26002 37490 26014
rect 45502 26066 45554 26078
rect 45502 26002 45554 26014
rect 45838 26066 45890 26078
rect 45838 26002 45890 26014
rect 47070 26066 47122 26078
rect 60386 26014 60398 26066
rect 60450 26014 60462 26066
rect 47070 26002 47122 26014
rect 1344 25898 62608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 62608 25898
rect 1344 25812 62608 25846
rect 16494 25730 16546 25742
rect 16494 25666 16546 25678
rect 20302 25730 20354 25742
rect 24222 25730 24274 25742
rect 22754 25678 22766 25730
rect 22818 25678 22830 25730
rect 20302 25666 20354 25678
rect 24222 25666 24274 25678
rect 26462 25730 26514 25742
rect 31390 25730 31442 25742
rect 44830 25730 44882 25742
rect 27570 25678 27582 25730
rect 27634 25678 27646 25730
rect 34402 25678 34414 25730
rect 34466 25727 34478 25730
rect 34738 25727 34750 25730
rect 34466 25681 34750 25727
rect 34466 25678 34478 25681
rect 34738 25678 34750 25681
rect 34802 25678 34814 25730
rect 26462 25666 26514 25678
rect 31390 25666 31442 25678
rect 44830 25666 44882 25678
rect 45390 25730 45442 25742
rect 45390 25666 45442 25678
rect 45614 25730 45666 25742
rect 45614 25666 45666 25678
rect 46062 25730 46114 25742
rect 54562 25678 54574 25730
rect 54626 25678 54638 25730
rect 58594 25678 58606 25730
rect 58658 25678 58670 25730
rect 46062 25666 46114 25678
rect 10334 25618 10386 25630
rect 9650 25566 9662 25618
rect 9714 25566 9726 25618
rect 10334 25554 10386 25566
rect 10670 25618 10722 25630
rect 28702 25618 28754 25630
rect 17938 25566 17950 25618
rect 18002 25566 18014 25618
rect 25666 25566 25678 25618
rect 25730 25566 25742 25618
rect 10670 25554 10722 25566
rect 28702 25554 28754 25566
rect 34862 25618 34914 25630
rect 54238 25618 54290 25630
rect 39106 25566 39118 25618
rect 39170 25566 39182 25618
rect 45154 25566 45166 25618
rect 45218 25566 45230 25618
rect 46610 25566 46622 25618
rect 46674 25566 46686 25618
rect 48738 25566 48750 25618
rect 48802 25566 48814 25618
rect 34862 25554 34914 25566
rect 54238 25554 54290 25566
rect 55134 25618 55186 25630
rect 60958 25618 61010 25630
rect 58706 25566 58718 25618
rect 58770 25566 58782 25618
rect 55134 25554 55186 25566
rect 60958 25554 61010 25566
rect 5742 25506 5794 25518
rect 12014 25506 12066 25518
rect 4946 25454 4958 25506
rect 5010 25454 5022 25506
rect 6402 25454 6414 25506
rect 6466 25454 6478 25506
rect 6738 25454 6750 25506
rect 6802 25454 6814 25506
rect 5742 25442 5794 25454
rect 12014 25442 12066 25454
rect 12686 25506 12738 25518
rect 12686 25442 12738 25454
rect 13470 25506 13522 25518
rect 13470 25442 13522 25454
rect 17054 25506 17106 25518
rect 18510 25506 18562 25518
rect 17602 25454 17614 25506
rect 17666 25454 17678 25506
rect 17054 25442 17106 25454
rect 18510 25442 18562 25454
rect 18846 25506 18898 25518
rect 21870 25506 21922 25518
rect 26238 25506 26290 25518
rect 19618 25454 19630 25506
rect 19682 25454 19694 25506
rect 22418 25454 22430 25506
rect 22482 25454 22494 25506
rect 23538 25454 23550 25506
rect 23602 25454 23614 25506
rect 24770 25454 24782 25506
rect 24834 25454 24846 25506
rect 25218 25454 25230 25506
rect 25282 25454 25294 25506
rect 26002 25454 26014 25506
rect 26066 25454 26078 25506
rect 18846 25442 18898 25454
rect 21870 25442 21922 25454
rect 26238 25442 26290 25454
rect 27022 25506 27074 25518
rect 35422 25506 35474 25518
rect 32386 25454 32398 25506
rect 32450 25454 32462 25506
rect 33058 25454 33070 25506
rect 33122 25454 33134 25506
rect 34178 25454 34190 25506
rect 34242 25454 34254 25506
rect 27022 25442 27074 25454
rect 35422 25442 35474 25454
rect 36990 25506 37042 25518
rect 36990 25442 37042 25454
rect 37662 25506 37714 25518
rect 39566 25506 39618 25518
rect 38546 25454 38558 25506
rect 38610 25454 38622 25506
rect 37662 25442 37714 25454
rect 39566 25442 39618 25454
rect 41358 25506 41410 25518
rect 41358 25442 41410 25454
rect 41694 25506 41746 25518
rect 41694 25442 41746 25454
rect 42590 25506 42642 25518
rect 42590 25442 42642 25454
rect 42926 25506 42978 25518
rect 42926 25442 42978 25454
rect 44270 25506 44322 25518
rect 44270 25442 44322 25454
rect 45054 25506 45106 25518
rect 52782 25506 52834 25518
rect 49410 25454 49422 25506
rect 49474 25454 49486 25506
rect 50866 25454 50878 25506
rect 50930 25454 50942 25506
rect 45054 25442 45106 25454
rect 52782 25442 52834 25454
rect 54014 25506 54066 25518
rect 54014 25442 54066 25454
rect 54910 25506 54962 25518
rect 54910 25442 54962 25454
rect 55806 25506 55858 25518
rect 55806 25442 55858 25454
rect 56030 25506 56082 25518
rect 57138 25454 57150 25506
rect 57202 25454 57214 25506
rect 58594 25454 58606 25506
rect 58658 25454 58670 25506
rect 56030 25442 56082 25454
rect 4286 25394 4338 25406
rect 2370 25342 2382 25394
rect 2434 25342 2446 25394
rect 4286 25330 4338 25342
rect 4398 25394 4450 25406
rect 4398 25330 4450 25342
rect 5966 25394 6018 25406
rect 10782 25394 10834 25406
rect 7522 25342 7534 25394
rect 7586 25342 7598 25394
rect 5966 25330 6018 25342
rect 10782 25330 10834 25342
rect 11230 25394 11282 25406
rect 11230 25330 11282 25342
rect 11342 25394 11394 25406
rect 11342 25330 11394 25342
rect 11678 25394 11730 25406
rect 11678 25330 11730 25342
rect 12350 25394 12402 25406
rect 12350 25330 12402 25342
rect 12910 25394 12962 25406
rect 18286 25394 18338 25406
rect 22206 25394 22258 25406
rect 14690 25342 14702 25394
rect 14754 25342 14766 25394
rect 19506 25342 19518 25394
rect 19570 25342 19582 25394
rect 21522 25342 21534 25394
rect 21586 25342 21598 25394
rect 12910 25330 12962 25342
rect 18286 25330 18338 25342
rect 22206 25330 22258 25342
rect 23886 25394 23938 25406
rect 23886 25330 23938 25342
rect 24334 25394 24386 25406
rect 24334 25330 24386 25342
rect 28142 25394 28194 25406
rect 36094 25394 36146 25406
rect 33506 25342 33518 25394
rect 33570 25342 33582 25394
rect 35074 25342 35086 25394
rect 35138 25342 35150 25394
rect 28142 25330 28194 25342
rect 36094 25330 36146 25342
rect 37326 25394 37378 25406
rect 37326 25330 37378 25342
rect 38222 25394 38274 25406
rect 46174 25394 46226 25406
rect 43138 25342 43150 25394
rect 43202 25342 43214 25394
rect 43474 25342 43486 25394
rect 43538 25342 43550 25394
rect 38222 25330 38274 25342
rect 46174 25330 46226 25342
rect 50318 25394 50370 25406
rect 50318 25330 50370 25342
rect 50542 25394 50594 25406
rect 50542 25330 50594 25342
rect 50654 25394 50706 25406
rect 50654 25330 50706 25342
rect 51102 25394 51154 25406
rect 51102 25330 51154 25342
rect 52894 25394 52946 25406
rect 60622 25394 60674 25406
rect 57250 25342 57262 25394
rect 57314 25342 57326 25394
rect 61282 25342 61294 25394
rect 61346 25342 61358 25394
rect 61506 25342 61518 25394
rect 61570 25342 61582 25394
rect 52894 25330 52946 25342
rect 60622 25330 60674 25342
rect 3726 25282 3778 25294
rect 3726 25218 3778 25230
rect 4062 25282 4114 25294
rect 4062 25218 4114 25230
rect 4734 25282 4786 25294
rect 4734 25218 4786 25230
rect 5630 25282 5682 25294
rect 5630 25218 5682 25230
rect 5854 25282 5906 25294
rect 5854 25218 5906 25230
rect 11006 25282 11058 25294
rect 11006 25218 11058 25230
rect 12462 25282 12514 25294
rect 17166 25282 17218 25294
rect 13794 25230 13806 25282
rect 13858 25230 13870 25282
rect 12462 25218 12514 25230
rect 17166 25218 17218 25230
rect 17390 25282 17442 25294
rect 17390 25218 17442 25230
rect 18510 25282 18562 25294
rect 18510 25218 18562 25230
rect 20638 25282 20690 25294
rect 35758 25282 35810 25294
rect 30034 25230 30046 25282
rect 30098 25230 30110 25282
rect 20638 25218 20690 25230
rect 35758 25218 35810 25230
rect 49758 25282 49810 25294
rect 49758 25218 49810 25230
rect 49870 25282 49922 25294
rect 49870 25218 49922 25230
rect 50094 25282 50146 25294
rect 51774 25282 51826 25294
rect 51426 25230 51438 25282
rect 51490 25230 51502 25282
rect 50094 25218 50146 25230
rect 51774 25218 51826 25230
rect 53006 25282 53058 25294
rect 53006 25218 53058 25230
rect 53230 25282 53282 25294
rect 53666 25230 53678 25282
rect 53730 25230 53742 25282
rect 55458 25230 55470 25282
rect 55522 25230 55534 25282
rect 53230 25218 53282 25230
rect 1344 25114 62608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 62608 25114
rect 1344 25028 62608 25062
rect 6414 24946 6466 24958
rect 6414 24882 6466 24894
rect 7534 24946 7586 24958
rect 7534 24882 7586 24894
rect 8990 24946 9042 24958
rect 8990 24882 9042 24894
rect 15038 24946 15090 24958
rect 16606 24946 16658 24958
rect 30382 24946 30434 24958
rect 16146 24894 16158 24946
rect 16210 24894 16222 24946
rect 24658 24894 24670 24946
rect 24722 24894 24734 24946
rect 15038 24882 15090 24894
rect 16606 24882 16658 24894
rect 30382 24882 30434 24894
rect 30494 24946 30546 24958
rect 30494 24882 30546 24894
rect 30606 24946 30658 24958
rect 30606 24882 30658 24894
rect 37550 24946 37602 24958
rect 37550 24882 37602 24894
rect 38334 24946 38386 24958
rect 38334 24882 38386 24894
rect 41022 24946 41074 24958
rect 41022 24882 41074 24894
rect 43150 24946 43202 24958
rect 43150 24882 43202 24894
rect 49310 24946 49362 24958
rect 49310 24882 49362 24894
rect 56814 24946 56866 24958
rect 56814 24882 56866 24894
rect 57038 24946 57090 24958
rect 57038 24882 57090 24894
rect 58830 24946 58882 24958
rect 58830 24882 58882 24894
rect 8430 24834 8482 24846
rect 5618 24782 5630 24834
rect 5682 24782 5694 24834
rect 6962 24782 6974 24834
rect 7026 24782 7038 24834
rect 8430 24770 8482 24782
rect 13134 24834 13186 24846
rect 17838 24834 17890 24846
rect 14018 24782 14030 24834
rect 14082 24782 14094 24834
rect 13134 24770 13186 24782
rect 17838 24770 17890 24782
rect 18062 24834 18114 24846
rect 22766 24834 22818 24846
rect 31950 24834 32002 24846
rect 19618 24782 19630 24834
rect 19682 24782 19694 24834
rect 21298 24782 21310 24834
rect 21362 24782 21374 24834
rect 25890 24782 25902 24834
rect 25954 24782 25966 24834
rect 29138 24782 29150 24834
rect 29202 24782 29214 24834
rect 18062 24770 18114 24782
rect 22766 24770 22818 24782
rect 31950 24770 32002 24782
rect 32062 24834 32114 24846
rect 38110 24834 38162 24846
rect 33394 24782 33406 24834
rect 33458 24782 33470 24834
rect 36306 24782 36318 24834
rect 36370 24782 36382 24834
rect 32062 24770 32114 24782
rect 38110 24770 38162 24782
rect 38894 24834 38946 24846
rect 48078 24834 48130 24846
rect 57150 24834 57202 24846
rect 40226 24782 40238 24834
rect 40290 24782 40302 24834
rect 41906 24782 41918 24834
rect 41970 24782 41982 24834
rect 47058 24782 47070 24834
rect 47122 24782 47134 24834
rect 47282 24782 47294 24834
rect 47346 24782 47358 24834
rect 51314 24782 51326 24834
rect 51378 24782 51390 24834
rect 51874 24782 51886 24834
rect 51938 24782 51950 24834
rect 55234 24782 55246 24834
rect 55298 24782 55310 24834
rect 57810 24782 57822 24834
rect 57874 24782 57886 24834
rect 58258 24782 58270 24834
rect 58322 24782 58334 24834
rect 60050 24782 60062 24834
rect 60114 24782 60126 24834
rect 38894 24770 38946 24782
rect 48078 24770 48130 24782
rect 57150 24770 57202 24782
rect 5070 24722 5122 24734
rect 7198 24722 7250 24734
rect 3826 24670 3838 24722
rect 3890 24670 3902 24722
rect 5842 24670 5854 24722
rect 5906 24670 5918 24722
rect 6626 24670 6638 24722
rect 6690 24670 6702 24722
rect 5070 24658 5122 24670
rect 7198 24658 7250 24670
rect 7870 24722 7922 24734
rect 7870 24658 7922 24670
rect 8206 24722 8258 24734
rect 13022 24722 13074 24734
rect 9538 24670 9550 24722
rect 9602 24670 9614 24722
rect 8206 24658 8258 24670
rect 13022 24658 13074 24670
rect 13358 24722 13410 24734
rect 13358 24658 13410 24670
rect 13470 24722 13522 24734
rect 15822 24722 15874 24734
rect 17502 24722 17554 24734
rect 18846 24722 18898 24734
rect 13906 24670 13918 24722
rect 13970 24670 13982 24722
rect 16818 24670 16830 24722
rect 16882 24670 16894 24722
rect 18386 24670 18398 24722
rect 18450 24670 18462 24722
rect 13470 24658 13522 24670
rect 15822 24658 15874 24670
rect 17502 24658 17554 24670
rect 18846 24658 18898 24670
rect 19182 24722 19234 24734
rect 19182 24658 19234 24670
rect 19966 24722 20018 24734
rect 22206 24722 22258 24734
rect 21410 24670 21422 24722
rect 21474 24670 21486 24722
rect 19966 24658 20018 24670
rect 22206 24658 22258 24670
rect 23662 24722 23714 24734
rect 32174 24722 32226 24734
rect 24434 24670 24446 24722
rect 24498 24670 24510 24722
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 25778 24670 25790 24722
rect 25842 24670 25854 24722
rect 26786 24670 26798 24722
rect 26850 24670 26862 24722
rect 27906 24670 27918 24722
rect 27970 24670 27982 24722
rect 29810 24670 29822 24722
rect 29874 24670 29886 24722
rect 30930 24670 30942 24722
rect 30994 24670 31006 24722
rect 31378 24670 31390 24722
rect 31442 24670 31454 24722
rect 31714 24670 31726 24722
rect 31778 24670 31790 24722
rect 23662 24658 23714 24670
rect 32174 24658 32226 24670
rect 37998 24722 38050 24734
rect 46398 24722 46450 24734
rect 38658 24670 38670 24722
rect 38722 24670 38734 24722
rect 39330 24670 39342 24722
rect 39394 24670 39406 24722
rect 44482 24670 44494 24722
rect 44546 24670 44558 24722
rect 45042 24670 45054 24722
rect 45106 24670 45118 24722
rect 45490 24670 45502 24722
rect 45554 24670 45566 24722
rect 37998 24658 38050 24670
rect 46398 24658 46450 24670
rect 47966 24722 48018 24734
rect 47966 24658 48018 24670
rect 48302 24722 48354 24734
rect 48302 24658 48354 24670
rect 49534 24722 49586 24734
rect 49534 24658 49586 24670
rect 49758 24722 49810 24734
rect 57262 24722 57314 24734
rect 50978 24670 50990 24722
rect 51042 24670 51054 24722
rect 51986 24670 51998 24722
rect 52050 24670 52062 24722
rect 52994 24670 53006 24722
rect 53058 24670 53070 24722
rect 53330 24670 53342 24722
rect 53394 24670 53406 24722
rect 54674 24670 54686 24722
rect 54738 24670 54750 24722
rect 55122 24670 55134 24722
rect 55186 24670 55198 24722
rect 55458 24670 55470 24722
rect 55522 24670 55534 24722
rect 49758 24658 49810 24670
rect 57262 24658 57314 24670
rect 58494 24722 58546 24734
rect 59266 24670 59278 24722
rect 59330 24670 59342 24722
rect 58494 24658 58546 24670
rect 15598 24610 15650 24622
rect 10322 24558 10334 24610
rect 10386 24558 10398 24610
rect 12450 24558 12462 24610
rect 12514 24558 12526 24610
rect 15598 24546 15650 24558
rect 17614 24610 17666 24622
rect 17614 24546 17666 24558
rect 19070 24610 19122 24622
rect 48862 24610 48914 24622
rect 25666 24558 25678 24610
rect 25730 24558 25742 24610
rect 30930 24558 30942 24610
rect 30994 24607 31006 24610
rect 31154 24607 31166 24610
rect 30994 24561 31166 24607
rect 30994 24558 31006 24561
rect 31154 24558 31166 24561
rect 31218 24558 31230 24610
rect 44706 24558 44718 24610
rect 44770 24558 44782 24610
rect 19070 24546 19122 24558
rect 48862 24546 48914 24558
rect 49646 24610 49698 24622
rect 49646 24546 49698 24558
rect 52446 24610 52498 24622
rect 62178 24558 62190 24610
rect 62242 24558 62254 24610
rect 52446 24546 52498 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 4734 24498 4786 24510
rect 4734 24434 4786 24446
rect 6750 24498 6802 24510
rect 6750 24434 6802 24446
rect 7646 24498 7698 24510
rect 7646 24434 7698 24446
rect 14702 24498 14754 24510
rect 14702 24434 14754 24446
rect 16494 24498 16546 24510
rect 16494 24434 16546 24446
rect 18734 24498 18786 24510
rect 18734 24434 18786 24446
rect 20414 24498 20466 24510
rect 20414 24434 20466 24446
rect 20750 24498 20802 24510
rect 23438 24498 23490 24510
rect 35310 24498 35362 24510
rect 46734 24498 46786 24510
rect 23090 24446 23102 24498
rect 23154 24446 23166 24498
rect 27122 24446 27134 24498
rect 27186 24446 27198 24498
rect 40114 24446 40126 24498
rect 40178 24446 40190 24498
rect 20750 24434 20802 24446
rect 23438 24434 23490 24446
rect 35310 24434 35362 24446
rect 46734 24434 46786 24446
rect 50206 24498 50258 24510
rect 50206 24434 50258 24446
rect 50542 24498 50594 24510
rect 50542 24434 50594 24446
rect 1344 24330 62608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 62608 24330
rect 1344 24244 62608 24278
rect 3502 24162 3554 24174
rect 3502 24098 3554 24110
rect 6526 24162 6578 24174
rect 6526 24098 6578 24110
rect 8094 24162 8146 24174
rect 8094 24098 8146 24110
rect 11790 24162 11842 24174
rect 11790 24098 11842 24110
rect 12238 24162 12290 24174
rect 12238 24098 12290 24110
rect 12462 24162 12514 24174
rect 15374 24162 15426 24174
rect 13682 24110 13694 24162
rect 13746 24110 13758 24162
rect 12462 24098 12514 24110
rect 15374 24098 15426 24110
rect 18062 24162 18114 24174
rect 18062 24098 18114 24110
rect 26014 24162 26066 24174
rect 26014 24098 26066 24110
rect 26350 24162 26402 24174
rect 33182 24162 33234 24174
rect 27570 24110 27582 24162
rect 27634 24110 27646 24162
rect 26350 24098 26402 24110
rect 33182 24098 33234 24110
rect 35198 24162 35250 24174
rect 44382 24162 44434 24174
rect 60062 24162 60114 24174
rect 39218 24110 39230 24162
rect 39282 24110 39294 24162
rect 53554 24110 53566 24162
rect 53618 24110 53630 24162
rect 35198 24098 35250 24110
rect 44382 24098 44434 24110
rect 60062 24098 60114 24110
rect 5070 24050 5122 24062
rect 5070 23986 5122 23998
rect 5854 24050 5906 24062
rect 5854 23986 5906 23998
rect 6974 24050 7026 24062
rect 6974 23986 7026 23998
rect 10894 24050 10946 24062
rect 10894 23986 10946 23998
rect 24334 24050 24386 24062
rect 24334 23986 24386 23998
rect 29262 24050 29314 24062
rect 44942 24050 44994 24062
rect 40114 23998 40126 24050
rect 40178 23998 40190 24050
rect 47842 23998 47854 24050
rect 47906 23998 47918 24050
rect 54898 23998 54910 24050
rect 54962 23998 54974 24050
rect 57138 23998 57150 24050
rect 57202 23998 57214 24050
rect 29262 23986 29314 23998
rect 44942 23986 44994 23998
rect 4062 23938 4114 23950
rect 4062 23874 4114 23886
rect 4286 23938 4338 23950
rect 4286 23874 4338 23886
rect 6750 23938 6802 23950
rect 6750 23874 6802 23886
rect 7086 23938 7138 23950
rect 7086 23874 7138 23886
rect 7310 23938 7362 23950
rect 7310 23874 7362 23886
rect 11902 23938 11954 23950
rect 14254 23938 14306 23950
rect 18398 23938 18450 23950
rect 19630 23938 19682 23950
rect 13570 23886 13582 23938
rect 13634 23886 13646 23938
rect 15026 23886 15038 23938
rect 15090 23886 15102 23938
rect 19170 23886 19182 23938
rect 19234 23886 19246 23938
rect 11902 23874 11954 23886
rect 14254 23874 14306 23886
rect 18398 23874 18450 23886
rect 19630 23874 19682 23886
rect 19966 23938 20018 23950
rect 19966 23874 20018 23886
rect 20078 23938 20130 23950
rect 24446 23938 24498 23950
rect 26126 23938 26178 23950
rect 28366 23938 28418 23950
rect 31614 23938 31666 23950
rect 20178 23886 20190 23938
rect 20242 23886 20254 23938
rect 24098 23886 24110 23938
rect 24162 23886 24174 23938
rect 24658 23886 24670 23938
rect 24722 23886 24734 23938
rect 25666 23886 25678 23938
rect 25730 23886 25742 23938
rect 27010 23886 27022 23938
rect 27074 23886 27086 23938
rect 29810 23886 29822 23938
rect 29874 23886 29886 23938
rect 20078 23874 20130 23886
rect 24446 23874 24498 23886
rect 26126 23874 26178 23886
rect 28366 23874 28418 23886
rect 31614 23874 31666 23886
rect 32062 23938 32114 23950
rect 33518 23938 33570 23950
rect 39342 23938 39394 23950
rect 41582 23938 41634 23950
rect 51102 23938 51154 23950
rect 32162 23886 32174 23938
rect 32226 23886 32238 23938
rect 34178 23886 34190 23938
rect 34242 23886 34254 23938
rect 38994 23886 39006 23938
rect 39058 23886 39070 23938
rect 39778 23886 39790 23938
rect 39842 23886 39854 23938
rect 45938 23886 45950 23938
rect 46002 23886 46014 23938
rect 46722 23886 46734 23938
rect 46786 23886 46798 23938
rect 47506 23886 47518 23938
rect 47570 23886 47582 23938
rect 48626 23886 48638 23938
rect 48690 23886 48702 23938
rect 49410 23886 49422 23938
rect 49474 23886 49486 23938
rect 50642 23886 50654 23938
rect 50706 23886 50718 23938
rect 32062 23874 32114 23886
rect 33518 23874 33570 23886
rect 39342 23874 39394 23886
rect 41582 23874 41634 23886
rect 51102 23874 51154 23886
rect 51438 23938 51490 23950
rect 51438 23874 51490 23886
rect 51662 23938 51714 23950
rect 60958 23938 61010 23950
rect 52882 23886 52894 23938
rect 52946 23886 52958 23938
rect 54786 23886 54798 23938
rect 54850 23886 54862 23938
rect 57026 23886 57038 23938
rect 57090 23886 57102 23938
rect 51662 23874 51714 23886
rect 60958 23874 61010 23886
rect 6302 23826 6354 23838
rect 2370 23774 2382 23826
rect 2434 23774 2446 23826
rect 6302 23762 6354 23774
rect 7758 23826 7810 23838
rect 7758 23762 7810 23774
rect 7982 23826 8034 23838
rect 7982 23762 8034 23774
rect 9774 23826 9826 23838
rect 9774 23762 9826 23774
rect 11118 23826 11170 23838
rect 11118 23762 11170 23774
rect 11454 23826 11506 23838
rect 11454 23762 11506 23774
rect 11678 23826 11730 23838
rect 25454 23826 25506 23838
rect 14018 23774 14030 23826
rect 14082 23774 14094 23826
rect 17266 23774 17278 23826
rect 17330 23774 17342 23826
rect 18946 23774 18958 23826
rect 19010 23774 19022 23826
rect 21858 23774 21870 23826
rect 21922 23774 21934 23826
rect 24882 23774 24894 23826
rect 24946 23774 24958 23826
rect 11678 23762 11730 23774
rect 25454 23762 25506 23774
rect 25902 23826 25954 23838
rect 28478 23826 28530 23838
rect 27906 23774 27918 23826
rect 27970 23774 27982 23826
rect 25902 23762 25954 23774
rect 28478 23762 28530 23774
rect 29486 23826 29538 23838
rect 45278 23826 45330 23838
rect 49982 23826 50034 23838
rect 31826 23774 31838 23826
rect 31890 23774 31902 23826
rect 34290 23774 34302 23826
rect 34354 23774 34366 23826
rect 35410 23774 35422 23826
rect 35474 23774 35486 23826
rect 35746 23774 35758 23826
rect 35810 23774 35822 23826
rect 37314 23774 37326 23826
rect 37378 23774 37390 23826
rect 42578 23774 42590 23826
rect 42642 23774 42654 23826
rect 46834 23774 46846 23826
rect 46898 23774 46910 23826
rect 47618 23774 47630 23826
rect 47682 23774 47694 23826
rect 49298 23774 49310 23826
rect 49362 23774 49374 23826
rect 29486 23762 29538 23774
rect 45278 23762 45330 23774
rect 49982 23762 50034 23774
rect 50878 23826 50930 23838
rect 56590 23826 56642 23838
rect 53442 23774 53454 23826
rect 53506 23774 53518 23826
rect 50878 23762 50930 23774
rect 56590 23762 56642 23774
rect 56702 23826 56754 23838
rect 60622 23826 60674 23838
rect 58146 23774 58158 23826
rect 58210 23774 58222 23826
rect 61170 23774 61182 23826
rect 61234 23774 61246 23826
rect 61618 23774 61630 23826
rect 61682 23774 61694 23826
rect 56702 23762 56754 23774
rect 60622 23762 60674 23774
rect 6414 23714 6466 23726
rect 4610 23662 4622 23714
rect 4674 23662 4686 23714
rect 6414 23650 6466 23662
rect 8766 23714 8818 23726
rect 8766 23650 8818 23662
rect 9214 23714 9266 23726
rect 9214 23650 9266 23662
rect 9438 23714 9490 23726
rect 9438 23650 9490 23662
rect 9662 23714 9714 23726
rect 9662 23650 9714 23662
rect 10334 23714 10386 23726
rect 10334 23650 10386 23662
rect 11230 23714 11282 23726
rect 11230 23650 11282 23662
rect 14142 23714 14194 23726
rect 19742 23714 19794 23726
rect 14802 23662 14814 23714
rect 14866 23662 14878 23714
rect 14142 23650 14194 23662
rect 19742 23650 19794 23662
rect 23102 23714 23154 23726
rect 23102 23650 23154 23662
rect 28702 23714 28754 23726
rect 28702 23650 28754 23662
rect 29150 23714 29202 23726
rect 29150 23650 29202 23662
rect 29374 23714 29426 23726
rect 29374 23650 29426 23662
rect 30382 23714 30434 23726
rect 30382 23650 30434 23662
rect 30606 23714 30658 23726
rect 30606 23650 30658 23662
rect 30718 23714 30770 23726
rect 30718 23650 30770 23662
rect 30830 23714 30882 23726
rect 30830 23650 30882 23662
rect 31390 23714 31442 23726
rect 31390 23650 31442 23662
rect 32398 23714 32450 23726
rect 32398 23650 32450 23662
rect 34862 23714 34914 23726
rect 34862 23650 34914 23662
rect 36990 23714 37042 23726
rect 36990 23650 37042 23662
rect 41694 23714 41746 23726
rect 41694 23650 41746 23662
rect 41918 23714 41970 23726
rect 41918 23650 41970 23662
rect 44830 23714 44882 23726
rect 44830 23650 44882 23662
rect 45054 23714 45106 23726
rect 51326 23714 51378 23726
rect 45938 23662 45950 23714
rect 46002 23662 46014 23714
rect 45054 23650 45106 23662
rect 51326 23650 51378 23662
rect 56366 23714 56418 23726
rect 56366 23650 56418 23662
rect 1344 23546 62608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 62608 23546
rect 1344 23460 62608 23494
rect 2046 23378 2098 23390
rect 9774 23378 9826 23390
rect 6850 23326 6862 23378
rect 6914 23326 6926 23378
rect 2046 23314 2098 23326
rect 9774 23314 9826 23326
rect 17614 23378 17666 23390
rect 17614 23314 17666 23326
rect 18174 23378 18226 23390
rect 25230 23378 25282 23390
rect 19394 23326 19406 23378
rect 19458 23326 19470 23378
rect 18174 23314 18226 23326
rect 25230 23314 25282 23326
rect 29934 23378 29986 23390
rect 35422 23378 35474 23390
rect 34290 23326 34302 23378
rect 34354 23326 34366 23378
rect 29934 23314 29986 23326
rect 35422 23314 35474 23326
rect 36766 23378 36818 23390
rect 36766 23314 36818 23326
rect 37438 23378 37490 23390
rect 37438 23314 37490 23326
rect 40126 23378 40178 23390
rect 40126 23314 40178 23326
rect 40238 23378 40290 23390
rect 47518 23378 47570 23390
rect 46274 23326 46286 23378
rect 46338 23326 46350 23378
rect 56578 23326 56590 23378
rect 56642 23326 56654 23378
rect 40238 23314 40290 23326
rect 47518 23314 47570 23326
rect 1710 23266 1762 23278
rect 1710 23202 1762 23214
rect 2606 23266 2658 23278
rect 16046 23266 16098 23278
rect 11554 23214 11566 23266
rect 11618 23214 11630 23266
rect 14802 23214 14814 23266
rect 14866 23214 14878 23266
rect 15362 23214 15374 23266
rect 15426 23214 15438 23266
rect 2606 23202 2658 23214
rect 16046 23202 16098 23214
rect 16830 23266 16882 23278
rect 16830 23202 16882 23214
rect 17838 23266 17890 23278
rect 23438 23266 23490 23278
rect 20514 23214 20526 23266
rect 20578 23214 20590 23266
rect 17838 23202 17890 23214
rect 23438 23202 23490 23214
rect 23662 23266 23714 23278
rect 33182 23266 33234 23278
rect 36990 23266 37042 23278
rect 31714 23214 31726 23266
rect 31778 23214 31790 23266
rect 35858 23214 35870 23266
rect 35922 23214 35934 23266
rect 23662 23202 23714 23214
rect 33182 23202 33234 23214
rect 36990 23202 37042 23214
rect 37550 23266 37602 23278
rect 40014 23266 40066 23278
rect 39106 23214 39118 23266
rect 39170 23214 39182 23266
rect 37550 23202 37602 23214
rect 40014 23202 40066 23214
rect 44606 23266 44658 23278
rect 47182 23266 47234 23278
rect 46610 23214 46622 23266
rect 46674 23214 46686 23266
rect 44606 23202 44658 23214
rect 47182 23202 47234 23214
rect 47406 23266 47458 23278
rect 47406 23202 47458 23214
rect 49646 23266 49698 23278
rect 53554 23214 53566 23266
rect 53618 23214 53630 23266
rect 60946 23214 60958 23266
rect 61010 23214 61022 23266
rect 49646 23202 49698 23214
rect 2830 23154 2882 23166
rect 6190 23154 6242 23166
rect 7534 23154 7586 23166
rect 3490 23102 3502 23154
rect 3554 23102 3566 23154
rect 5954 23102 5966 23154
rect 6018 23102 6030 23154
rect 7074 23102 7086 23154
rect 7138 23102 7150 23154
rect 2830 23090 2882 23102
rect 6190 23090 6242 23102
rect 7534 23090 7586 23102
rect 8430 23154 8482 23166
rect 16158 23154 16210 23166
rect 18286 23154 18338 23166
rect 10098 23102 10110 23154
rect 10162 23102 10174 23154
rect 14354 23102 14366 23154
rect 14418 23102 14430 23154
rect 15138 23102 15150 23154
rect 15202 23102 15214 23154
rect 16594 23102 16606 23154
rect 16658 23102 16670 23154
rect 8430 23090 8482 23102
rect 16158 23090 16210 23102
rect 18286 23090 18338 23102
rect 18510 23154 18562 23166
rect 18510 23090 18562 23102
rect 18958 23154 19010 23166
rect 22990 23154 23042 23166
rect 19618 23102 19630 23154
rect 19682 23102 19694 23154
rect 21074 23102 21086 23154
rect 21138 23102 21150 23154
rect 22418 23102 22430 23154
rect 22482 23102 22494 23154
rect 18958 23090 19010 23102
rect 22990 23090 23042 23102
rect 23214 23154 23266 23166
rect 25790 23154 25842 23166
rect 27806 23154 27858 23166
rect 36654 23154 36706 23166
rect 24546 23102 24558 23154
rect 24610 23102 24622 23154
rect 27570 23102 27582 23154
rect 27634 23102 27646 23154
rect 28466 23102 28478 23154
rect 28530 23102 28542 23154
rect 29586 23102 29598 23154
rect 29650 23102 29662 23154
rect 36082 23102 36094 23154
rect 36146 23102 36158 23154
rect 23214 23090 23266 23102
rect 25790 23090 25842 23102
rect 27806 23090 27858 23102
rect 36654 23090 36706 23102
rect 38334 23154 38386 23166
rect 40350 23154 40402 23166
rect 42366 23154 42418 23166
rect 44942 23154 44994 23166
rect 47854 23154 47906 23166
rect 51550 23154 51602 23166
rect 56926 23154 56978 23166
rect 38994 23102 39006 23154
rect 39058 23102 39070 23154
rect 39554 23102 39566 23154
rect 39618 23102 39630 23154
rect 41794 23102 41806 23154
rect 41858 23102 41870 23154
rect 43026 23102 43038 23154
rect 43090 23102 43102 23154
rect 44258 23102 44270 23154
rect 44322 23102 44334 23154
rect 45714 23102 45726 23154
rect 45778 23102 45790 23154
rect 46834 23102 46846 23154
rect 46898 23102 46910 23154
rect 48738 23102 48750 23154
rect 48802 23102 48814 23154
rect 49858 23102 49870 23154
rect 49922 23102 49934 23154
rect 52210 23102 52222 23154
rect 52274 23102 52286 23154
rect 52882 23102 52894 23154
rect 52946 23102 52958 23154
rect 54562 23102 54574 23154
rect 54626 23102 54638 23154
rect 58594 23102 58606 23154
rect 58658 23102 58670 23154
rect 59042 23102 59054 23154
rect 59106 23102 59118 23154
rect 59938 23102 59950 23154
rect 60002 23102 60014 23154
rect 38334 23090 38386 23102
rect 40350 23090 40402 23102
rect 42366 23090 42418 23102
rect 44942 23090 44994 23102
rect 47854 23090 47906 23102
rect 51550 23090 51602 23102
rect 56926 23090 56978 23102
rect 3166 23042 3218 23054
rect 8094 23042 8146 23054
rect 3826 22990 3838 23042
rect 3890 22990 3902 23042
rect 3166 22978 3218 22990
rect 8094 22978 8146 22990
rect 8990 23042 9042 23054
rect 8990 22978 9042 22990
rect 10558 23042 10610 23054
rect 48190 23042 48242 23054
rect 57150 23042 57202 23054
rect 14690 22990 14702 23042
rect 14754 22990 14766 23042
rect 21634 22990 21646 23042
rect 21698 22990 21710 23042
rect 24434 22990 24446 23042
rect 24498 22990 24510 23042
rect 45938 22990 45950 23042
rect 46002 22990 46014 23042
rect 54786 22990 54798 23042
rect 54850 22990 54862 23042
rect 57810 22990 57822 23042
rect 57874 22990 57886 23042
rect 10558 22978 10610 22990
rect 48190 22978 48242 22990
rect 57150 22978 57202 22990
rect 13470 22930 13522 22942
rect 13470 22866 13522 22878
rect 16046 22930 16098 22942
rect 16046 22866 16098 22878
rect 17502 22930 17554 22942
rect 17502 22866 17554 22878
rect 19070 22930 19122 22942
rect 33070 22930 33122 22942
rect 29250 22878 29262 22930
rect 29314 22878 29326 22930
rect 19070 22866 19122 22878
rect 33070 22866 33122 22878
rect 37998 22930 38050 22942
rect 62078 22930 62130 22942
rect 41010 22878 41022 22930
rect 41074 22878 41086 22930
rect 52770 22878 52782 22930
rect 52834 22878 52846 22930
rect 37998 22866 38050 22878
rect 62078 22866 62130 22878
rect 1344 22762 62608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 62608 22762
rect 1344 22676 62608 22710
rect 22318 22594 22370 22606
rect 22318 22530 22370 22542
rect 24782 22594 24834 22606
rect 32622 22594 32674 22606
rect 25666 22542 25678 22594
rect 25730 22542 25742 22594
rect 24782 22530 24834 22542
rect 32622 22530 32674 22542
rect 39006 22594 39058 22606
rect 39006 22530 39058 22542
rect 49982 22594 50034 22606
rect 60622 22594 60674 22606
rect 51090 22542 51102 22594
rect 51154 22542 51166 22594
rect 49982 22530 50034 22542
rect 60622 22530 60674 22542
rect 60958 22594 61010 22606
rect 60958 22530 61010 22542
rect 9102 22482 9154 22494
rect 12462 22482 12514 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 9538 22430 9550 22482
rect 9602 22430 9614 22482
rect 10658 22430 10670 22482
rect 10722 22430 10734 22482
rect 9102 22418 9154 22430
rect 12462 22418 12514 22430
rect 13582 22482 13634 22494
rect 13582 22418 13634 22430
rect 14030 22482 14082 22494
rect 14030 22418 14082 22430
rect 14926 22482 14978 22494
rect 45278 22482 45330 22494
rect 18386 22430 18398 22482
rect 18450 22430 18462 22482
rect 20514 22430 20526 22482
rect 20578 22430 20590 22482
rect 21410 22430 21422 22482
rect 21474 22430 21486 22482
rect 29362 22430 29374 22482
rect 29426 22430 29438 22482
rect 39778 22430 39790 22482
rect 39842 22430 39854 22482
rect 14926 22418 14978 22430
rect 45278 22418 45330 22430
rect 45838 22482 45890 22494
rect 45838 22418 45890 22430
rect 47966 22482 48018 22494
rect 47966 22418 48018 22430
rect 54238 22482 54290 22494
rect 54238 22418 54290 22430
rect 13022 22370 13074 22382
rect 5618 22318 5630 22370
rect 5682 22318 5694 22370
rect 6962 22318 6974 22370
rect 7026 22318 7038 22370
rect 8642 22318 8654 22370
rect 8706 22318 8718 22370
rect 9762 22318 9774 22370
rect 9826 22318 9838 22370
rect 10210 22318 10222 22370
rect 10274 22318 10286 22370
rect 10994 22318 11006 22370
rect 11058 22318 11070 22370
rect 11778 22318 11790 22370
rect 11842 22318 11854 22370
rect 13022 22306 13074 22318
rect 13918 22370 13970 22382
rect 13918 22306 13970 22318
rect 14142 22370 14194 22382
rect 14142 22306 14194 22318
rect 14478 22370 14530 22382
rect 14478 22306 14530 22318
rect 15038 22370 15090 22382
rect 15038 22306 15090 22318
rect 15374 22370 15426 22382
rect 21870 22370 21922 22382
rect 15698 22318 15710 22370
rect 15762 22318 15774 22370
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 15374 22306 15426 22318
rect 21870 22306 21922 22318
rect 22430 22370 22482 22382
rect 32062 22370 32114 22382
rect 25218 22318 25230 22370
rect 25282 22318 25294 22370
rect 26450 22318 26462 22370
rect 26514 22318 26526 22370
rect 27346 22318 27358 22370
rect 27410 22318 27422 22370
rect 30034 22318 30046 22370
rect 30098 22318 30110 22370
rect 30482 22318 30494 22370
rect 30546 22318 30558 22370
rect 31490 22318 31502 22370
rect 31554 22318 31566 22370
rect 22430 22306 22482 22318
rect 32062 22306 32114 22318
rect 32398 22370 32450 22382
rect 32398 22306 32450 22318
rect 33518 22370 33570 22382
rect 35198 22370 35250 22382
rect 33842 22318 33854 22370
rect 33906 22318 33918 22370
rect 33518 22306 33570 22318
rect 35198 22306 35250 22318
rect 35870 22370 35922 22382
rect 35870 22306 35922 22318
rect 36318 22370 36370 22382
rect 45166 22370 45218 22382
rect 39442 22318 39454 22370
rect 39506 22318 39518 22370
rect 40674 22318 40686 22370
rect 40738 22318 40750 22370
rect 41682 22318 41694 22370
rect 41746 22318 41758 22370
rect 44818 22318 44830 22370
rect 44882 22318 44894 22370
rect 36318 22306 36370 22318
rect 45166 22306 45218 22318
rect 45390 22370 45442 22382
rect 47854 22370 47906 22382
rect 49758 22370 49810 22382
rect 47618 22318 47630 22370
rect 47682 22318 47694 22370
rect 49298 22318 49310 22370
rect 49362 22318 49374 22370
rect 45390 22306 45442 22318
rect 47854 22306 47906 22318
rect 49758 22306 49810 22318
rect 50542 22370 50594 22382
rect 53454 22370 53506 22382
rect 52658 22318 52670 22370
rect 52722 22318 52734 22370
rect 50542 22306 50594 22318
rect 53454 22306 53506 22318
rect 53790 22370 53842 22382
rect 53790 22306 53842 22318
rect 54350 22370 54402 22382
rect 58158 22370 58210 22382
rect 57474 22318 57486 22370
rect 57538 22318 57550 22370
rect 54350 22306 54402 22318
rect 58158 22306 58210 22318
rect 12350 22258 12402 22270
rect 3490 22206 3502 22258
rect 3554 22206 3566 22258
rect 6402 22206 6414 22258
rect 6466 22206 6478 22258
rect 7522 22206 7534 22258
rect 7586 22206 7598 22258
rect 9538 22206 9550 22258
rect 9602 22206 9614 22258
rect 10882 22206 10894 22258
rect 10946 22206 10958 22258
rect 12350 22194 12402 22206
rect 14814 22258 14866 22270
rect 22318 22258 22370 22270
rect 31838 22258 31890 22270
rect 17266 22206 17278 22258
rect 17330 22206 17342 22258
rect 28018 22206 28030 22258
rect 28082 22206 28094 22258
rect 14814 22194 14866 22206
rect 22318 22194 22370 22206
rect 31838 22194 31890 22206
rect 32174 22258 32226 22270
rect 32174 22194 32226 22206
rect 33070 22258 33122 22270
rect 53118 22258 53170 22270
rect 33282 22206 33294 22258
rect 33346 22206 33358 22258
rect 34514 22206 34526 22258
rect 34578 22206 34590 22258
rect 37538 22206 37550 22258
rect 37602 22206 37614 22258
rect 40898 22206 40910 22258
rect 40962 22206 40974 22258
rect 42690 22206 42702 22258
rect 42754 22206 42766 22258
rect 48850 22206 48862 22258
rect 48914 22206 48926 22258
rect 51538 22206 51550 22258
rect 51602 22206 51614 22258
rect 33070 22194 33122 22206
rect 53118 22194 53170 22206
rect 54014 22258 54066 22270
rect 55122 22206 55134 22258
rect 55186 22206 55198 22258
rect 57250 22206 57262 22258
rect 57314 22206 57326 22258
rect 59378 22206 59390 22258
rect 59442 22206 59454 22258
rect 61282 22206 61294 22258
rect 61346 22206 61358 22258
rect 61506 22206 61518 22258
rect 61570 22206 61582 22258
rect 54014 22194 54066 22206
rect 1710 22146 1762 22158
rect 1710 22082 1762 22094
rect 5070 22146 5122 22158
rect 12574 22146 12626 22158
rect 12002 22094 12014 22146
rect 12066 22094 12078 22146
rect 5070 22082 5122 22094
rect 12574 22082 12626 22094
rect 15822 22146 15874 22158
rect 15822 22082 15874 22094
rect 16942 22146 16994 22158
rect 33854 22146 33906 22158
rect 23426 22094 23438 22146
rect 23490 22094 23502 22146
rect 16942 22082 16994 22094
rect 33854 22082 33906 22094
rect 34190 22146 34242 22158
rect 34190 22082 34242 22094
rect 34862 22146 34914 22158
rect 34862 22082 34914 22094
rect 35982 22146 36034 22158
rect 35982 22082 36034 22094
rect 36430 22146 36482 22158
rect 44158 22146 44210 22158
rect 41570 22094 41582 22146
rect 41634 22094 41646 22146
rect 36430 22082 36482 22094
rect 44158 22082 44210 22094
rect 52110 22146 52162 22158
rect 52110 22082 52162 22094
rect 53230 22146 53282 22158
rect 53230 22082 53282 22094
rect 53342 22146 53394 22158
rect 53342 22082 53394 22094
rect 57038 22146 57090 22158
rect 57038 22082 57090 22094
rect 1344 21978 62608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 62608 21978
rect 1344 21892 62608 21926
rect 4622 21810 4674 21822
rect 2370 21758 2382 21810
rect 2434 21758 2446 21810
rect 4622 21746 4674 21758
rect 4846 21810 4898 21822
rect 4846 21746 4898 21758
rect 7646 21810 7698 21822
rect 14926 21810 14978 21822
rect 19518 21810 19570 21822
rect 11330 21758 11342 21810
rect 11394 21758 11406 21810
rect 17714 21758 17726 21810
rect 17778 21758 17790 21810
rect 7646 21746 7698 21758
rect 14926 21746 14978 21758
rect 19518 21746 19570 21758
rect 19630 21810 19682 21822
rect 19630 21746 19682 21758
rect 20302 21810 20354 21822
rect 20302 21746 20354 21758
rect 22654 21810 22706 21822
rect 22654 21746 22706 21758
rect 23886 21810 23938 21822
rect 31054 21810 31106 21822
rect 29698 21758 29710 21810
rect 29762 21758 29774 21810
rect 23886 21746 23938 21758
rect 31054 21746 31106 21758
rect 33294 21810 33346 21822
rect 41918 21810 41970 21822
rect 33954 21758 33966 21810
rect 34018 21758 34030 21810
rect 40002 21758 40014 21810
rect 40066 21758 40078 21810
rect 41570 21758 41582 21810
rect 41634 21758 41646 21810
rect 33294 21746 33346 21758
rect 41918 21746 41970 21758
rect 42142 21810 42194 21822
rect 44494 21810 44546 21822
rect 45838 21810 45890 21822
rect 43250 21758 43262 21810
rect 43314 21758 43326 21810
rect 45378 21758 45390 21810
rect 45442 21758 45454 21810
rect 42142 21746 42194 21758
rect 44494 21746 44546 21758
rect 45838 21746 45890 21758
rect 46622 21810 46674 21822
rect 46622 21746 46674 21758
rect 55358 21810 55410 21822
rect 55682 21758 55694 21810
rect 55746 21758 55758 21810
rect 61506 21758 61518 21810
rect 61570 21758 61582 21810
rect 55358 21746 55410 21758
rect 3502 21698 3554 21710
rect 3502 21634 3554 21646
rect 4398 21698 4450 21710
rect 4398 21634 4450 21646
rect 5182 21698 5234 21710
rect 19406 21698 19458 21710
rect 21310 21698 21362 21710
rect 8306 21646 8318 21698
rect 8370 21646 8382 21698
rect 8754 21646 8766 21698
rect 8818 21646 8830 21698
rect 11778 21646 11790 21698
rect 11842 21646 11854 21698
rect 15586 21646 15598 21698
rect 15650 21646 15662 21698
rect 17602 21646 17614 21698
rect 17666 21646 17678 21698
rect 18386 21646 18398 21698
rect 18450 21646 18462 21698
rect 19954 21646 19966 21698
rect 20018 21646 20030 21698
rect 20962 21646 20974 21698
rect 21026 21646 21038 21698
rect 5182 21634 5234 21646
rect 19406 21634 19458 21646
rect 21310 21634 21362 21646
rect 21646 21698 21698 21710
rect 21646 21634 21698 21646
rect 23550 21698 23602 21710
rect 23550 21634 23602 21646
rect 23662 21698 23714 21710
rect 30270 21698 30322 21710
rect 33630 21698 33682 21710
rect 26450 21646 26462 21698
rect 26514 21646 26526 21698
rect 28018 21646 28030 21698
rect 28082 21646 28094 21698
rect 31602 21646 31614 21698
rect 31666 21646 31678 21698
rect 32162 21646 32174 21698
rect 32226 21646 32238 21698
rect 23662 21634 23714 21646
rect 30270 21634 30322 21646
rect 33630 21634 33682 21646
rect 39678 21698 39730 21710
rect 39678 21634 39730 21646
rect 42366 21698 42418 21710
rect 42366 21634 42418 21646
rect 43822 21698 43874 21710
rect 48750 21698 48802 21710
rect 44146 21646 44158 21698
rect 44210 21646 44222 21698
rect 47730 21646 47742 21698
rect 47794 21646 47806 21698
rect 43822 21634 43874 21646
rect 48750 21634 48802 21646
rect 48974 21698 49026 21710
rect 48974 21634 49026 21646
rect 49086 21698 49138 21710
rect 59614 21698 59666 21710
rect 49298 21646 49310 21698
rect 49362 21646 49374 21698
rect 51314 21646 51326 21698
rect 51378 21646 51390 21698
rect 58370 21646 58382 21698
rect 58434 21646 58446 21698
rect 49086 21634 49138 21646
rect 59614 21634 59666 21646
rect 6190 21586 6242 21598
rect 13582 21586 13634 21598
rect 5394 21534 5406 21586
rect 5458 21534 5470 21586
rect 6626 21534 6638 21586
rect 6690 21534 6702 21586
rect 11106 21534 11118 21586
rect 11170 21534 11182 21586
rect 12002 21534 12014 21586
rect 12066 21534 12078 21586
rect 6190 21522 6242 21534
rect 13582 21522 13634 21534
rect 13806 21586 13858 21598
rect 13806 21522 13858 21534
rect 14478 21586 14530 21598
rect 14478 21522 14530 21534
rect 14702 21586 14754 21598
rect 17390 21586 17442 21598
rect 20638 21586 20690 21598
rect 15474 21534 15486 21586
rect 15538 21534 15550 21586
rect 18834 21534 18846 21586
rect 18898 21534 18910 21586
rect 19170 21534 19182 21586
rect 19234 21534 19246 21586
rect 14702 21522 14754 21534
rect 17390 21522 17442 21534
rect 20638 21522 20690 21534
rect 22318 21586 22370 21598
rect 22318 21522 22370 21534
rect 22878 21586 22930 21598
rect 22878 21522 22930 21534
rect 23326 21586 23378 21598
rect 25342 21586 25394 21598
rect 24546 21534 24558 21586
rect 24610 21534 24622 21586
rect 23326 21522 23378 21534
rect 25342 21522 25394 21534
rect 33070 21586 33122 21598
rect 33070 21522 33122 21534
rect 33294 21586 33346 21598
rect 33294 21522 33346 21534
rect 34526 21586 34578 21598
rect 39118 21586 39170 21598
rect 41022 21586 41074 21598
rect 34962 21534 34974 21586
rect 35026 21534 35038 21586
rect 35746 21534 35758 21586
rect 35810 21534 35822 21586
rect 38658 21534 38670 21586
rect 38722 21534 38734 21586
rect 40226 21534 40238 21586
rect 40290 21534 40302 21586
rect 34526 21522 34578 21534
rect 39118 21522 39170 21534
rect 41022 21522 41074 21534
rect 42030 21586 42082 21598
rect 42030 21522 42082 21534
rect 43598 21586 43650 21598
rect 43598 21522 43650 21534
rect 44830 21586 44882 21598
rect 44830 21522 44882 21534
rect 45054 21586 45106 21598
rect 46958 21586 47010 21598
rect 53006 21586 53058 21598
rect 45714 21534 45726 21586
rect 45778 21534 45790 21586
rect 47618 21534 47630 21586
rect 47682 21534 47694 21586
rect 49858 21534 49870 21586
rect 49922 21534 49934 21586
rect 45054 21522 45106 21534
rect 46958 21522 47010 21534
rect 53006 21522 53058 21534
rect 54686 21586 54738 21598
rect 54686 21522 54738 21534
rect 55022 21586 55074 21598
rect 55022 21522 55074 21534
rect 55246 21586 55298 21598
rect 59278 21586 59330 21598
rect 55906 21534 55918 21586
rect 55970 21534 55982 21586
rect 57250 21534 57262 21586
rect 57314 21534 57326 21586
rect 58258 21534 58270 21586
rect 58322 21534 58334 21586
rect 59042 21534 59054 21586
rect 59106 21534 59118 21586
rect 55246 21522 55298 21534
rect 59278 21522 59330 21534
rect 4734 21474 4786 21486
rect 9886 21474 9938 21486
rect 6066 21422 6078 21474
rect 6130 21422 6142 21474
rect 4734 21410 4786 21422
rect 9886 21410 9938 21422
rect 10782 21474 10834 21486
rect 10782 21410 10834 21422
rect 12574 21474 12626 21486
rect 14590 21474 14642 21486
rect 22766 21474 22818 21486
rect 29262 21474 29314 21486
rect 14130 21422 14142 21474
rect 14194 21422 14206 21474
rect 21970 21422 21982 21474
rect 22034 21422 22046 21474
rect 24210 21422 24222 21474
rect 24274 21422 24286 21474
rect 12574 21410 12626 21422
rect 14590 21410 14642 21422
rect 22766 21410 22818 21422
rect 29262 21410 29314 21422
rect 30046 21474 30098 21486
rect 30046 21410 30098 21422
rect 34302 21474 34354 21486
rect 38222 21474 38274 21486
rect 37874 21422 37886 21474
rect 37938 21422 37950 21474
rect 34302 21410 34354 21422
rect 38222 21410 38274 21422
rect 42926 21474 42978 21486
rect 42926 21410 42978 21422
rect 48862 21474 48914 21486
rect 54014 21474 54066 21486
rect 59502 21474 59554 21486
rect 49970 21422 49982 21474
rect 50034 21422 50046 21474
rect 53442 21422 53454 21474
rect 53506 21422 53518 21474
rect 57586 21422 57598 21474
rect 57650 21422 57662 21474
rect 58370 21422 58382 21474
rect 58434 21422 58446 21474
rect 48862 21410 48914 21422
rect 54014 21410 54066 21422
rect 59502 21410 59554 21422
rect 7982 21362 8034 21374
rect 10558 21362 10610 21374
rect 10210 21310 10222 21362
rect 10274 21310 10286 21362
rect 7982 21298 8034 21310
rect 10558 21298 10610 21310
rect 12798 21362 12850 21374
rect 12798 21298 12850 21310
rect 13134 21362 13186 21374
rect 13134 21298 13186 21310
rect 16270 21362 16322 21374
rect 16270 21298 16322 21310
rect 16606 21362 16658 21374
rect 16606 21298 16658 21310
rect 31390 21362 31442 21374
rect 31390 21298 31442 21310
rect 41246 21362 41298 21374
rect 41246 21298 41298 21310
rect 52558 21362 52610 21374
rect 52558 21298 52610 21310
rect 54126 21362 54178 21374
rect 54126 21298 54178 21310
rect 54462 21362 54514 21374
rect 60174 21362 60226 21374
rect 59042 21310 59054 21362
rect 59106 21310 59118 21362
rect 54462 21298 54514 21310
rect 60174 21298 60226 21310
rect 1344 21194 62608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 62608 21194
rect 1344 21108 62608 21142
rect 3278 21026 3330 21038
rect 3278 20962 3330 20974
rect 4174 21026 4226 21038
rect 4174 20962 4226 20974
rect 4510 21026 4562 21038
rect 4510 20962 4562 20974
rect 5630 21026 5682 21038
rect 5630 20962 5682 20974
rect 12014 21026 12066 21038
rect 27134 21026 27186 21038
rect 17378 20974 17390 21026
rect 17442 20974 17454 21026
rect 12014 20962 12066 20974
rect 27134 20962 27186 20974
rect 27470 21026 27522 21038
rect 27470 20962 27522 20974
rect 29374 21026 29426 21038
rect 60510 21026 60562 21038
rect 61966 21026 62018 21038
rect 48290 20974 48302 21026
rect 48354 20974 48366 21026
rect 58594 20974 58606 21026
rect 58658 20974 58670 21026
rect 61618 20974 61630 21026
rect 61682 20974 61694 21026
rect 29374 20962 29426 20974
rect 60510 20962 60562 20974
rect 61966 20962 62018 20974
rect 5742 20914 5794 20926
rect 9214 20914 9266 20926
rect 7746 20862 7758 20914
rect 7810 20862 7822 20914
rect 5742 20850 5794 20862
rect 9214 20850 9266 20862
rect 12462 20914 12514 20926
rect 15598 20914 15650 20926
rect 21310 20914 21362 20926
rect 29934 20914 29986 20926
rect 31950 20914 32002 20926
rect 39454 20914 39506 20926
rect 14018 20862 14030 20914
rect 14082 20862 14094 20914
rect 17826 20862 17838 20914
rect 17890 20862 17902 20914
rect 22530 20862 22542 20914
rect 22594 20862 22606 20914
rect 24658 20862 24670 20914
rect 24722 20862 24734 20914
rect 31714 20862 31726 20914
rect 31778 20862 31790 20914
rect 33058 20862 33070 20914
rect 33122 20862 33134 20914
rect 35186 20862 35198 20914
rect 35250 20862 35262 20914
rect 36306 20862 36318 20914
rect 36370 20862 36382 20914
rect 38434 20862 38446 20914
rect 38498 20862 38510 20914
rect 12462 20850 12514 20862
rect 15598 20850 15650 20862
rect 21310 20850 21362 20862
rect 29934 20850 29986 20862
rect 31950 20850 32002 20862
rect 39454 20850 39506 20862
rect 49534 20914 49586 20926
rect 54238 20914 54290 20926
rect 53106 20862 53118 20914
rect 53170 20862 53182 20914
rect 49534 20850 49586 20862
rect 54238 20850 54290 20862
rect 62190 20914 62242 20926
rect 62190 20850 62242 20862
rect 1822 20802 1874 20814
rect 3054 20802 3106 20814
rect 2706 20750 2718 20802
rect 2770 20750 2782 20802
rect 1822 20738 1874 20750
rect 3054 20738 3106 20750
rect 3950 20802 4002 20814
rect 3950 20738 4002 20750
rect 4846 20802 4898 20814
rect 4846 20738 4898 20750
rect 6974 20802 7026 20814
rect 8990 20802 9042 20814
rect 7858 20750 7870 20802
rect 7922 20750 7934 20802
rect 8082 20750 8094 20802
rect 8146 20750 8158 20802
rect 6974 20738 7026 20750
rect 8990 20738 9042 20750
rect 9550 20802 9602 20814
rect 20414 20802 20466 20814
rect 13682 20750 13694 20802
rect 13746 20750 13758 20802
rect 14578 20750 14590 20802
rect 14642 20750 14654 20802
rect 17266 20750 17278 20802
rect 17330 20750 17342 20802
rect 17938 20750 17950 20802
rect 18002 20750 18014 20802
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 9550 20738 9602 20750
rect 20414 20738 20466 20750
rect 20638 20802 20690 20814
rect 20638 20738 20690 20750
rect 21422 20802 21474 20814
rect 24894 20802 24946 20814
rect 21858 20750 21870 20802
rect 21922 20750 21934 20802
rect 21422 20738 21474 20750
rect 24894 20738 24946 20750
rect 25678 20802 25730 20814
rect 31054 20802 31106 20814
rect 40574 20802 40626 20814
rect 27906 20750 27918 20802
rect 27970 20750 27982 20802
rect 29250 20750 29262 20802
rect 29314 20750 29326 20802
rect 31602 20750 31614 20802
rect 31666 20750 31678 20802
rect 32386 20750 32398 20802
rect 32450 20750 32462 20802
rect 36194 20750 36206 20802
rect 36258 20750 36270 20802
rect 37090 20750 37102 20802
rect 37154 20750 37166 20802
rect 38098 20750 38110 20802
rect 38162 20750 38174 20802
rect 38994 20750 39006 20802
rect 39058 20750 39070 20802
rect 40114 20750 40126 20802
rect 40178 20750 40190 20802
rect 25678 20738 25730 20750
rect 31054 20738 31106 20750
rect 40574 20738 40626 20750
rect 40910 20802 40962 20814
rect 40910 20738 40962 20750
rect 43038 20802 43090 20814
rect 53902 20802 53954 20814
rect 45154 20750 45166 20802
rect 45218 20750 45230 20802
rect 46274 20750 46286 20802
rect 46338 20750 46350 20802
rect 47618 20750 47630 20802
rect 47682 20750 47694 20802
rect 52658 20750 52670 20802
rect 52722 20750 52734 20802
rect 43038 20738 43090 20750
rect 53902 20738 53954 20750
rect 54014 20802 54066 20814
rect 54014 20738 54066 20750
rect 54462 20802 54514 20814
rect 56142 20802 56194 20814
rect 55682 20750 55694 20802
rect 55746 20750 55758 20802
rect 54462 20738 54514 20750
rect 56142 20738 56194 20750
rect 56366 20802 56418 20814
rect 58830 20802 58882 20814
rect 56578 20750 56590 20802
rect 56642 20750 56654 20802
rect 58370 20750 58382 20802
rect 58434 20750 58446 20802
rect 56366 20738 56418 20750
rect 58830 20738 58882 20750
rect 59054 20802 59106 20814
rect 59054 20738 59106 20750
rect 59166 20802 59218 20814
rect 59166 20738 59218 20750
rect 59838 20802 59890 20814
rect 59838 20738 59890 20750
rect 60734 20802 60786 20814
rect 60734 20738 60786 20750
rect 8318 20690 8370 20702
rect 6290 20638 6302 20690
rect 6354 20638 6366 20690
rect 6626 20638 6638 20690
rect 6690 20638 6702 20690
rect 8318 20626 8370 20638
rect 9438 20690 9490 20702
rect 15374 20690 15426 20702
rect 14466 20638 14478 20690
rect 14530 20638 14542 20690
rect 15138 20638 15150 20690
rect 15202 20638 15214 20690
rect 9438 20626 9490 20638
rect 15374 20626 15426 20638
rect 15486 20690 15538 20702
rect 15486 20626 15538 20638
rect 15710 20690 15762 20702
rect 25118 20690 25170 20702
rect 16594 20638 16606 20690
rect 16658 20638 16670 20690
rect 15710 20626 15762 20638
rect 25118 20626 25170 20638
rect 25230 20690 25282 20702
rect 29822 20690 29874 20702
rect 26114 20638 26126 20690
rect 26178 20638 26190 20690
rect 26562 20638 26574 20690
rect 26626 20638 26638 20690
rect 28242 20638 28254 20690
rect 28306 20638 28318 20690
rect 25230 20626 25282 20638
rect 29822 20626 29874 20638
rect 30158 20690 30210 20702
rect 30158 20626 30210 20638
rect 30382 20690 30434 20702
rect 30382 20626 30434 20638
rect 30718 20690 30770 20702
rect 30718 20626 30770 20638
rect 31278 20690 31330 20702
rect 31278 20626 31330 20638
rect 35870 20690 35922 20702
rect 35870 20626 35922 20638
rect 40798 20690 40850 20702
rect 40798 20626 40850 20638
rect 41358 20690 41410 20702
rect 56254 20690 56306 20702
rect 42242 20638 42254 20690
rect 42306 20638 42318 20690
rect 42802 20638 42814 20690
rect 42866 20638 42878 20690
rect 47506 20638 47518 20690
rect 47570 20638 47582 20690
rect 50978 20638 50990 20690
rect 51042 20638 51054 20690
rect 59490 20638 59502 20690
rect 59554 20638 59566 20690
rect 41358 20626 41410 20638
rect 56254 20626 56306 20638
rect 1934 20578 1986 20590
rect 1934 20514 1986 20526
rect 2158 20578 2210 20590
rect 2158 20514 2210 20526
rect 2606 20578 2658 20590
rect 4958 20578 5010 20590
rect 3602 20526 3614 20578
rect 3666 20526 3678 20578
rect 2606 20514 2658 20526
rect 4958 20514 5010 20526
rect 5182 20578 5234 20590
rect 5182 20514 5234 20526
rect 7310 20578 7362 20590
rect 7310 20514 7362 20526
rect 8542 20578 8594 20590
rect 12574 20578 12626 20590
rect 10658 20526 10670 20578
rect 10722 20526 10734 20578
rect 8542 20514 8594 20526
rect 12574 20514 12626 20526
rect 20526 20578 20578 20590
rect 30942 20578 30994 20590
rect 25890 20526 25902 20578
rect 25954 20526 25966 20578
rect 20526 20514 20578 20526
rect 30942 20514 30994 20526
rect 35534 20578 35586 20590
rect 35534 20514 35586 20526
rect 35758 20578 35810 20590
rect 35758 20514 35810 20526
rect 37214 20578 37266 20590
rect 41694 20578 41746 20590
rect 40338 20526 40350 20578
rect 40402 20526 40414 20578
rect 37214 20514 37266 20526
rect 41694 20514 41746 20526
rect 43374 20578 43426 20590
rect 43374 20514 43426 20526
rect 43822 20578 43874 20590
rect 48750 20578 48802 20590
rect 51998 20578 52050 20590
rect 44146 20526 44158 20578
rect 44210 20526 44222 20578
rect 49074 20526 49086 20578
rect 49138 20526 49150 20578
rect 43822 20514 43874 20526
rect 48750 20514 48802 20526
rect 51998 20514 52050 20526
rect 60958 20578 61010 20590
rect 60958 20514 61010 20526
rect 61070 20578 61122 20590
rect 61070 20514 61122 20526
rect 61182 20578 61234 20590
rect 61182 20514 61234 20526
rect 1344 20410 62608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 62608 20410
rect 1344 20324 62608 20358
rect 43038 20242 43090 20254
rect 57598 20242 57650 20254
rect 44146 20190 44158 20242
rect 44210 20190 44222 20242
rect 50530 20190 50542 20242
rect 50594 20190 50606 20242
rect 43038 20178 43090 20190
rect 57598 20178 57650 20190
rect 5182 20130 5234 20142
rect 2482 20078 2494 20130
rect 2546 20078 2558 20130
rect 5182 20066 5234 20078
rect 5294 20130 5346 20142
rect 5294 20066 5346 20078
rect 5518 20130 5570 20142
rect 5518 20066 5570 20078
rect 6078 20130 6130 20142
rect 7758 20130 7810 20142
rect 7522 20078 7534 20130
rect 7586 20078 7598 20130
rect 6078 20066 6130 20078
rect 7758 20066 7810 20078
rect 8430 20130 8482 20142
rect 8430 20066 8482 20078
rect 8766 20130 8818 20142
rect 8766 20066 8818 20078
rect 8990 20130 9042 20142
rect 8990 20066 9042 20078
rect 11230 20130 11282 20142
rect 25902 20130 25954 20142
rect 30494 20130 30546 20142
rect 11778 20078 11790 20130
rect 11842 20078 11854 20130
rect 22082 20078 22094 20130
rect 22146 20078 22158 20130
rect 29698 20078 29710 20130
rect 29762 20078 29774 20130
rect 11230 20066 11282 20078
rect 25902 20066 25954 20078
rect 30494 20066 30546 20078
rect 30718 20130 30770 20142
rect 45950 20130 46002 20142
rect 31042 20078 31054 20130
rect 31106 20078 31118 20130
rect 31714 20078 31726 20130
rect 31778 20078 31790 20130
rect 34850 20078 34862 20130
rect 34914 20078 34926 20130
rect 39890 20078 39902 20130
rect 39954 20078 39966 20130
rect 41794 20078 41806 20130
rect 41858 20078 41870 20130
rect 30718 20066 30770 20078
rect 45950 20066 46002 20078
rect 47854 20130 47906 20142
rect 47854 20066 47906 20078
rect 47966 20130 48018 20142
rect 47966 20066 48018 20078
rect 48862 20130 48914 20142
rect 48862 20066 48914 20078
rect 51662 20130 51714 20142
rect 51662 20066 51714 20078
rect 52222 20130 52274 20142
rect 54350 20130 54402 20142
rect 53890 20078 53902 20130
rect 53954 20078 53966 20130
rect 52222 20066 52274 20078
rect 54350 20066 54402 20078
rect 54574 20130 54626 20142
rect 54574 20066 54626 20078
rect 57710 20130 57762 20142
rect 61518 20130 61570 20142
rect 58930 20078 58942 20130
rect 58994 20078 59006 20130
rect 57710 20066 57762 20078
rect 61518 20066 61570 20078
rect 8542 20018 8594 20030
rect 1698 19966 1710 20018
rect 1762 19966 1774 20018
rect 5730 19966 5742 20018
rect 5794 19966 5806 20018
rect 6290 19966 6302 20018
rect 6354 19966 6366 20018
rect 7186 19966 7198 20018
rect 7250 19966 7262 20018
rect 8542 19954 8594 19966
rect 9550 20018 9602 20030
rect 15374 20018 15426 20030
rect 20526 20018 20578 20030
rect 24782 20018 24834 20030
rect 28254 20018 28306 20030
rect 30382 20018 30434 20030
rect 45502 20018 45554 20030
rect 9762 19966 9774 20018
rect 9826 19966 9838 20018
rect 10658 19966 10670 20018
rect 10722 19966 10734 20018
rect 12002 19966 12014 20018
rect 12066 19966 12078 20018
rect 12674 19966 12686 20018
rect 12738 19966 12750 20018
rect 13458 19966 13470 20018
rect 13522 19966 13534 20018
rect 14690 19966 14702 20018
rect 14754 19966 14766 20018
rect 16482 19966 16494 20018
rect 16546 19966 16558 20018
rect 17378 19966 17390 20018
rect 17442 19966 17454 20018
rect 20290 19966 20302 20018
rect 20354 19966 20366 20018
rect 21410 19966 21422 20018
rect 21474 19966 21486 20018
rect 25442 19966 25454 20018
rect 25506 19966 25518 20018
rect 26338 19966 26350 20018
rect 26402 19966 26414 20018
rect 29810 19966 29822 20018
rect 29874 19966 29886 20018
rect 30930 19966 30942 20018
rect 30994 19966 31006 20018
rect 31938 19966 31950 20018
rect 32002 19966 32014 20018
rect 32498 19966 32510 20018
rect 32562 19966 32574 20018
rect 33618 19966 33630 20018
rect 33682 19966 33694 20018
rect 34178 19966 34190 20018
rect 34242 19966 34254 20018
rect 36082 19966 36094 20018
rect 36146 19966 36158 20018
rect 37314 19966 37326 20018
rect 37378 19966 37390 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 39106 19966 39118 20018
rect 39170 19966 39182 20018
rect 39442 19966 39454 20018
rect 39506 19966 39518 20018
rect 9550 19954 9602 19966
rect 15374 19954 15426 19966
rect 20526 19954 20578 19966
rect 24782 19954 24834 19966
rect 28254 19954 28306 19966
rect 30382 19954 30434 19966
rect 45502 19954 45554 19966
rect 47070 20018 47122 20030
rect 47070 19954 47122 19966
rect 48750 20018 48802 20030
rect 48750 19954 48802 19966
rect 48974 20018 49026 20030
rect 55022 20018 55074 20030
rect 61406 20018 61458 20030
rect 49298 19966 49310 20018
rect 49362 19966 49374 20018
rect 53666 19966 53678 20018
rect 53730 19966 53742 20018
rect 55906 19966 55918 20018
rect 55970 19966 55982 20018
rect 57026 19966 57038 20018
rect 57090 19966 57102 20018
rect 58146 19966 58158 20018
rect 58210 19966 58222 20018
rect 48974 19954 49026 19966
rect 55022 19954 55074 19966
rect 61406 19954 61458 19966
rect 61630 20018 61682 20030
rect 61630 19954 61682 19966
rect 61966 20018 62018 20030
rect 61966 19954 62018 19966
rect 12238 19906 12290 19918
rect 4610 19854 4622 19906
rect 4674 19854 4686 19906
rect 10098 19854 10110 19906
rect 10162 19854 10174 19906
rect 12238 19842 12290 19854
rect 12350 19906 12402 19918
rect 20078 19906 20130 19918
rect 27246 19906 27298 19918
rect 18050 19854 18062 19906
rect 18114 19854 18126 19906
rect 24210 19854 24222 19906
rect 24274 19854 24286 19906
rect 25554 19854 25566 19906
rect 25618 19854 25630 19906
rect 26226 19854 26238 19906
rect 26290 19854 26302 19906
rect 12350 19842 12402 19854
rect 20078 19842 20130 19854
rect 27246 19842 27298 19854
rect 27694 19906 27746 19918
rect 46846 19906 46898 19918
rect 33506 19854 33518 19906
rect 33570 19854 33582 19906
rect 46386 19854 46398 19906
rect 46450 19854 46462 19906
rect 27694 19842 27746 19854
rect 46846 19842 46898 19854
rect 54462 19906 54514 19918
rect 56590 19906 56642 19918
rect 55458 19854 55470 19906
rect 55522 19854 55534 19906
rect 61058 19854 61070 19906
rect 61122 19854 61134 19906
rect 54462 19842 54514 19854
rect 56590 19842 56642 19854
rect 16606 19794 16658 19806
rect 16606 19730 16658 19742
rect 27358 19794 27410 19806
rect 27358 19730 27410 19742
rect 28702 19794 28754 19806
rect 28702 19730 28754 19742
rect 29038 19794 29090 19806
rect 47854 19794 47906 19806
rect 34066 19742 34078 19794
rect 34130 19742 34142 19794
rect 47394 19742 47406 19794
rect 47458 19742 47470 19794
rect 29038 19730 29090 19742
rect 47854 19730 47906 19742
rect 52110 19794 52162 19806
rect 52110 19730 52162 19742
rect 52782 19794 52834 19806
rect 52782 19730 52834 19742
rect 53118 19794 53170 19806
rect 53118 19730 53170 19742
rect 57486 19794 57538 19806
rect 57486 19730 57538 19742
rect 1344 19626 62608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 62608 19626
rect 1344 19540 62608 19574
rect 21422 19458 21474 19470
rect 21422 19394 21474 19406
rect 21758 19458 21810 19470
rect 21758 19394 21810 19406
rect 26686 19458 26738 19470
rect 26686 19394 26738 19406
rect 42030 19458 42082 19470
rect 52782 19458 52834 19470
rect 59838 19458 59890 19470
rect 45042 19406 45054 19458
rect 45106 19406 45118 19458
rect 56802 19406 56814 19458
rect 56866 19406 56878 19458
rect 60498 19406 60510 19458
rect 60562 19406 60574 19458
rect 42030 19394 42082 19406
rect 52782 19394 52834 19406
rect 59838 19394 59890 19406
rect 19518 19346 19570 19358
rect 5954 19294 5966 19346
rect 6018 19294 6030 19346
rect 14130 19294 14142 19346
rect 14194 19294 14206 19346
rect 16930 19294 16942 19346
rect 16994 19294 17006 19346
rect 19518 19282 19570 19294
rect 23214 19346 23266 19358
rect 23214 19282 23266 19294
rect 29374 19346 29426 19358
rect 29374 19282 29426 19294
rect 30158 19346 30210 19358
rect 51662 19346 51714 19358
rect 36194 19294 36206 19346
rect 36258 19294 36270 19346
rect 42242 19294 42254 19346
rect 42306 19294 42318 19346
rect 47170 19294 47182 19346
rect 47234 19294 47246 19346
rect 50530 19294 50542 19346
rect 50594 19294 50606 19346
rect 53218 19294 53230 19346
rect 53282 19294 53294 19346
rect 30158 19282 30210 19294
rect 51662 19282 51714 19294
rect 6414 19234 6466 19246
rect 4722 19182 4734 19234
rect 4786 19182 4798 19234
rect 6414 19170 6466 19182
rect 6638 19234 6690 19246
rect 6638 19170 6690 19182
rect 6974 19234 7026 19246
rect 7758 19234 7810 19246
rect 9886 19234 9938 19246
rect 15710 19234 15762 19246
rect 19630 19234 19682 19246
rect 26686 19234 26738 19246
rect 7298 19182 7310 19234
rect 7362 19182 7374 19234
rect 9650 19182 9662 19234
rect 9714 19182 9726 19234
rect 10322 19182 10334 19234
rect 10386 19182 10398 19234
rect 11778 19182 11790 19234
rect 11842 19182 11854 19234
rect 12338 19182 12350 19234
rect 12402 19182 12414 19234
rect 13906 19182 13918 19234
rect 13970 19182 13982 19234
rect 14578 19182 14590 19234
rect 14642 19182 14654 19234
rect 16818 19182 16830 19234
rect 16882 19182 16894 19234
rect 20402 19182 20414 19234
rect 20466 19182 20478 19234
rect 24210 19182 24222 19234
rect 24274 19182 24286 19234
rect 25554 19182 25566 19234
rect 25618 19182 25630 19234
rect 6974 19170 7026 19182
rect 7758 19170 7810 19182
rect 9886 19170 9938 19182
rect 15710 19170 15762 19182
rect 19630 19170 19682 19182
rect 26686 19170 26738 19182
rect 27022 19234 27074 19246
rect 29598 19234 29650 19246
rect 34190 19234 34242 19246
rect 35758 19234 35810 19246
rect 43038 19234 43090 19246
rect 27122 19182 27134 19234
rect 27186 19182 27198 19234
rect 33058 19182 33070 19234
rect 33122 19182 33134 19234
rect 34962 19182 34974 19234
rect 35026 19182 35038 19234
rect 36082 19182 36094 19234
rect 36146 19182 36158 19234
rect 42354 19182 42366 19234
rect 42418 19182 42430 19234
rect 27022 19170 27074 19182
rect 29598 19170 29650 19182
rect 34190 19170 34242 19182
rect 35758 19170 35810 19182
rect 43038 19170 43090 19182
rect 44270 19234 44322 19246
rect 45950 19234 46002 19246
rect 51214 19234 51266 19246
rect 44818 19182 44830 19234
rect 44882 19182 44894 19234
rect 46386 19182 46398 19234
rect 46450 19182 46462 19234
rect 47730 19182 47742 19234
rect 47794 19182 47806 19234
rect 44270 19170 44322 19182
rect 45950 19170 46002 19182
rect 51214 19170 51266 19182
rect 52222 19234 52274 19246
rect 56254 19234 56306 19246
rect 52546 19182 52558 19234
rect 52610 19182 52622 19234
rect 53554 19182 53566 19234
rect 53618 19182 53630 19234
rect 54338 19182 54350 19234
rect 54402 19182 54414 19234
rect 55682 19182 55694 19234
rect 55746 19182 55758 19234
rect 56466 19182 56478 19234
rect 56530 19182 56542 19234
rect 58146 19182 58158 19234
rect 58210 19182 58222 19234
rect 58482 19182 58494 19234
rect 58546 19182 58558 19234
rect 59490 19182 59502 19234
rect 59554 19182 59566 19234
rect 60722 19182 60734 19234
rect 60786 19182 60798 19234
rect 52222 19170 52274 19182
rect 56254 19170 56306 19182
rect 5630 19122 5682 19134
rect 2930 19070 2942 19122
rect 2994 19070 3006 19122
rect 5630 19058 5682 19070
rect 11118 19122 11170 19134
rect 11118 19058 11170 19070
rect 11454 19122 11506 19134
rect 15374 19122 15426 19134
rect 12562 19070 12574 19122
rect 12626 19070 12638 19122
rect 14242 19070 14254 19122
rect 14306 19070 14318 19122
rect 14914 19070 14926 19122
rect 14978 19070 14990 19122
rect 11454 19058 11506 19070
rect 15374 19058 15426 19070
rect 15486 19122 15538 19134
rect 15486 19058 15538 19070
rect 16494 19122 16546 19134
rect 23774 19122 23826 19134
rect 21970 19070 21982 19122
rect 22034 19070 22046 19122
rect 22306 19070 22318 19122
rect 22370 19070 22382 19122
rect 16494 19058 16546 19070
rect 23774 19058 23826 19070
rect 24558 19122 24610 19134
rect 24558 19058 24610 19070
rect 24670 19122 24722 19134
rect 34750 19122 34802 19134
rect 42702 19122 42754 19134
rect 31154 19070 31166 19122
rect 31218 19070 31230 19122
rect 33282 19070 33294 19122
rect 33346 19070 33358 19122
rect 33842 19070 33854 19122
rect 33906 19070 33918 19122
rect 38546 19070 38558 19122
rect 38610 19070 38622 19122
rect 40226 19070 40238 19122
rect 40290 19070 40302 19122
rect 24670 19058 24722 19070
rect 34750 19058 34802 19070
rect 42702 19058 42754 19070
rect 43710 19122 43762 19134
rect 43710 19058 43762 19070
rect 44046 19122 44098 19134
rect 45502 19122 45554 19134
rect 45378 19070 45390 19122
rect 45442 19070 45454 19122
rect 44046 19058 44098 19070
rect 45502 19058 45554 19070
rect 45614 19122 45666 19134
rect 45614 19058 45666 19070
rect 46846 19122 46898 19134
rect 59726 19122 59778 19134
rect 48402 19070 48414 19122
rect 48466 19070 48478 19122
rect 50866 19070 50878 19122
rect 50930 19070 50942 19122
rect 58594 19070 58606 19122
rect 58658 19070 58670 19122
rect 46846 19058 46898 19070
rect 59726 19058 59778 19070
rect 61406 19122 61458 19134
rect 61842 19070 61854 19122
rect 61906 19070 61918 19122
rect 61406 19058 61458 19070
rect 2046 19010 2098 19022
rect 2046 18946 2098 18958
rect 6750 19010 6802 19022
rect 15934 19010 15986 19022
rect 11890 18958 11902 19010
rect 11954 18958 11966 19010
rect 6750 18946 6802 18958
rect 15934 18946 15986 18958
rect 23662 19010 23714 19022
rect 23662 18946 23714 18958
rect 24782 19010 24834 19022
rect 24782 18946 24834 18958
rect 24894 19010 24946 19022
rect 24894 18946 24946 18958
rect 32510 19010 32562 19022
rect 32510 18946 32562 18958
rect 37102 19010 37154 19022
rect 37102 18946 37154 18958
rect 42814 19010 42866 19022
rect 42814 18946 42866 18958
rect 43934 19010 43986 19022
rect 43934 18946 43986 18958
rect 47070 19010 47122 19022
rect 47070 18946 47122 18958
rect 51550 19010 51602 19022
rect 51550 18946 51602 18958
rect 51774 19010 51826 19022
rect 51774 18946 51826 18958
rect 59838 19010 59890 19022
rect 59838 18946 59890 18958
rect 61518 19010 61570 19022
rect 61518 18946 61570 18958
rect 62190 19010 62242 19022
rect 62190 18946 62242 18958
rect 1344 18842 62608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 62608 18842
rect 1344 18756 62608 18790
rect 8430 18674 8482 18686
rect 8430 18610 8482 18622
rect 10334 18674 10386 18686
rect 10334 18610 10386 18622
rect 13358 18674 13410 18686
rect 13358 18610 13410 18622
rect 13582 18674 13634 18686
rect 13582 18610 13634 18622
rect 24110 18674 24162 18686
rect 24110 18610 24162 18622
rect 24334 18674 24386 18686
rect 36878 18674 36930 18686
rect 33170 18622 33182 18674
rect 33234 18622 33246 18674
rect 24334 18610 24386 18622
rect 36878 18610 36930 18622
rect 41022 18674 41074 18686
rect 41022 18610 41074 18622
rect 50206 18674 50258 18686
rect 50206 18610 50258 18622
rect 53790 18674 53842 18686
rect 60846 18674 60898 18686
rect 57698 18622 57710 18674
rect 57762 18622 57774 18674
rect 53790 18610 53842 18622
rect 60846 18610 60898 18622
rect 8654 18562 8706 18574
rect 4834 18510 4846 18562
rect 4898 18510 4910 18562
rect 8654 18498 8706 18510
rect 10558 18562 10610 18574
rect 22430 18562 22482 18574
rect 35758 18562 35810 18574
rect 49422 18562 49474 18574
rect 11330 18510 11342 18562
rect 11394 18510 11406 18562
rect 13906 18510 13918 18562
rect 13970 18510 13982 18562
rect 16034 18510 16046 18562
rect 16098 18510 16110 18562
rect 16594 18510 16606 18562
rect 16658 18510 16670 18562
rect 25778 18510 25790 18562
rect 25842 18510 25854 18562
rect 33730 18510 33742 18562
rect 33794 18510 33806 18562
rect 42018 18510 42030 18562
rect 42082 18510 42094 18562
rect 44930 18510 44942 18562
rect 44994 18510 45006 18562
rect 46050 18510 46062 18562
rect 46114 18510 46126 18562
rect 10558 18498 10610 18510
rect 22430 18498 22482 18510
rect 35758 18498 35810 18510
rect 49422 18498 49474 18510
rect 49534 18562 49586 18574
rect 51326 18562 51378 18574
rect 50978 18510 50990 18562
rect 51042 18510 51054 18562
rect 49534 18498 49586 18510
rect 51326 18498 51378 18510
rect 53678 18562 53730 18574
rect 53678 18498 53730 18510
rect 54014 18562 54066 18574
rect 61854 18562 61906 18574
rect 57026 18510 57038 18562
rect 57090 18510 57102 18562
rect 59938 18510 59950 18562
rect 60002 18510 60014 18562
rect 54014 18498 54066 18510
rect 61854 18498 61906 18510
rect 2718 18450 2770 18462
rect 2718 18386 2770 18398
rect 3054 18450 3106 18462
rect 3054 18386 3106 18398
rect 3614 18450 3666 18462
rect 7534 18450 7586 18462
rect 13470 18450 13522 18462
rect 16718 18450 16770 18462
rect 6514 18398 6526 18450
rect 6578 18398 6590 18450
rect 7858 18398 7870 18450
rect 7922 18398 7934 18450
rect 8194 18398 8206 18450
rect 8258 18398 8270 18450
rect 9986 18398 9998 18450
rect 10050 18398 10062 18450
rect 13794 18398 13806 18450
rect 13858 18398 13870 18450
rect 15362 18398 15374 18450
rect 15426 18398 15438 18450
rect 3614 18386 3666 18398
rect 7534 18386 7586 18398
rect 13470 18386 13522 18398
rect 16718 18386 16770 18398
rect 18062 18450 18114 18462
rect 19854 18450 19906 18462
rect 18946 18398 18958 18450
rect 19010 18398 19022 18450
rect 18062 18386 18114 18398
rect 19854 18386 19906 18398
rect 20190 18450 20242 18462
rect 22766 18450 22818 18462
rect 20514 18398 20526 18450
rect 20578 18398 20590 18450
rect 22194 18398 22206 18450
rect 22258 18398 22270 18450
rect 20190 18386 20242 18398
rect 22766 18386 22818 18398
rect 24222 18450 24274 18462
rect 28254 18450 28306 18462
rect 24658 18398 24670 18450
rect 24722 18398 24734 18450
rect 24222 18386 24274 18398
rect 28254 18386 28306 18398
rect 28366 18450 28418 18462
rect 28366 18386 28418 18398
rect 30494 18450 30546 18462
rect 42702 18450 42754 18462
rect 30706 18398 30718 18450
rect 30770 18398 30782 18450
rect 32386 18398 32398 18450
rect 32450 18398 32462 18450
rect 33058 18398 33070 18450
rect 33122 18398 33134 18450
rect 33618 18398 33630 18450
rect 33682 18398 33694 18450
rect 35074 18398 35086 18450
rect 35138 18398 35150 18450
rect 36194 18398 36206 18450
rect 36258 18398 36270 18450
rect 37426 18398 37438 18450
rect 37490 18398 37502 18450
rect 42130 18398 42142 18450
rect 42194 18398 42206 18450
rect 30494 18386 30546 18398
rect 42702 18386 42754 18398
rect 42814 18450 42866 18462
rect 42814 18386 42866 18398
rect 43150 18450 43202 18462
rect 43150 18386 43202 18398
rect 44046 18450 44098 18462
rect 49758 18450 49810 18462
rect 45154 18398 45166 18450
rect 45218 18398 45230 18450
rect 46274 18398 46286 18450
rect 46338 18398 46350 18450
rect 47618 18398 47630 18450
rect 47682 18398 47694 18450
rect 48738 18398 48750 18450
rect 48802 18398 48814 18450
rect 44046 18386 44098 18398
rect 49758 18386 49810 18398
rect 49982 18450 50034 18462
rect 49982 18386 50034 18398
rect 50654 18450 50706 18462
rect 52334 18450 52386 18462
rect 53342 18450 53394 18462
rect 51986 18398 51998 18450
rect 52050 18398 52062 18450
rect 53106 18398 53118 18450
rect 53170 18398 53182 18450
rect 50654 18386 50706 18398
rect 52334 18386 52386 18398
rect 53342 18386 53394 18398
rect 54126 18450 54178 18462
rect 54126 18386 54178 18398
rect 54910 18450 54962 18462
rect 54910 18386 54962 18398
rect 56030 18450 56082 18462
rect 61182 18450 61234 18462
rect 57362 18398 57374 18450
rect 57426 18398 57438 18450
rect 57922 18398 57934 18450
rect 57986 18398 57998 18450
rect 62066 18398 62078 18450
rect 62130 18398 62142 18450
rect 56030 18386 56082 18398
rect 61182 18386 61234 18398
rect 2270 18338 2322 18350
rect 2270 18274 2322 18286
rect 3950 18338 4002 18350
rect 9774 18338 9826 18350
rect 8306 18286 8318 18338
rect 8370 18286 8382 18338
rect 3950 18274 4002 18286
rect 9774 18274 9826 18286
rect 10446 18338 10498 18350
rect 16942 18338 16994 18350
rect 23326 18338 23378 18350
rect 15026 18286 15038 18338
rect 15090 18286 15102 18338
rect 17602 18286 17614 18338
rect 17666 18286 17678 18338
rect 10446 18274 10498 18286
rect 16942 18274 16994 18286
rect 23326 18274 23378 18286
rect 23886 18338 23938 18350
rect 23886 18274 23938 18286
rect 27022 18338 27074 18350
rect 27022 18274 27074 18286
rect 28702 18338 28754 18350
rect 28702 18274 28754 18286
rect 31950 18338 32002 18350
rect 43038 18338 43090 18350
rect 35410 18286 35422 18338
rect 35474 18286 35486 18338
rect 38210 18286 38222 18338
rect 38274 18286 38286 18338
rect 40338 18286 40350 18338
rect 40402 18286 40414 18338
rect 31950 18274 32002 18286
rect 43038 18274 43090 18286
rect 43598 18338 43650 18350
rect 50094 18338 50146 18350
rect 46386 18286 46398 18338
rect 46450 18286 46462 18338
rect 48850 18286 48862 18338
rect 48914 18286 48926 18338
rect 43598 18274 43650 18286
rect 50094 18274 50146 18286
rect 13134 18226 13186 18238
rect 41358 18226 41410 18238
rect 18498 18174 18510 18226
rect 18562 18174 18574 18226
rect 35074 18174 35086 18226
rect 35138 18174 35150 18226
rect 13134 18162 13186 18174
rect 41358 18162 41410 18174
rect 44382 18226 44434 18238
rect 54350 18226 54402 18238
rect 58494 18226 58546 18238
rect 52210 18174 52222 18226
rect 52274 18174 52286 18226
rect 55794 18174 55806 18226
rect 55858 18174 55870 18226
rect 44382 18162 44434 18174
rect 54350 18162 54402 18174
rect 58494 18162 58546 18174
rect 1344 18058 62608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 62608 18058
rect 1344 17972 62608 18006
rect 12014 17890 12066 17902
rect 12014 17826 12066 17838
rect 14702 17890 14754 17902
rect 14702 17826 14754 17838
rect 15262 17890 15314 17902
rect 15262 17826 15314 17838
rect 15822 17890 15874 17902
rect 25678 17890 25730 17902
rect 39566 17890 39618 17902
rect 18722 17838 18734 17890
rect 18786 17838 18798 17890
rect 33954 17838 33966 17890
rect 34018 17838 34030 17890
rect 15822 17826 15874 17838
rect 25678 17826 25730 17838
rect 39566 17826 39618 17838
rect 40014 17890 40066 17902
rect 40014 17826 40066 17838
rect 41470 17890 41522 17902
rect 41470 17826 41522 17838
rect 44830 17890 44882 17902
rect 44830 17826 44882 17838
rect 45278 17890 45330 17902
rect 45278 17826 45330 17838
rect 51774 17890 51826 17902
rect 60622 17890 60674 17902
rect 55794 17838 55806 17890
rect 55858 17838 55870 17890
rect 51774 17826 51826 17838
rect 60622 17826 60674 17838
rect 2046 17778 2098 17790
rect 2046 17714 2098 17726
rect 5966 17778 6018 17790
rect 5966 17714 6018 17726
rect 6862 17778 6914 17790
rect 6862 17714 6914 17726
rect 11342 17778 11394 17790
rect 11342 17714 11394 17726
rect 14366 17778 14418 17790
rect 35758 17778 35810 17790
rect 19618 17726 19630 17778
rect 19682 17726 19694 17778
rect 20066 17726 20078 17778
rect 20130 17726 20142 17778
rect 24882 17726 24894 17778
rect 24946 17726 24958 17778
rect 29586 17726 29598 17778
rect 29650 17726 29662 17778
rect 30370 17726 30382 17778
rect 30434 17726 30446 17778
rect 30706 17726 30718 17778
rect 30770 17726 30782 17778
rect 14366 17714 14418 17726
rect 35758 17714 35810 17726
rect 37886 17778 37938 17790
rect 37886 17714 37938 17726
rect 44942 17778 44994 17790
rect 44942 17714 44994 17726
rect 48302 17778 48354 17790
rect 52558 17778 52610 17790
rect 50306 17726 50318 17778
rect 50370 17726 50382 17778
rect 48302 17714 48354 17726
rect 52558 17714 52610 17726
rect 56814 17778 56866 17790
rect 56814 17714 56866 17726
rect 7982 17666 8034 17678
rect 9886 17666 9938 17678
rect 19070 17666 19122 17678
rect 26686 17666 26738 17678
rect 29150 17666 29202 17678
rect 34974 17666 35026 17678
rect 7298 17614 7310 17666
rect 7362 17614 7374 17666
rect 9650 17614 9662 17666
rect 9714 17614 9726 17666
rect 10098 17614 10110 17666
rect 10162 17614 10174 17666
rect 12674 17614 12686 17666
rect 12738 17614 12750 17666
rect 18162 17614 18174 17666
rect 18226 17614 18238 17666
rect 19282 17614 19294 17666
rect 19346 17614 19358 17666
rect 20178 17614 20190 17666
rect 20242 17614 20254 17666
rect 21970 17614 21982 17666
rect 22034 17614 22046 17666
rect 26338 17614 26350 17666
rect 26402 17614 26414 17666
rect 27122 17614 27134 17666
rect 27186 17614 27198 17666
rect 28466 17614 28478 17666
rect 28530 17614 28542 17666
rect 30258 17614 30270 17666
rect 30322 17614 30334 17666
rect 30818 17614 30830 17666
rect 30882 17614 30894 17666
rect 7982 17602 8034 17614
rect 9886 17602 9938 17614
rect 19070 17602 19122 17614
rect 26686 17602 26738 17614
rect 29150 17602 29202 17614
rect 34974 17602 35026 17614
rect 36990 17666 37042 17678
rect 36990 17602 37042 17614
rect 37550 17666 37602 17678
rect 37550 17602 37602 17614
rect 38222 17666 38274 17678
rect 38222 17602 38274 17614
rect 40238 17666 40290 17678
rect 40238 17602 40290 17614
rect 41134 17666 41186 17678
rect 41134 17602 41186 17614
rect 41358 17666 41410 17678
rect 41358 17602 41410 17614
rect 42814 17666 42866 17678
rect 42814 17602 42866 17614
rect 43822 17666 43874 17678
rect 48190 17666 48242 17678
rect 47842 17614 47854 17666
rect 47906 17614 47918 17666
rect 43822 17602 43874 17614
rect 48190 17602 48242 17614
rect 49086 17666 49138 17678
rect 54238 17666 54290 17678
rect 61630 17666 61682 17678
rect 49410 17614 49422 17666
rect 49474 17614 49486 17666
rect 50642 17614 50654 17666
rect 50706 17614 50718 17666
rect 51650 17614 51662 17666
rect 51714 17614 51726 17666
rect 51874 17614 51886 17666
rect 51938 17614 51950 17666
rect 53778 17614 53790 17666
rect 53842 17614 53854 17666
rect 54674 17614 54686 17666
rect 54738 17614 54750 17666
rect 55010 17614 55022 17666
rect 55074 17614 55086 17666
rect 56354 17614 56366 17666
rect 56418 17614 56430 17666
rect 57026 17614 57038 17666
rect 57090 17614 57102 17666
rect 60498 17614 60510 17666
rect 60562 17614 60574 17666
rect 60722 17614 60734 17666
rect 60786 17614 60798 17666
rect 49086 17602 49138 17614
rect 54238 17602 54290 17614
rect 61630 17602 61682 17614
rect 61854 17666 61906 17678
rect 61854 17602 61906 17614
rect 62190 17666 62242 17678
rect 62190 17602 62242 17614
rect 15262 17554 15314 17566
rect 3826 17502 3838 17554
rect 3890 17502 3902 17554
rect 12786 17502 12798 17554
rect 12850 17502 12862 17554
rect 13570 17502 13582 17554
rect 13634 17502 13646 17554
rect 14130 17502 14142 17554
rect 14194 17502 14206 17554
rect 15262 17490 15314 17502
rect 15374 17554 15426 17566
rect 21310 17554 21362 17566
rect 17042 17502 17054 17554
rect 17106 17502 17118 17554
rect 15374 17490 15426 17502
rect 21310 17490 21362 17502
rect 21646 17554 21698 17566
rect 36094 17554 36146 17566
rect 22754 17502 22766 17554
rect 22818 17502 22830 17554
rect 32386 17502 32398 17554
rect 32450 17502 32462 17554
rect 21646 17490 21698 17502
rect 36094 17490 36146 17502
rect 38446 17554 38498 17566
rect 38446 17490 38498 17502
rect 39454 17554 39506 17566
rect 39454 17490 39506 17502
rect 39678 17554 39730 17566
rect 39678 17490 39730 17502
rect 40798 17554 40850 17566
rect 40798 17490 40850 17502
rect 40910 17554 40962 17566
rect 43710 17554 43762 17566
rect 48414 17554 48466 17566
rect 52110 17554 52162 17566
rect 54462 17554 54514 17566
rect 42242 17502 42254 17554
rect 42306 17502 42318 17554
rect 42578 17502 42590 17554
rect 42642 17502 42654 17554
rect 47170 17502 47182 17554
rect 47234 17502 47246 17554
rect 49522 17502 49534 17554
rect 49586 17502 49598 17554
rect 53218 17502 53230 17554
rect 53282 17502 53294 17554
rect 53666 17502 53678 17554
rect 53730 17502 53742 17554
rect 40910 17490 40962 17502
rect 43710 17490 43762 17502
rect 48414 17490 48466 17502
rect 52110 17490 52162 17502
rect 54462 17490 54514 17502
rect 55358 17554 55410 17566
rect 60958 17554 61010 17566
rect 59378 17502 59390 17554
rect 59442 17502 59454 17554
rect 61282 17502 61294 17554
rect 61346 17502 61358 17554
rect 55358 17490 55410 17502
rect 60958 17490 61010 17502
rect 2494 17442 2546 17454
rect 2494 17378 2546 17390
rect 2830 17442 2882 17454
rect 2830 17378 2882 17390
rect 4958 17442 5010 17454
rect 4958 17378 5010 17390
rect 5854 17442 5906 17454
rect 5854 17378 5906 17390
rect 6302 17442 6354 17454
rect 6302 17378 6354 17390
rect 11678 17442 11730 17454
rect 11678 17378 11730 17390
rect 35086 17442 35138 17454
rect 35086 17378 35138 17390
rect 35310 17442 35362 17454
rect 35310 17378 35362 17390
rect 35646 17442 35698 17454
rect 35646 17378 35698 17390
rect 35870 17442 35922 17454
rect 35870 17378 35922 17390
rect 38894 17442 38946 17454
rect 38894 17378 38946 17390
rect 41470 17442 41522 17454
rect 41470 17378 41522 17390
rect 43150 17442 43202 17454
rect 43150 17378 43202 17390
rect 43598 17442 43650 17454
rect 43598 17378 43650 17390
rect 44046 17442 44098 17454
rect 44046 17378 44098 17390
rect 48862 17442 48914 17454
rect 48862 17378 48914 17390
rect 48974 17442 49026 17454
rect 54350 17442 54402 17454
rect 49970 17390 49982 17442
rect 50034 17390 50046 17442
rect 48974 17378 49026 17390
rect 54350 17378 54402 17390
rect 57934 17442 57986 17454
rect 57934 17378 57986 17390
rect 62078 17442 62130 17454
rect 62078 17378 62130 17390
rect 1344 17274 62608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 62608 17274
rect 1344 17188 62608 17222
rect 2606 17106 2658 17118
rect 2606 17042 2658 17054
rect 2942 17106 2994 17118
rect 2942 17042 2994 17054
rect 3950 17106 4002 17118
rect 3950 17042 4002 17054
rect 4398 17106 4450 17118
rect 4398 17042 4450 17054
rect 5630 17106 5682 17118
rect 5630 17042 5682 17054
rect 5854 17106 5906 17118
rect 5854 17042 5906 17054
rect 8878 17106 8930 17118
rect 13918 17106 13970 17118
rect 10994 17054 11006 17106
rect 11058 17054 11070 17106
rect 8878 17042 8930 17054
rect 13918 17042 13970 17054
rect 15486 17106 15538 17118
rect 15486 17042 15538 17054
rect 16606 17106 16658 17118
rect 16606 17042 16658 17054
rect 17614 17106 17666 17118
rect 17614 17042 17666 17054
rect 18734 17106 18786 17118
rect 18734 17042 18786 17054
rect 18958 17106 19010 17118
rect 18958 17042 19010 17054
rect 24334 17106 24386 17118
rect 24334 17042 24386 17054
rect 24558 17106 24610 17118
rect 24558 17042 24610 17054
rect 26014 17106 26066 17118
rect 33854 17106 33906 17118
rect 30370 17054 30382 17106
rect 30434 17054 30446 17106
rect 26014 17042 26066 17054
rect 33854 17042 33906 17054
rect 34078 17106 34130 17118
rect 34078 17042 34130 17054
rect 36766 17106 36818 17118
rect 36766 17042 36818 17054
rect 40350 17106 40402 17118
rect 40350 17042 40402 17054
rect 46174 17106 46226 17118
rect 53790 17106 53842 17118
rect 47058 17054 47070 17106
rect 47122 17054 47134 17106
rect 49298 17054 49310 17106
rect 49362 17054 49374 17106
rect 46174 17042 46226 17054
rect 53790 17042 53842 17054
rect 54574 17106 54626 17118
rect 54574 17042 54626 17054
rect 56030 17106 56082 17118
rect 60846 17106 60898 17118
rect 56578 17054 56590 17106
rect 56642 17054 56654 17106
rect 60498 17054 60510 17106
rect 60562 17054 60574 17106
rect 56030 17042 56082 17054
rect 60846 17042 60898 17054
rect 61182 17106 61234 17118
rect 62190 17106 62242 17118
rect 61506 17054 61518 17106
rect 61570 17054 61582 17106
rect 61182 17042 61234 17054
rect 62190 17042 62242 17054
rect 4846 16994 4898 17006
rect 4846 16930 4898 16942
rect 5070 16994 5122 17006
rect 6974 16994 7026 17006
rect 16270 16994 16322 17006
rect 6402 16942 6414 16994
rect 6466 16942 6478 16994
rect 7970 16942 7982 16994
rect 8034 16942 8046 16994
rect 8306 16942 8318 16994
rect 8370 16942 8382 16994
rect 14466 16942 14478 16994
rect 14530 16942 14542 16994
rect 14914 16942 14926 16994
rect 14978 16942 14990 16994
rect 5070 16930 5122 16942
rect 6974 16930 7026 16942
rect 16270 16930 16322 16942
rect 16718 16994 16770 17006
rect 16718 16930 16770 16942
rect 17950 16994 18002 17006
rect 17950 16930 18002 16942
rect 19070 16994 19122 17006
rect 23886 16994 23938 17006
rect 20402 16942 20414 16994
rect 20466 16942 20478 16994
rect 19070 16930 19122 16942
rect 23886 16930 23938 16942
rect 24670 16994 24722 17006
rect 25790 16994 25842 17006
rect 31614 16994 31666 17006
rect 25442 16942 25454 16994
rect 25506 16942 25518 16994
rect 26674 16942 26686 16994
rect 26738 16942 26750 16994
rect 27010 16942 27022 16994
rect 27074 16942 27086 16994
rect 28130 16942 28142 16994
rect 28194 16942 28206 16994
rect 24670 16930 24722 16942
rect 25790 16930 25842 16942
rect 31614 16930 31666 16942
rect 32062 16994 32114 17006
rect 32062 16930 32114 16942
rect 32174 16994 32226 17006
rect 34750 16994 34802 17006
rect 38894 16994 38946 17006
rect 33506 16942 33518 16994
rect 33570 16942 33582 16994
rect 37202 16942 37214 16994
rect 37266 16942 37278 16994
rect 32174 16930 32226 16942
rect 34750 16930 34802 16942
rect 38894 16930 38946 16942
rect 39006 16994 39058 17006
rect 39006 16930 39058 16942
rect 41358 16994 41410 17006
rect 41358 16930 41410 16942
rect 41918 16994 41970 17006
rect 46510 16994 46562 17006
rect 43250 16942 43262 16994
rect 43314 16942 43326 16994
rect 41918 16930 41970 16942
rect 46510 16930 46562 16942
rect 47406 16994 47458 17006
rect 47406 16930 47458 16942
rect 54798 16994 54850 17006
rect 55806 16994 55858 17006
rect 55458 16942 55470 16994
rect 55522 16942 55534 16994
rect 54798 16930 54850 16942
rect 55806 16930 55858 16942
rect 55918 16994 55970 17006
rect 55918 16930 55970 16942
rect 57598 16994 57650 17006
rect 57598 16930 57650 16942
rect 57710 16994 57762 17006
rect 59378 16942 59390 16994
rect 59442 16942 59454 16994
rect 61842 16942 61854 16994
rect 61906 16942 61918 16994
rect 57710 16930 57762 16942
rect 5182 16882 5234 16894
rect 5182 16818 5234 16830
rect 5518 16882 5570 16894
rect 6862 16882 6914 16894
rect 6178 16830 6190 16882
rect 6242 16830 6254 16882
rect 5518 16818 5570 16830
rect 6862 16818 6914 16830
rect 7422 16882 7474 16894
rect 7422 16818 7474 16830
rect 10110 16882 10162 16894
rect 10110 16818 10162 16830
rect 12910 16882 12962 16894
rect 12910 16818 12962 16830
rect 14254 16882 14306 16894
rect 15934 16882 15986 16894
rect 15474 16830 15486 16882
rect 15538 16830 15550 16882
rect 14254 16818 14306 16830
rect 15934 16818 15986 16830
rect 18174 16882 18226 16894
rect 18174 16818 18226 16830
rect 18398 16882 18450 16894
rect 24110 16882 24162 16894
rect 27246 16882 27298 16894
rect 19506 16830 19518 16882
rect 19570 16830 19582 16882
rect 20514 16830 20526 16882
rect 20578 16830 20590 16882
rect 21970 16830 21982 16882
rect 22034 16830 22046 16882
rect 23538 16830 23550 16882
rect 23602 16830 23614 16882
rect 25554 16830 25566 16882
rect 25618 16830 25630 16882
rect 18398 16818 18450 16830
rect 24110 16818 24162 16830
rect 27246 16818 27298 16830
rect 27582 16882 27634 16894
rect 29934 16882 29986 16894
rect 31278 16882 31330 16894
rect 34526 16882 34578 16894
rect 29026 16830 29038 16882
rect 29090 16830 29102 16882
rect 30930 16830 30942 16882
rect 30994 16830 31006 16882
rect 33282 16830 33294 16882
rect 33346 16830 33358 16882
rect 27582 16818 27634 16830
rect 29934 16818 29986 16830
rect 31278 16818 31330 16830
rect 34526 16818 34578 16830
rect 34974 16882 35026 16894
rect 34974 16818 35026 16830
rect 35310 16882 35362 16894
rect 35310 16818 35362 16830
rect 35534 16882 35586 16894
rect 35534 16818 35586 16830
rect 35870 16882 35922 16894
rect 35870 16818 35922 16830
rect 36094 16882 36146 16894
rect 36094 16818 36146 16830
rect 37550 16882 37602 16894
rect 37550 16818 37602 16830
rect 37886 16882 37938 16894
rect 37886 16818 37938 16830
rect 39230 16882 39282 16894
rect 39230 16818 39282 16830
rect 39678 16882 39730 16894
rect 39678 16818 39730 16830
rect 39902 16882 39954 16894
rect 39902 16818 39954 16830
rect 41134 16882 41186 16894
rect 41134 16818 41186 16830
rect 41470 16882 41522 16894
rect 41470 16818 41522 16830
rect 41806 16882 41858 16894
rect 41806 16818 41858 16830
rect 42142 16882 42194 16894
rect 47966 16882 48018 16894
rect 42578 16830 42590 16882
rect 42642 16830 42654 16882
rect 44258 16830 44270 16882
rect 44322 16830 44334 16882
rect 45714 16830 45726 16882
rect 45778 16830 45790 16882
rect 47618 16830 47630 16882
rect 47682 16830 47694 16882
rect 42142 16818 42194 16830
rect 47966 16818 48018 16830
rect 48750 16882 48802 16894
rect 48750 16818 48802 16830
rect 49758 16882 49810 16894
rect 54350 16882 54402 16894
rect 57374 16882 57426 16894
rect 50194 16830 50206 16882
rect 50258 16830 50270 16882
rect 53666 16830 53678 16882
rect 53730 16830 53742 16882
rect 55570 16830 55582 16882
rect 55634 16830 55646 16882
rect 57138 16830 57150 16882
rect 57202 16830 57214 16882
rect 49758 16818 49810 16830
rect 54350 16818 54402 16830
rect 57374 16818 57426 16830
rect 2158 16770 2210 16782
rect 2158 16706 2210 16718
rect 3502 16770 3554 16782
rect 3502 16706 3554 16718
rect 7198 16770 7250 16782
rect 7198 16706 7250 16718
rect 8542 16770 8594 16782
rect 8542 16706 8594 16718
rect 18286 16770 18338 16782
rect 23998 16770 24050 16782
rect 33966 16770 34018 16782
rect 19058 16718 19070 16770
rect 19122 16718 19134 16770
rect 21858 16718 21870 16770
rect 21922 16718 21934 16770
rect 25666 16718 25678 16770
rect 25730 16718 25742 16770
rect 18286 16706 18338 16718
rect 23998 16706 24050 16718
rect 33966 16706 34018 16718
rect 34862 16770 34914 16782
rect 34862 16706 34914 16718
rect 35758 16770 35810 16782
rect 35758 16706 35810 16718
rect 39790 16770 39842 16782
rect 39790 16706 39842 16718
rect 46734 16770 46786 16782
rect 54462 16770 54514 16782
rect 50866 16718 50878 16770
rect 50930 16718 50942 16770
rect 52994 16718 53006 16770
rect 53058 16718 53070 16770
rect 46734 16706 46786 16718
rect 54462 16706 54514 16718
rect 15822 16658 15874 16670
rect 2146 16606 2158 16658
rect 2210 16655 2222 16658
rect 3266 16655 3278 16658
rect 2210 16609 3278 16655
rect 2210 16606 2222 16609
rect 3266 16606 3278 16609
rect 3330 16606 3342 16658
rect 15822 16594 15874 16606
rect 20302 16658 20354 16670
rect 29710 16658 29762 16670
rect 28242 16606 28254 16658
rect 28306 16606 28318 16658
rect 20302 16594 20354 16606
rect 29710 16594 29762 16606
rect 32062 16658 32114 16670
rect 32062 16594 32114 16606
rect 38110 16658 38162 16670
rect 38894 16658 38946 16670
rect 47294 16658 47346 16670
rect 38434 16606 38446 16658
rect 38498 16606 38510 16658
rect 42914 16606 42926 16658
rect 42978 16606 42990 16658
rect 38110 16594 38162 16606
rect 38894 16594 38946 16606
rect 47294 16594 47346 16606
rect 48974 16658 49026 16670
rect 48974 16594 49026 16606
rect 58158 16658 58210 16670
rect 58158 16594 58210 16606
rect 1344 16490 62608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 62608 16490
rect 1344 16404 62608 16438
rect 12126 16322 12178 16334
rect 10210 16270 10222 16322
rect 10274 16270 10286 16322
rect 12126 16258 12178 16270
rect 12350 16322 12402 16334
rect 12350 16258 12402 16270
rect 12910 16322 12962 16334
rect 12910 16258 12962 16270
rect 13918 16322 13970 16334
rect 13918 16258 13970 16270
rect 15374 16322 15426 16334
rect 15374 16258 15426 16270
rect 30270 16322 30322 16334
rect 49086 16322 49138 16334
rect 45042 16270 45054 16322
rect 45106 16270 45118 16322
rect 30270 16258 30322 16270
rect 49086 16258 49138 16270
rect 50206 16322 50258 16334
rect 55458 16270 55470 16322
rect 55522 16270 55534 16322
rect 50206 16258 50258 16270
rect 2270 16210 2322 16222
rect 2270 16146 2322 16158
rect 3166 16210 3218 16222
rect 3166 16146 3218 16158
rect 3614 16210 3666 16222
rect 13582 16210 13634 16222
rect 26686 16210 26738 16222
rect 6626 16158 6638 16210
rect 6690 16158 6702 16210
rect 10658 16158 10670 16210
rect 10722 16158 10734 16210
rect 20626 16158 20638 16210
rect 20690 16158 20702 16210
rect 3614 16146 3666 16158
rect 13582 16146 13634 16158
rect 26686 16146 26738 16158
rect 30718 16210 30770 16222
rect 49870 16210 49922 16222
rect 36418 16158 36430 16210
rect 36482 16158 36494 16210
rect 39330 16158 39342 16210
rect 39394 16158 39406 16210
rect 41458 16158 41470 16210
rect 41522 16158 41534 16210
rect 41906 16158 41918 16210
rect 41970 16158 41982 16210
rect 47394 16158 47406 16210
rect 47458 16158 47470 16210
rect 49522 16158 49534 16210
rect 49586 16158 49598 16210
rect 30718 16146 30770 16158
rect 49870 16146 49922 16158
rect 50766 16210 50818 16222
rect 50766 16146 50818 16158
rect 51438 16210 51490 16222
rect 51438 16146 51490 16158
rect 51886 16210 51938 16222
rect 58046 16210 58098 16222
rect 54562 16158 54574 16210
rect 54626 16158 54638 16210
rect 51886 16146 51938 16158
rect 58046 16146 58098 16158
rect 58382 16210 58434 16222
rect 60622 16210 60674 16222
rect 59266 16158 59278 16210
rect 59330 16158 59342 16210
rect 58382 16146 58434 16158
rect 60622 16146 60674 16158
rect 61518 16210 61570 16222
rect 61518 16146 61570 16158
rect 61966 16210 62018 16222
rect 61966 16146 62018 16158
rect 4622 16098 4674 16110
rect 3938 16046 3950 16098
rect 4002 16046 4014 16098
rect 4622 16034 4674 16046
rect 4734 16098 4786 16110
rect 4734 16034 4786 16046
rect 5182 16098 5234 16110
rect 12686 16098 12738 16110
rect 6066 16046 6078 16098
rect 6130 16046 6142 16098
rect 7410 16046 7422 16098
rect 7474 16046 7486 16098
rect 8978 16046 8990 16098
rect 9042 16046 9054 16098
rect 9874 16046 9886 16098
rect 9938 16046 9950 16098
rect 11106 16046 11118 16098
rect 11170 16046 11182 16098
rect 5182 16034 5234 16046
rect 12686 16034 12738 16046
rect 13470 16098 13522 16110
rect 13470 16034 13522 16046
rect 14030 16098 14082 16110
rect 14030 16034 14082 16046
rect 14478 16098 14530 16110
rect 14478 16034 14530 16046
rect 14702 16098 14754 16110
rect 14702 16034 14754 16046
rect 15710 16098 15762 16110
rect 15710 16034 15762 16046
rect 15934 16098 15986 16110
rect 26126 16098 26178 16110
rect 18946 16046 18958 16098
rect 19010 16046 19022 16098
rect 20290 16046 20302 16098
rect 20354 16046 20366 16098
rect 21298 16046 21310 16098
rect 21362 16046 21374 16098
rect 23090 16046 23102 16098
rect 23154 16046 23166 16098
rect 15934 16034 15986 16046
rect 26126 16034 26178 16046
rect 28366 16098 28418 16110
rect 28366 16034 28418 16046
rect 28478 16098 28530 16110
rect 28478 16034 28530 16046
rect 29150 16098 29202 16110
rect 29150 16034 29202 16046
rect 29486 16098 29538 16110
rect 29486 16034 29538 16046
rect 29598 16098 29650 16110
rect 31726 16098 31778 16110
rect 29922 16046 29934 16098
rect 29986 16046 29998 16098
rect 31490 16046 31502 16098
rect 31554 16046 31566 16098
rect 29598 16034 29650 16046
rect 31726 16034 31778 16046
rect 32062 16098 32114 16110
rect 32062 16034 32114 16046
rect 32622 16098 32674 16110
rect 32622 16034 32674 16046
rect 32958 16098 33010 16110
rect 42366 16098 42418 16110
rect 33506 16046 33518 16098
rect 33570 16046 33582 16098
rect 37538 16046 37550 16098
rect 37602 16046 37614 16098
rect 38546 16046 38558 16098
rect 38610 16046 38622 16098
rect 32958 16034 33010 16046
rect 42366 16034 42418 16046
rect 43038 16098 43090 16110
rect 43038 16034 43090 16046
rect 43150 16098 43202 16110
rect 43150 16034 43202 16046
rect 44270 16098 44322 16110
rect 45614 16098 45666 16110
rect 48190 16098 48242 16110
rect 44818 16046 44830 16098
rect 44882 16046 44894 16098
rect 46610 16046 46622 16098
rect 46674 16046 46686 16098
rect 47058 16046 47070 16098
rect 47122 16046 47134 16098
rect 44270 16034 44322 16046
rect 45614 16034 45666 16046
rect 48190 16034 48242 16046
rect 49310 16098 49362 16110
rect 49310 16034 49362 16046
rect 50430 16098 50482 16110
rect 55358 16098 55410 16110
rect 54674 16046 54686 16098
rect 54738 16046 54750 16098
rect 56578 16046 56590 16098
rect 56642 16046 56654 16098
rect 57586 16046 57598 16098
rect 57650 16046 57662 16098
rect 58818 16046 58830 16098
rect 58882 16046 58894 16098
rect 59490 16046 59502 16098
rect 59554 16046 59566 16098
rect 50430 16034 50482 16046
rect 55358 16034 55410 16046
rect 9662 15986 9714 15998
rect 4162 15934 4174 15986
rect 4226 15934 4238 15986
rect 6178 15934 6190 15986
rect 6242 15934 6254 15986
rect 9662 15922 9714 15934
rect 12574 15986 12626 15998
rect 12574 15922 12626 15934
rect 16382 15986 16434 15998
rect 27694 15986 27746 15998
rect 17378 15934 17390 15986
rect 17442 15934 17454 15986
rect 21746 15934 21758 15986
rect 21810 15934 21822 15986
rect 23426 15934 23438 15986
rect 23490 15934 23502 15986
rect 27346 15934 27358 15986
rect 27410 15934 27422 15986
rect 16382 15922 16434 15934
rect 27694 15922 27746 15934
rect 28030 15986 28082 15998
rect 28030 15922 28082 15934
rect 29262 15986 29314 15998
rect 29262 15922 29314 15934
rect 30158 15986 30210 15998
rect 30158 15922 30210 15934
rect 30942 15986 30994 15998
rect 30942 15922 30994 15934
rect 33070 15986 33122 15998
rect 37102 15986 37154 15998
rect 34290 15934 34302 15986
rect 34354 15934 34366 15986
rect 33070 15922 33122 15934
rect 37102 15922 37154 15934
rect 37774 15986 37826 15998
rect 37774 15922 37826 15934
rect 38110 15986 38162 15998
rect 38110 15922 38162 15934
rect 42142 15986 42194 15998
rect 42142 15922 42194 15934
rect 42814 15986 42866 15998
rect 47854 15986 47906 15998
rect 45378 15934 45390 15986
rect 45442 15934 45454 15986
rect 42814 15922 42866 15934
rect 47854 15922 47906 15934
rect 48414 15986 48466 15998
rect 48414 15922 48466 15934
rect 49646 15986 49698 15998
rect 49646 15922 49698 15934
rect 50878 15986 50930 15998
rect 50878 15922 50930 15934
rect 53118 15986 53170 15998
rect 53118 15922 53170 15934
rect 2718 15874 2770 15886
rect 2718 15810 2770 15822
rect 4958 15874 5010 15886
rect 4958 15810 5010 15822
rect 14814 15874 14866 15886
rect 14814 15810 14866 15822
rect 16270 15874 16322 15886
rect 16270 15810 16322 15822
rect 24110 15874 24162 15886
rect 26574 15874 26626 15886
rect 25218 15822 25230 15874
rect 25282 15822 25294 15874
rect 24110 15810 24162 15822
rect 26574 15810 26626 15822
rect 26798 15874 26850 15886
rect 26798 15810 26850 15822
rect 28142 15874 28194 15886
rect 28142 15810 28194 15822
rect 33294 15874 33346 15886
rect 33294 15810 33346 15822
rect 36990 15874 37042 15886
rect 36990 15810 37042 15822
rect 38222 15874 38274 15886
rect 38222 15810 38274 15822
rect 44830 15874 44882 15886
rect 48078 15874 48130 15886
rect 46050 15822 46062 15874
rect 46114 15822 46126 15874
rect 44830 15810 44882 15822
rect 48078 15810 48130 15822
rect 50654 15874 50706 15886
rect 50654 15810 50706 15822
rect 52782 15874 52834 15886
rect 52782 15810 52834 15822
rect 61070 15874 61122 15886
rect 61070 15810 61122 15822
rect 1344 15706 62608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 62608 15706
rect 1344 15620 62608 15654
rect 2046 15538 2098 15550
rect 2046 15474 2098 15486
rect 2494 15538 2546 15550
rect 2494 15474 2546 15486
rect 3838 15538 3890 15550
rect 3838 15474 3890 15486
rect 4286 15538 4338 15550
rect 4286 15474 4338 15486
rect 5630 15538 5682 15550
rect 5630 15474 5682 15486
rect 13022 15538 13074 15550
rect 13022 15474 13074 15486
rect 13918 15538 13970 15550
rect 13918 15474 13970 15486
rect 16494 15538 16546 15550
rect 16494 15474 16546 15486
rect 22542 15538 22594 15550
rect 25566 15538 25618 15550
rect 32062 15538 32114 15550
rect 24658 15486 24670 15538
rect 24722 15486 24734 15538
rect 25218 15486 25230 15538
rect 25282 15486 25294 15538
rect 30706 15486 30718 15538
rect 30770 15486 30782 15538
rect 22542 15474 22594 15486
rect 25566 15474 25618 15486
rect 32062 15474 32114 15486
rect 34414 15538 34466 15550
rect 34414 15474 34466 15486
rect 37662 15538 37714 15550
rect 41806 15538 41858 15550
rect 38770 15486 38782 15538
rect 38834 15486 38846 15538
rect 37662 15474 37714 15486
rect 41806 15474 41858 15486
rect 49310 15538 49362 15550
rect 49310 15474 49362 15486
rect 50430 15538 50482 15550
rect 50430 15474 50482 15486
rect 55918 15538 55970 15550
rect 55918 15474 55970 15486
rect 59950 15538 60002 15550
rect 59950 15474 60002 15486
rect 60398 15538 60450 15550
rect 60398 15474 60450 15486
rect 60846 15538 60898 15550
rect 60846 15474 60898 15486
rect 61406 15538 61458 15550
rect 61406 15474 61458 15486
rect 61742 15538 61794 15550
rect 61742 15474 61794 15486
rect 62190 15538 62242 15550
rect 62190 15474 62242 15486
rect 5294 15426 5346 15438
rect 4498 15374 4510 15426
rect 4562 15374 4574 15426
rect 5294 15362 5346 15374
rect 5518 15426 5570 15438
rect 12014 15426 12066 15438
rect 7074 15374 7086 15426
rect 7138 15374 7150 15426
rect 9650 15374 9662 15426
rect 9714 15374 9726 15426
rect 5518 15362 5570 15374
rect 12014 15362 12066 15374
rect 13806 15426 13858 15438
rect 17390 15426 17442 15438
rect 33182 15426 33234 15438
rect 14802 15374 14814 15426
rect 14866 15374 14878 15426
rect 20178 15374 20190 15426
rect 20242 15374 20254 15426
rect 21522 15374 21534 15426
rect 21586 15374 21598 15426
rect 28690 15374 28702 15426
rect 28754 15374 28766 15426
rect 13806 15362 13858 15374
rect 17390 15362 17442 15374
rect 33182 15362 33234 15374
rect 33518 15426 33570 15438
rect 41694 15426 41746 15438
rect 47854 15426 47906 15438
rect 35522 15374 35534 15426
rect 35586 15374 35598 15426
rect 41458 15374 41470 15426
rect 41522 15374 41534 15426
rect 42914 15374 42926 15426
rect 42978 15374 42990 15426
rect 46610 15374 46622 15426
rect 46674 15374 46686 15426
rect 33518 15362 33570 15374
rect 41694 15362 41746 15374
rect 47854 15362 47906 15374
rect 50094 15426 50146 15438
rect 51214 15426 51266 15438
rect 50978 15374 50990 15426
rect 51042 15374 51054 15426
rect 51538 15374 51550 15426
rect 51602 15374 51614 15426
rect 53554 15374 53566 15426
rect 53618 15374 53630 15426
rect 54898 15374 54910 15426
rect 54962 15374 54974 15426
rect 55346 15374 55358 15426
rect 55410 15374 55422 15426
rect 50094 15362 50146 15374
rect 51214 15362 51266 15374
rect 4846 15314 4898 15326
rect 4846 15250 4898 15262
rect 5742 15314 5794 15326
rect 5742 15250 5794 15262
rect 6078 15314 6130 15326
rect 8430 15314 8482 15326
rect 11454 15314 11506 15326
rect 6290 15262 6302 15314
rect 6354 15262 6366 15314
rect 7298 15262 7310 15314
rect 7362 15262 7374 15314
rect 8866 15262 8878 15314
rect 8930 15262 8942 15314
rect 9538 15262 9550 15314
rect 9602 15262 9614 15314
rect 10770 15262 10782 15314
rect 10834 15262 10846 15314
rect 10994 15262 11006 15314
rect 11058 15262 11070 15314
rect 6078 15250 6130 15262
rect 8430 15250 8482 15262
rect 11454 15250 11506 15262
rect 11790 15314 11842 15326
rect 11790 15250 11842 15262
rect 12574 15314 12626 15326
rect 13246 15314 13298 15326
rect 23438 15314 23490 15326
rect 12898 15262 12910 15314
rect 12962 15262 12974 15314
rect 21410 15262 21422 15314
rect 21474 15262 21486 15314
rect 12574 15250 12626 15262
rect 13246 15250 13298 15262
rect 23438 15250 23490 15262
rect 24334 15314 24386 15326
rect 33630 15314 33682 15326
rect 27458 15262 27470 15314
rect 27522 15262 27534 15314
rect 28914 15262 28926 15314
rect 28978 15262 28990 15314
rect 24334 15250 24386 15262
rect 33630 15250 33682 15262
rect 34078 15314 34130 15326
rect 39790 15314 39842 15326
rect 34514 15262 34526 15314
rect 34578 15311 34590 15314
rect 34850 15311 34862 15314
rect 34578 15265 34862 15311
rect 34578 15262 34590 15265
rect 34850 15262 34862 15265
rect 34914 15262 34926 15314
rect 34078 15250 34130 15262
rect 39790 15250 39842 15262
rect 40014 15314 40066 15326
rect 40014 15250 40066 15262
rect 40462 15314 40514 15326
rect 40462 15250 40514 15262
rect 42030 15314 42082 15326
rect 44046 15314 44098 15326
rect 48862 15314 48914 15326
rect 43586 15262 43598 15314
rect 43650 15262 43662 15314
rect 44258 15262 44270 15314
rect 44322 15262 44334 15314
rect 42030 15250 42082 15262
rect 44046 15250 44098 15262
rect 48862 15250 48914 15262
rect 48974 15314 49026 15326
rect 51886 15314 51938 15326
rect 49298 15262 49310 15314
rect 49362 15262 49374 15314
rect 49858 15262 49870 15314
rect 49922 15262 49934 15314
rect 50418 15262 50430 15314
rect 50482 15262 50494 15314
rect 56578 15262 56590 15314
rect 56642 15262 56654 15314
rect 48974 15250 49026 15262
rect 51886 15250 51938 15262
rect 2830 15202 2882 15214
rect 2830 15138 2882 15150
rect 3390 15202 3442 15214
rect 11902 15202 11954 15214
rect 7074 15150 7086 15202
rect 7138 15150 7150 15202
rect 10098 15150 10110 15202
rect 10162 15150 10174 15202
rect 3390 15138 3442 15150
rect 11902 15138 11954 15150
rect 13134 15202 13186 15214
rect 18734 15202 18786 15214
rect 17826 15150 17838 15202
rect 17890 15150 17902 15202
rect 13134 15138 13186 15150
rect 18734 15138 18786 15150
rect 23214 15202 23266 15214
rect 24110 15202 24162 15214
rect 39902 15202 39954 15214
rect 49646 15202 49698 15214
rect 23762 15150 23774 15202
rect 23826 15150 23838 15202
rect 27682 15150 27694 15202
rect 27746 15150 27758 15202
rect 41682 15150 41694 15202
rect 41746 15150 41758 15202
rect 23214 15138 23266 15150
rect 24110 15138 24162 15150
rect 39902 15138 39954 15150
rect 49646 15138 49698 15150
rect 52334 15202 52386 15214
rect 52334 15138 52386 15150
rect 55582 15202 55634 15214
rect 57362 15150 57374 15202
rect 57426 15150 57438 15202
rect 59490 15150 59502 15202
rect 59554 15150 59566 15202
rect 55582 15138 55634 15150
rect 14030 15090 14082 15102
rect 14030 15026 14082 15038
rect 22206 15090 22258 15102
rect 33070 15090 33122 15102
rect 26898 15038 26910 15090
rect 26962 15038 26974 15090
rect 22206 15026 22258 15038
rect 33070 15026 33122 15038
rect 34302 15090 34354 15102
rect 34302 15026 34354 15038
rect 37326 15090 37378 15102
rect 45266 15038 45278 15090
rect 45330 15038 45342 15090
rect 50642 15038 50654 15090
rect 50706 15038 50718 15090
rect 37326 15026 37378 15038
rect 1344 14922 62608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 62608 14922
rect 1344 14836 62608 14870
rect 13582 14754 13634 14766
rect 22654 14754 22706 14766
rect 22418 14702 22430 14754
rect 22482 14702 22494 14754
rect 13582 14690 13634 14702
rect 22654 14690 22706 14702
rect 31166 14754 31218 14766
rect 34526 14754 34578 14766
rect 44942 14754 44994 14766
rect 33394 14702 33406 14754
rect 33458 14702 33470 14754
rect 35522 14702 35534 14754
rect 35586 14702 35598 14754
rect 31166 14690 31218 14702
rect 34526 14690 34578 14702
rect 44942 14690 44994 14702
rect 47182 14754 47234 14766
rect 47182 14690 47234 14702
rect 53118 14754 53170 14766
rect 53118 14690 53170 14702
rect 53454 14754 53506 14766
rect 53890 14702 53902 14754
rect 53954 14702 53966 14754
rect 53454 14690 53506 14702
rect 2494 14642 2546 14654
rect 2494 14578 2546 14590
rect 3838 14642 3890 14654
rect 3838 14578 3890 14590
rect 4286 14642 4338 14654
rect 4286 14578 4338 14590
rect 4958 14642 5010 14654
rect 4958 14578 5010 14590
rect 6302 14642 6354 14654
rect 13694 14642 13746 14654
rect 10882 14590 10894 14642
rect 10946 14590 10958 14642
rect 6302 14578 6354 14590
rect 13694 14578 13746 14590
rect 18622 14642 18674 14654
rect 18622 14578 18674 14590
rect 21870 14642 21922 14654
rect 21870 14578 21922 14590
rect 29262 14642 29314 14654
rect 35982 14642 36034 14654
rect 44270 14642 44322 14654
rect 33282 14590 33294 14642
rect 33346 14590 33358 14642
rect 37090 14590 37102 14642
rect 37154 14590 37166 14642
rect 41234 14590 41246 14642
rect 41298 14590 41310 14642
rect 43362 14590 43374 14642
rect 43426 14590 43438 14642
rect 29262 14578 29314 14590
rect 35982 14578 36034 14590
rect 44270 14578 44322 14590
rect 48190 14642 48242 14654
rect 57598 14642 57650 14654
rect 48402 14590 48414 14642
rect 48466 14590 48478 14642
rect 55794 14590 55806 14642
rect 55858 14590 55870 14642
rect 48190 14578 48242 14590
rect 57598 14578 57650 14590
rect 58718 14642 58770 14654
rect 58718 14578 58770 14590
rect 61070 14642 61122 14654
rect 61070 14578 61122 14590
rect 61630 14642 61682 14654
rect 61630 14578 61682 14590
rect 62190 14642 62242 14654
rect 62190 14578 62242 14590
rect 3278 14530 3330 14542
rect 3278 14466 3330 14478
rect 5966 14530 6018 14542
rect 5966 14466 6018 14478
rect 6190 14530 6242 14542
rect 12238 14530 12290 14542
rect 6850 14478 6862 14530
rect 6914 14478 6926 14530
rect 7074 14478 7086 14530
rect 7138 14478 7150 14530
rect 9426 14478 9438 14530
rect 9490 14478 9502 14530
rect 11218 14478 11230 14530
rect 11282 14478 11294 14530
rect 11778 14478 11790 14530
rect 11842 14478 11854 14530
rect 6190 14466 6242 14478
rect 12238 14466 12290 14478
rect 14926 14530 14978 14542
rect 21310 14530 21362 14542
rect 16258 14478 16270 14530
rect 16322 14478 16334 14530
rect 17938 14478 17950 14530
rect 18002 14478 18014 14530
rect 14926 14466 14978 14478
rect 21310 14466 21362 14478
rect 21646 14530 21698 14542
rect 21646 14466 21698 14478
rect 22094 14530 22146 14542
rect 28142 14530 28194 14542
rect 25218 14478 25230 14530
rect 25282 14478 25294 14530
rect 26114 14478 26126 14530
rect 26178 14478 26190 14530
rect 26562 14478 26574 14530
rect 26626 14478 26638 14530
rect 22094 14466 22146 14478
rect 28142 14466 28194 14478
rect 28366 14530 28418 14542
rect 29934 14530 29986 14542
rect 37550 14530 37602 14542
rect 40910 14530 40962 14542
rect 28578 14478 28590 14530
rect 28642 14478 28654 14530
rect 29586 14478 29598 14530
rect 29650 14478 29662 14530
rect 31826 14478 31838 14530
rect 31890 14478 31902 14530
rect 32274 14478 32286 14530
rect 32338 14478 32350 14530
rect 33058 14478 33070 14530
rect 33122 14478 33134 14530
rect 34402 14478 34414 14530
rect 34466 14478 34478 14530
rect 35522 14478 35534 14530
rect 35586 14478 35598 14530
rect 38434 14478 38446 14530
rect 38498 14478 38510 14530
rect 39218 14478 39230 14530
rect 39282 14478 39294 14530
rect 28366 14466 28418 14478
rect 29934 14466 29986 14478
rect 37550 14466 37602 14478
rect 40910 14466 40962 14478
rect 41918 14530 41970 14542
rect 41918 14466 41970 14478
rect 42590 14530 42642 14542
rect 55246 14530 55298 14542
rect 57486 14530 57538 14542
rect 47506 14478 47518 14530
rect 47570 14478 47582 14530
rect 48514 14478 48526 14530
rect 48578 14478 48590 14530
rect 55010 14478 55022 14530
rect 55074 14478 55086 14530
rect 55906 14478 55918 14530
rect 55970 14478 55982 14530
rect 42590 14466 42642 14478
rect 55246 14466 55298 14478
rect 57486 14466 57538 14478
rect 60622 14530 60674 14542
rect 60622 14466 60674 14478
rect 4622 14418 4674 14430
rect 12574 14418 12626 14430
rect 9874 14366 9886 14418
rect 9938 14366 9950 14418
rect 4622 14354 4674 14366
rect 12574 14354 12626 14366
rect 12686 14418 12738 14430
rect 12686 14354 12738 14366
rect 13806 14418 13858 14430
rect 30382 14418 30434 14430
rect 34974 14418 35026 14430
rect 36094 14418 36146 14430
rect 41246 14418 41298 14430
rect 42366 14418 42418 14430
rect 47070 14418 47122 14430
rect 52894 14418 52946 14430
rect 15586 14366 15598 14418
rect 15650 14366 15662 14418
rect 19506 14366 19518 14418
rect 19570 14366 19582 14418
rect 24434 14366 24446 14418
rect 24498 14366 24510 14418
rect 30146 14366 30158 14418
rect 30210 14366 30222 14418
rect 31714 14366 31726 14418
rect 31778 14366 31790 14418
rect 34738 14366 34750 14418
rect 34802 14366 34814 14418
rect 35858 14366 35870 14418
rect 35922 14366 35934 14418
rect 40114 14366 40126 14418
rect 40178 14366 40190 14418
rect 41346 14366 41358 14418
rect 41410 14366 41422 14418
rect 43698 14366 43710 14418
rect 43762 14366 43774 14418
rect 46162 14366 46174 14418
rect 46226 14366 46238 14418
rect 47618 14366 47630 14418
rect 47682 14366 47694 14418
rect 49746 14366 49758 14418
rect 49810 14366 49822 14418
rect 13806 14354 13858 14366
rect 30382 14354 30434 14366
rect 34974 14354 35026 14366
rect 36094 14354 36146 14366
rect 41246 14354 41298 14366
rect 42366 14354 42418 14366
rect 47070 14354 47122 14366
rect 52894 14354 52946 14366
rect 57710 14418 57762 14430
rect 57710 14354 57762 14366
rect 1934 14306 1986 14318
rect 1934 14242 1986 14254
rect 2942 14306 2994 14318
rect 2942 14242 2994 14254
rect 4846 14306 4898 14318
rect 4846 14242 4898 14254
rect 5070 14306 5122 14318
rect 5070 14242 5122 14254
rect 6302 14306 6354 14318
rect 14590 14306 14642 14318
rect 9202 14254 9214 14306
rect 9266 14254 9278 14306
rect 14242 14254 14254 14306
rect 14306 14254 14318 14306
rect 6302 14242 6354 14254
rect 14590 14242 14642 14254
rect 15262 14306 15314 14318
rect 15262 14242 15314 14254
rect 17838 14306 17890 14318
rect 17838 14242 17890 14254
rect 20638 14306 20690 14318
rect 20638 14242 20690 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 25342 14306 25394 14318
rect 25342 14242 25394 14254
rect 28478 14306 28530 14318
rect 28478 14242 28530 14254
rect 29150 14306 29202 14318
rect 29150 14242 29202 14254
rect 29598 14306 29650 14318
rect 29598 14242 29650 14254
rect 30830 14306 30882 14318
rect 30830 14242 30882 14254
rect 34190 14306 34242 14318
rect 34190 14242 34242 14254
rect 37998 14306 38050 14318
rect 37998 14242 38050 14254
rect 41134 14306 41186 14318
rect 41134 14242 41186 14254
rect 51662 14306 51714 14318
rect 51662 14242 51714 14254
rect 51998 14306 52050 14318
rect 51998 14242 52050 14254
rect 57934 14306 57986 14318
rect 57934 14242 57986 14254
rect 58606 14306 58658 14318
rect 58606 14242 58658 14254
rect 59278 14306 59330 14318
rect 59278 14242 59330 14254
rect 59726 14306 59778 14318
rect 59726 14242 59778 14254
rect 1344 14138 62608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 62608 14138
rect 1344 14052 62608 14086
rect 2158 13970 2210 13982
rect 2158 13906 2210 13918
rect 2718 13970 2770 13982
rect 2718 13906 2770 13918
rect 3054 13970 3106 13982
rect 3054 13906 3106 13918
rect 3614 13970 3666 13982
rect 3614 13906 3666 13918
rect 7198 13970 7250 13982
rect 7198 13906 7250 13918
rect 8878 13970 8930 13982
rect 23998 13970 24050 13982
rect 17938 13918 17950 13970
rect 18002 13918 18014 13970
rect 18946 13918 18958 13970
rect 19010 13918 19022 13970
rect 21746 13918 21758 13970
rect 21810 13918 21822 13970
rect 8878 13906 8930 13918
rect 23998 13906 24050 13918
rect 24334 13970 24386 13982
rect 24334 13906 24386 13918
rect 24558 13970 24610 13982
rect 24558 13906 24610 13918
rect 25454 13970 25506 13982
rect 25454 13906 25506 13918
rect 32286 13970 32338 13982
rect 41134 13970 41186 13982
rect 35634 13918 35646 13970
rect 35698 13918 35710 13970
rect 37202 13918 37214 13970
rect 37266 13918 37278 13970
rect 38434 13918 38446 13970
rect 38498 13918 38510 13970
rect 32286 13906 32338 13918
rect 41134 13906 41186 13918
rect 41358 13970 41410 13982
rect 47854 13970 47906 13982
rect 46722 13918 46734 13970
rect 46786 13918 46798 13970
rect 41358 13906 41410 13918
rect 47854 13906 47906 13918
rect 48862 13970 48914 13982
rect 48862 13906 48914 13918
rect 49758 13970 49810 13982
rect 49758 13906 49810 13918
rect 50654 13970 50706 13982
rect 50654 13906 50706 13918
rect 58046 13970 58098 13982
rect 58046 13906 58098 13918
rect 58494 13970 58546 13982
rect 58494 13906 58546 13918
rect 59390 13970 59442 13982
rect 59390 13906 59442 13918
rect 60286 13970 60338 13982
rect 60286 13906 60338 13918
rect 61182 13970 61234 13982
rect 61182 13906 61234 13918
rect 61742 13970 61794 13982
rect 61742 13906 61794 13918
rect 62190 13970 62242 13982
rect 62190 13906 62242 13918
rect 8542 13858 8594 13870
rect 18622 13858 18674 13870
rect 22318 13858 22370 13870
rect 24670 13858 24722 13870
rect 5618 13806 5630 13858
rect 5682 13806 5694 13858
rect 7298 13806 7310 13858
rect 7362 13806 7374 13858
rect 16258 13806 16270 13858
rect 16322 13806 16334 13858
rect 19730 13806 19742 13858
rect 19794 13806 19806 13858
rect 23090 13806 23102 13858
rect 23154 13806 23166 13858
rect 8542 13794 8594 13806
rect 18622 13794 18674 13806
rect 22318 13794 22370 13806
rect 24670 13794 24722 13806
rect 26462 13858 26514 13870
rect 49086 13858 49138 13870
rect 27570 13806 27582 13858
rect 27634 13806 27646 13858
rect 33394 13806 33406 13858
rect 33458 13806 33470 13858
rect 33954 13806 33966 13858
rect 34018 13806 34030 13858
rect 35410 13806 35422 13858
rect 35474 13806 35486 13858
rect 39330 13806 39342 13858
rect 39394 13806 39406 13858
rect 39554 13806 39566 13858
rect 39618 13806 39630 13858
rect 42130 13806 42142 13858
rect 42194 13806 42206 13858
rect 26462 13794 26514 13806
rect 49086 13794 49138 13806
rect 50206 13858 50258 13870
rect 60734 13858 60786 13870
rect 52322 13806 52334 13858
rect 52386 13806 52398 13858
rect 50206 13794 50258 13806
rect 60734 13794 60786 13806
rect 6302 13746 6354 13758
rect 4834 13694 4846 13746
rect 4898 13694 4910 13746
rect 5842 13694 5854 13746
rect 5906 13694 5918 13746
rect 6302 13682 6354 13694
rect 7086 13746 7138 13758
rect 7086 13682 7138 13694
rect 7534 13746 7586 13758
rect 8766 13746 8818 13758
rect 7858 13694 7870 13746
rect 7922 13694 7934 13746
rect 7534 13682 7586 13694
rect 8766 13682 8818 13694
rect 8990 13746 9042 13758
rect 15038 13746 15090 13758
rect 9650 13694 9662 13746
rect 9714 13694 9726 13746
rect 9986 13694 9998 13746
rect 10050 13694 10062 13746
rect 10994 13694 11006 13746
rect 11058 13694 11070 13746
rect 11554 13694 11566 13746
rect 11618 13694 11630 13746
rect 12338 13694 12350 13746
rect 12402 13694 12414 13746
rect 8990 13682 9042 13694
rect 15038 13682 15090 13694
rect 17390 13746 17442 13758
rect 17390 13682 17442 13694
rect 17614 13746 17666 13758
rect 17614 13682 17666 13694
rect 22094 13746 22146 13758
rect 29934 13746 29986 13758
rect 22866 13694 22878 13746
rect 22930 13694 22942 13746
rect 25666 13694 25678 13746
rect 25730 13694 25742 13746
rect 26226 13694 26238 13746
rect 26290 13694 26302 13746
rect 26898 13694 26910 13746
rect 26962 13694 26974 13746
rect 22094 13682 22146 13694
rect 29934 13682 29986 13694
rect 30494 13746 30546 13758
rect 31838 13746 31890 13758
rect 35198 13746 35250 13758
rect 36878 13746 36930 13758
rect 30818 13694 30830 13746
rect 30882 13694 30894 13746
rect 33282 13694 33294 13746
rect 33346 13694 33358 13746
rect 34514 13694 34526 13746
rect 34578 13694 34590 13746
rect 34850 13694 34862 13746
rect 34914 13694 34926 13746
rect 35970 13694 35982 13746
rect 36034 13694 36046 13746
rect 30494 13682 30546 13694
rect 31838 13682 31890 13694
rect 35198 13682 35250 13694
rect 36878 13682 36930 13694
rect 37550 13746 37602 13758
rect 37550 13682 37602 13694
rect 38110 13746 38162 13758
rect 38110 13682 38162 13694
rect 39902 13746 39954 13758
rect 39902 13682 39954 13694
rect 41022 13746 41074 13758
rect 43262 13746 43314 13758
rect 48750 13746 48802 13758
rect 42242 13694 42254 13746
rect 42306 13694 42318 13746
rect 43698 13694 43710 13746
rect 43762 13694 43774 13746
rect 41022 13682 41074 13694
rect 43262 13682 43314 13694
rect 48750 13682 48802 13694
rect 49198 13746 49250 13758
rect 49198 13682 49250 13694
rect 49534 13746 49586 13758
rect 49534 13682 49586 13694
rect 49982 13746 50034 13758
rect 51438 13746 51490 13758
rect 50978 13694 50990 13746
rect 51042 13743 51054 13746
rect 51202 13743 51214 13746
rect 51042 13697 51214 13743
rect 51042 13694 51054 13697
rect 51202 13694 51214 13697
rect 51266 13694 51278 13746
rect 49982 13682 50034 13694
rect 51438 13682 51490 13694
rect 51774 13746 51826 13758
rect 56590 13746 56642 13758
rect 52546 13694 52558 13746
rect 52610 13694 52622 13746
rect 53330 13694 53342 13746
rect 53394 13694 53406 13746
rect 54562 13694 54574 13746
rect 54626 13694 54638 13746
rect 55346 13694 55358 13746
rect 55410 13694 55422 13746
rect 51774 13682 51826 13694
rect 56590 13682 56642 13694
rect 56814 13746 56866 13758
rect 59838 13746 59890 13758
rect 57138 13694 57150 13746
rect 57202 13694 57214 13746
rect 56814 13682 56866 13694
rect 59838 13682 59890 13694
rect 4174 13634 4226 13646
rect 21534 13634 21586 13646
rect 3938 13582 3950 13634
rect 4002 13582 4014 13634
rect 4610 13582 4622 13634
rect 4674 13582 4686 13634
rect 14466 13582 14478 13634
rect 14530 13582 14542 13634
rect 4174 13570 4226 13582
rect 21534 13570 21586 13582
rect 23662 13634 23714 13646
rect 30382 13634 30434 13646
rect 29698 13582 29710 13634
rect 29762 13582 29774 13634
rect 23662 13570 23714 13582
rect 30382 13570 30434 13582
rect 37886 13634 37938 13646
rect 57598 13634 57650 13646
rect 53890 13582 53902 13634
rect 53954 13582 53966 13634
rect 37886 13570 37938 13582
rect 57598 13570 57650 13582
rect 58942 13634 58994 13646
rect 58942 13570 58994 13582
rect 6638 13522 6690 13534
rect 10782 13522 10834 13534
rect 7970 13470 7982 13522
rect 8034 13519 8046 13522
rect 8194 13519 8206 13522
rect 8034 13473 8206 13519
rect 8034 13470 8046 13473
rect 8194 13470 8206 13473
rect 8258 13470 8270 13522
rect 6638 13458 6690 13470
rect 10782 13458 10834 13470
rect 35646 13522 35698 13534
rect 36654 13522 36706 13534
rect 36306 13470 36318 13522
rect 36370 13470 36382 13522
rect 35646 13458 35698 13470
rect 36654 13458 36706 13470
rect 40238 13522 40290 13534
rect 45390 13522 45442 13534
rect 44482 13470 44494 13522
rect 44546 13470 44558 13522
rect 40238 13458 40290 13470
rect 45390 13458 45442 13470
rect 1344 13354 62608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 62608 13354
rect 1344 13268 62608 13302
rect 4958 13186 5010 13198
rect 38894 13186 38946 13198
rect 54686 13186 54738 13198
rect 1586 13134 1598 13186
rect 1650 13183 1662 13186
rect 2930 13183 2942 13186
rect 1650 13137 2942 13183
rect 1650 13134 1662 13137
rect 2930 13134 2942 13137
rect 2994 13134 3006 13186
rect 7522 13134 7534 13186
rect 7586 13134 7598 13186
rect 15586 13134 15598 13186
rect 15650 13134 15662 13186
rect 16818 13134 16830 13186
rect 16882 13134 16894 13186
rect 23202 13134 23214 13186
rect 23266 13134 23278 13186
rect 35522 13134 35534 13186
rect 35586 13134 35598 13186
rect 41906 13134 41918 13186
rect 41970 13134 41982 13186
rect 45378 13134 45390 13186
rect 45442 13183 45454 13186
rect 45826 13183 45838 13186
rect 45442 13137 45838 13183
rect 45442 13134 45454 13137
rect 45826 13134 45838 13137
rect 45890 13134 45902 13186
rect 4958 13122 5010 13134
rect 38894 13122 38946 13134
rect 54686 13122 54738 13134
rect 2046 13074 2098 13086
rect 2046 13010 2098 13022
rect 2942 13074 2994 13086
rect 18958 13074 19010 13086
rect 7634 13022 7646 13074
rect 7698 13022 7710 13074
rect 9202 13022 9214 13074
rect 9266 13022 9278 13074
rect 9874 13022 9886 13074
rect 9938 13022 9950 13074
rect 12002 13022 12014 13074
rect 12066 13022 12078 13074
rect 17938 13022 17950 13074
rect 18002 13022 18014 13074
rect 2942 13010 2994 13022
rect 18958 13010 19010 13022
rect 19854 13074 19906 13086
rect 29262 13074 29314 13086
rect 38670 13074 38722 13086
rect 21298 13022 21310 13074
rect 21362 13022 21374 13074
rect 30146 13022 30158 13074
rect 30210 13022 30222 13074
rect 34514 13022 34526 13074
rect 34578 13022 34590 13074
rect 35298 13022 35310 13074
rect 35362 13022 35374 13074
rect 19854 13010 19906 13022
rect 29262 13010 29314 13022
rect 38670 13010 38722 13022
rect 39230 13074 39282 13086
rect 45390 13074 45442 13086
rect 49982 13074 50034 13086
rect 40674 13022 40686 13074
rect 40738 13022 40750 13074
rect 43362 13022 43374 13074
rect 43426 13022 43438 13074
rect 46834 13022 46846 13074
rect 46898 13022 46910 13074
rect 39230 13010 39282 13022
rect 45390 13010 45442 13022
rect 49982 13010 50034 13022
rect 51438 13074 51490 13086
rect 51438 13010 51490 13022
rect 53342 13074 53394 13086
rect 53342 13010 53394 13022
rect 56926 13074 56978 13086
rect 56926 13010 56978 13022
rect 57374 13074 57426 13086
rect 57374 13010 57426 13022
rect 57822 13074 57874 13086
rect 57822 13010 57874 13022
rect 58830 13074 58882 13086
rect 58830 13010 58882 13022
rect 59166 13074 59218 13086
rect 59166 13010 59218 13022
rect 59614 13074 59666 13086
rect 59614 13010 59666 13022
rect 61854 13074 61906 13086
rect 61854 13010 61906 13022
rect 62302 13074 62354 13086
rect 62302 13010 62354 13022
rect 5966 12962 6018 12974
rect 17054 12962 17106 12974
rect 22654 12962 22706 12974
rect 23998 12962 24050 12974
rect 6178 12910 6190 12962
rect 6242 12910 6254 12962
rect 8642 12910 8654 12962
rect 8706 12910 8718 12962
rect 8978 12910 8990 12962
rect 9042 12910 9054 12962
rect 12674 12910 12686 12962
rect 12738 12910 12750 12962
rect 16594 12910 16606 12962
rect 16658 12910 16670 12962
rect 20626 12910 20638 12962
rect 20690 12910 20702 12962
rect 21410 12910 21422 12962
rect 21474 12910 21486 12962
rect 21634 12910 21646 12962
rect 21698 12910 21710 12962
rect 22866 12910 22878 12962
rect 22930 12910 22942 12962
rect 23426 12910 23438 12962
rect 23490 12910 23502 12962
rect 5966 12898 6018 12910
rect 17054 12898 17106 12910
rect 22654 12898 22706 12910
rect 23998 12898 24050 12910
rect 24334 12962 24386 12974
rect 24334 12898 24386 12910
rect 25006 12962 25058 12974
rect 35198 12962 35250 12974
rect 37438 12962 37490 12974
rect 41470 12962 41522 12974
rect 43822 12962 43874 12974
rect 47742 12962 47794 12974
rect 51662 12962 51714 12974
rect 55022 12962 55074 12974
rect 25890 12910 25902 12962
rect 25954 12910 25966 12962
rect 29698 12910 29710 12962
rect 29762 12910 29774 12962
rect 31042 12910 31054 12962
rect 31106 12910 31118 12962
rect 31266 12910 31278 12962
rect 31330 12910 31342 12962
rect 34402 12910 34414 12962
rect 34466 12910 34478 12962
rect 35522 12910 35534 12962
rect 35586 12910 35598 12962
rect 41010 12910 41022 12962
rect 41074 12910 41086 12962
rect 42690 12910 42702 12962
rect 42754 12910 42766 12962
rect 46722 12910 46734 12962
rect 46786 12910 46798 12962
rect 47282 12910 47294 12962
rect 47346 12910 47358 12962
rect 50978 12910 50990 12962
rect 51042 12910 51054 12962
rect 54114 12910 54126 12962
rect 54178 12910 54190 12962
rect 25006 12898 25058 12910
rect 35198 12898 35250 12910
rect 37438 12898 37490 12910
rect 41470 12898 41522 12910
rect 43822 12898 43874 12910
rect 47742 12898 47794 12910
rect 51662 12898 51714 12910
rect 55022 12898 55074 12910
rect 56590 12962 56642 12974
rect 56590 12898 56642 12910
rect 5630 12850 5682 12862
rect 3826 12798 3838 12850
rect 3890 12798 3902 12850
rect 5630 12786 5682 12798
rect 6526 12850 6578 12862
rect 6526 12786 6578 12798
rect 7982 12850 8034 12862
rect 17390 12850 17442 12862
rect 14018 12798 14030 12850
rect 14082 12798 14094 12850
rect 7982 12786 8034 12798
rect 17390 12786 17442 12798
rect 18174 12850 18226 12862
rect 18174 12786 18226 12798
rect 18510 12850 18562 12862
rect 18510 12786 18562 12798
rect 18734 12850 18786 12862
rect 18734 12786 18786 12798
rect 19070 12850 19122 12862
rect 19070 12786 19122 12798
rect 19518 12850 19570 12862
rect 21870 12850 21922 12862
rect 20402 12798 20414 12850
rect 20466 12798 20478 12850
rect 19518 12786 19570 12798
rect 21870 12786 21922 12798
rect 23774 12850 23826 12862
rect 23774 12786 23826 12798
rect 24670 12850 24722 12862
rect 30606 12850 30658 12862
rect 44270 12850 44322 12862
rect 27794 12798 27806 12850
rect 27858 12798 27870 12850
rect 34066 12798 34078 12850
rect 34130 12798 34142 12850
rect 37650 12798 37662 12850
rect 37714 12798 37726 12850
rect 37986 12798 37998 12850
rect 38050 12798 38062 12850
rect 24670 12786 24722 12798
rect 30606 12786 30658 12798
rect 44270 12786 44322 12798
rect 44942 12850 44994 12862
rect 47630 12850 47682 12862
rect 50542 12850 50594 12862
rect 46050 12798 46062 12850
rect 46114 12798 46126 12850
rect 48290 12798 48302 12850
rect 48354 12798 48366 12850
rect 48514 12798 48526 12850
rect 48578 12798 48590 12850
rect 49186 12798 49198 12850
rect 49250 12798 49262 12850
rect 44942 12786 44994 12798
rect 47630 12786 47682 12798
rect 50542 12786 50594 12798
rect 50654 12850 50706 12862
rect 56254 12850 56306 12862
rect 54002 12798 54014 12850
rect 54066 12798 54078 12850
rect 55234 12798 55246 12850
rect 55298 12798 55310 12850
rect 55794 12798 55806 12850
rect 55858 12798 55870 12850
rect 50654 12786 50706 12798
rect 56254 12786 56306 12798
rect 56366 12850 56418 12862
rect 56366 12786 56418 12798
rect 58270 12850 58322 12862
rect 58270 12786 58322 12798
rect 2494 12738 2546 12750
rect 2494 12674 2546 12686
rect 5742 12738 5794 12750
rect 5742 12674 5794 12686
rect 9662 12738 9714 12750
rect 22094 12738 22146 12750
rect 24222 12738 24274 12750
rect 16930 12686 16942 12738
rect 16994 12686 17006 12738
rect 23090 12686 23102 12738
rect 23154 12686 23166 12738
rect 9662 12674 9714 12686
rect 22094 12674 22146 12686
rect 24222 12674 24274 12686
rect 25790 12738 25842 12750
rect 25790 12674 25842 12686
rect 26350 12738 26402 12750
rect 26350 12674 26402 12686
rect 29150 12738 29202 12750
rect 29150 12674 29202 12686
rect 29374 12738 29426 12750
rect 29374 12674 29426 12686
rect 37102 12738 37154 12750
rect 37102 12674 37154 12686
rect 49534 12738 49586 12750
rect 49534 12674 49586 12686
rect 50318 12738 50370 12750
rect 50318 12674 50370 12686
rect 50430 12738 50482 12750
rect 53006 12738 53058 12750
rect 51986 12686 51998 12738
rect 52050 12686 52062 12738
rect 50430 12674 50482 12686
rect 53006 12674 53058 12686
rect 1344 12570 62608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 62608 12570
rect 1344 12484 62608 12518
rect 3278 12402 3330 12414
rect 3278 12338 3330 12350
rect 4510 12402 4562 12414
rect 16382 12402 16434 12414
rect 11218 12350 11230 12402
rect 11282 12350 11294 12402
rect 4510 12338 4562 12350
rect 16382 12338 16434 12350
rect 17614 12402 17666 12414
rect 17614 12338 17666 12350
rect 18398 12402 18450 12414
rect 18398 12338 18450 12350
rect 23774 12402 23826 12414
rect 23774 12338 23826 12350
rect 25342 12402 25394 12414
rect 28254 12402 28306 12414
rect 35870 12402 35922 12414
rect 27122 12350 27134 12402
rect 27186 12350 27198 12402
rect 29922 12350 29934 12402
rect 29986 12350 29998 12402
rect 25342 12338 25394 12350
rect 28254 12338 28306 12350
rect 35870 12338 35922 12350
rect 38334 12402 38386 12414
rect 38334 12338 38386 12350
rect 40014 12402 40066 12414
rect 40014 12338 40066 12350
rect 41470 12402 41522 12414
rect 41470 12338 41522 12350
rect 44158 12402 44210 12414
rect 49198 12402 49250 12414
rect 45042 12350 45054 12402
rect 45106 12350 45118 12402
rect 44158 12338 44210 12350
rect 49198 12338 49250 12350
rect 55134 12402 55186 12414
rect 56590 12402 56642 12414
rect 55458 12350 55470 12402
rect 55522 12350 55534 12402
rect 55134 12338 55186 12350
rect 56590 12338 56642 12350
rect 57934 12402 57986 12414
rect 57934 12338 57986 12350
rect 58830 12402 58882 12414
rect 58830 12338 58882 12350
rect 59614 12402 59666 12414
rect 59614 12338 59666 12350
rect 2046 12290 2098 12302
rect 2046 12226 2098 12238
rect 4062 12290 4114 12302
rect 13134 12290 13186 12302
rect 10322 12238 10334 12290
rect 10386 12238 10398 12290
rect 4062 12226 4114 12238
rect 13134 12226 13186 12238
rect 13582 12290 13634 12302
rect 16830 12290 16882 12302
rect 15250 12238 15262 12290
rect 15314 12238 15326 12290
rect 15922 12238 15934 12290
rect 15986 12238 15998 12290
rect 13582 12226 13634 12238
rect 16830 12226 16882 12238
rect 18622 12290 18674 12302
rect 18622 12226 18674 12238
rect 18734 12290 18786 12302
rect 18734 12226 18786 12238
rect 19630 12290 19682 12302
rect 22094 12290 22146 12302
rect 20178 12238 20190 12290
rect 20242 12238 20254 12290
rect 19630 12226 19682 12238
rect 22094 12226 22146 12238
rect 22318 12290 22370 12302
rect 22318 12226 22370 12238
rect 22990 12290 23042 12302
rect 24334 12290 24386 12302
rect 23202 12238 23214 12290
rect 23266 12238 23278 12290
rect 22990 12226 23042 12238
rect 24334 12226 24386 12238
rect 26126 12290 26178 12302
rect 33182 12290 33234 12302
rect 29250 12238 29262 12290
rect 29314 12238 29326 12290
rect 26126 12226 26178 12238
rect 33182 12226 33234 12238
rect 33294 12290 33346 12302
rect 41246 12290 41298 12302
rect 33954 12238 33966 12290
rect 34018 12238 34030 12290
rect 39106 12238 39118 12290
rect 39170 12238 39182 12290
rect 33294 12226 33346 12238
rect 41246 12226 41298 12238
rect 41694 12290 41746 12302
rect 47182 12290 47234 12302
rect 43362 12238 43374 12290
rect 43426 12238 43438 12290
rect 44706 12238 44718 12290
rect 44770 12238 44782 12290
rect 41694 12226 41746 12238
rect 47182 12226 47234 12238
rect 49758 12290 49810 12302
rect 56926 12290 56978 12302
rect 51202 12238 51214 12290
rect 51266 12238 51278 12290
rect 52658 12238 52670 12290
rect 52722 12238 52734 12290
rect 53330 12238 53342 12290
rect 53394 12238 53406 12290
rect 49758 12226 49810 12238
rect 56926 12226 56978 12238
rect 1710 12178 1762 12190
rect 8206 12178 8258 12190
rect 6066 12126 6078 12178
rect 6130 12126 6142 12178
rect 1710 12114 1762 12126
rect 8206 12114 8258 12126
rect 8542 12178 8594 12190
rect 13246 12178 13298 12190
rect 9538 12126 9550 12178
rect 9602 12126 9614 12178
rect 10210 12126 10222 12178
rect 10274 12126 10286 12178
rect 12450 12126 12462 12178
rect 12514 12126 12526 12178
rect 13010 12126 13022 12178
rect 13074 12126 13086 12178
rect 8542 12114 8594 12126
rect 13246 12114 13298 12126
rect 13806 12178 13858 12190
rect 13806 12114 13858 12126
rect 14254 12178 14306 12190
rect 14254 12114 14306 12126
rect 14590 12178 14642 12190
rect 15598 12178 15650 12190
rect 15026 12126 15038 12178
rect 15090 12126 15102 12178
rect 14590 12114 14642 12126
rect 15598 12114 15650 12126
rect 16270 12178 16322 12190
rect 16270 12114 16322 12126
rect 16494 12178 16546 12190
rect 16494 12114 16546 12126
rect 17390 12178 17442 12190
rect 17390 12114 17442 12126
rect 17838 12178 17890 12190
rect 17838 12114 17890 12126
rect 17950 12178 18002 12190
rect 19742 12178 19794 12190
rect 20750 12178 20802 12190
rect 22766 12178 22818 12190
rect 19058 12126 19070 12178
rect 19122 12126 19134 12178
rect 20066 12126 20078 12178
rect 20130 12126 20142 12178
rect 21074 12126 21086 12178
rect 21138 12126 21150 12178
rect 17950 12114 18002 12126
rect 19742 12114 19794 12126
rect 20750 12114 20802 12126
rect 22766 12114 22818 12126
rect 23438 12178 23490 12190
rect 24110 12178 24162 12190
rect 23650 12126 23662 12178
rect 23714 12126 23726 12178
rect 23438 12114 23490 12126
rect 24110 12114 24162 12126
rect 24782 12178 24834 12190
rect 25678 12178 25730 12190
rect 32958 12178 33010 12190
rect 39678 12178 39730 12190
rect 48190 12178 48242 12190
rect 25330 12126 25342 12178
rect 25394 12126 25406 12178
rect 25890 12126 25902 12178
rect 25954 12126 25966 12178
rect 28914 12126 28926 12178
rect 28978 12126 28990 12178
rect 30594 12126 30606 12178
rect 30658 12126 30670 12178
rect 31938 12126 31950 12178
rect 32002 12126 32014 12178
rect 36082 12126 36094 12178
rect 36146 12126 36158 12178
rect 37314 12126 37326 12178
rect 37378 12126 37390 12178
rect 37874 12126 37886 12178
rect 37938 12126 37950 12178
rect 38882 12126 38894 12178
rect 38946 12126 38958 12178
rect 41906 12126 41918 12178
rect 41970 12126 41982 12178
rect 42690 12126 42702 12178
rect 42754 12126 42766 12178
rect 44258 12126 44270 12178
rect 44322 12126 44334 12178
rect 45042 12126 45054 12178
rect 45106 12126 45118 12178
rect 45602 12126 45614 12178
rect 45666 12126 45678 12178
rect 46162 12126 46174 12178
rect 46226 12126 46238 12178
rect 46946 12126 46958 12178
rect 47010 12126 47022 12178
rect 47954 12126 47966 12178
rect 48018 12126 48030 12178
rect 24782 12114 24834 12126
rect 25678 12114 25730 12126
rect 32958 12114 33010 12126
rect 39678 12114 39730 12126
rect 48190 12114 48242 12126
rect 48750 12178 48802 12190
rect 48750 12114 48802 12126
rect 48974 12178 49026 12190
rect 48974 12114 49026 12126
rect 49310 12178 49362 12190
rect 58270 12178 58322 12190
rect 50530 12126 50542 12178
rect 50594 12126 50606 12178
rect 52210 12126 52222 12178
rect 52274 12126 52286 12178
rect 55682 12126 55694 12178
rect 55746 12126 55758 12178
rect 49310 12114 49362 12126
rect 58270 12114 58322 12126
rect 2830 12066 2882 12078
rect 2830 12002 2882 12014
rect 3726 12066 3778 12078
rect 11790 12066 11842 12078
rect 4946 12014 4958 12066
rect 5010 12014 5022 12066
rect 5954 12014 5966 12066
rect 6018 12014 6030 12066
rect 7858 12014 7870 12066
rect 7922 12014 7934 12066
rect 10098 12014 10110 12066
rect 10162 12014 10174 12066
rect 3726 12002 3778 12014
rect 11790 12002 11842 12014
rect 14030 12066 14082 12078
rect 20862 12066 20914 12078
rect 19170 12014 19182 12066
rect 19234 12014 19246 12066
rect 14030 12002 14082 12014
rect 20862 12002 20914 12014
rect 22542 12066 22594 12078
rect 22542 12002 22594 12014
rect 24558 12066 24610 12078
rect 24558 12002 24610 12014
rect 41806 12066 41858 12078
rect 57374 12066 57426 12078
rect 42578 12014 42590 12066
rect 42642 12014 42654 12066
rect 47058 12014 47070 12066
rect 47122 12014 47134 12066
rect 41806 12002 41858 12014
rect 57374 12002 57426 12014
rect 59166 12066 59218 12078
rect 59166 12002 59218 12014
rect 4174 11954 4226 11966
rect 4174 11890 4226 11902
rect 11566 11954 11618 11966
rect 14478 11954 14530 11966
rect 12674 11902 12686 11954
rect 12738 11902 12750 11954
rect 11566 11890 11618 11902
rect 14478 11890 14530 11902
rect 19630 11954 19682 11966
rect 19630 11890 19682 11902
rect 1344 11786 62608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 62608 11786
rect 1344 11700 62608 11734
rect 6862 11618 6914 11630
rect 6862 11554 6914 11566
rect 12126 11618 12178 11630
rect 12126 11554 12178 11566
rect 12798 11618 12850 11630
rect 12798 11554 12850 11566
rect 12910 11618 12962 11630
rect 12910 11554 12962 11566
rect 16830 11618 16882 11630
rect 16830 11554 16882 11566
rect 28030 11618 28082 11630
rect 28030 11554 28082 11566
rect 28366 11618 28418 11630
rect 34302 11618 34354 11630
rect 38110 11618 38162 11630
rect 55582 11618 55634 11630
rect 30594 11566 30606 11618
rect 30658 11566 30670 11618
rect 37538 11566 37550 11618
rect 37602 11566 37614 11618
rect 50530 11566 50542 11618
rect 50594 11566 50606 11618
rect 56242 11566 56254 11618
rect 56306 11615 56318 11618
rect 56690 11615 56702 11618
rect 56306 11569 56702 11615
rect 56306 11566 56318 11569
rect 56690 11566 56702 11569
rect 56754 11566 56766 11618
rect 28366 11554 28418 11566
rect 34302 11554 34354 11566
rect 38110 11554 38162 11566
rect 55582 11554 55634 11566
rect 2494 11506 2546 11518
rect 11790 11506 11842 11518
rect 9874 11454 9886 11506
rect 9938 11454 9950 11506
rect 2494 11442 2546 11454
rect 11790 11442 11842 11454
rect 16270 11506 16322 11518
rect 31838 11506 31890 11518
rect 17826 11454 17838 11506
rect 17890 11454 17902 11506
rect 25106 11454 25118 11506
rect 25170 11454 25182 11506
rect 29586 11454 29598 11506
rect 29650 11454 29662 11506
rect 16270 11442 16322 11454
rect 31838 11442 31890 11454
rect 33406 11506 33458 11518
rect 33406 11442 33458 11454
rect 35870 11506 35922 11518
rect 35870 11442 35922 11454
rect 36990 11506 37042 11518
rect 36990 11442 37042 11454
rect 37214 11506 37266 11518
rect 37214 11442 37266 11454
rect 42814 11506 42866 11518
rect 42814 11442 42866 11454
rect 44942 11506 44994 11518
rect 44942 11442 44994 11454
rect 46174 11506 46226 11518
rect 46174 11442 46226 11454
rect 46846 11506 46898 11518
rect 49422 11506 49474 11518
rect 49074 11454 49086 11506
rect 49138 11454 49150 11506
rect 46846 11442 46898 11454
rect 49422 11442 49474 11454
rect 56254 11506 56306 11518
rect 56254 11442 56306 11454
rect 56702 11506 56754 11518
rect 56702 11442 56754 11454
rect 57150 11506 57202 11518
rect 57150 11442 57202 11454
rect 57598 11506 57650 11518
rect 57598 11442 57650 11454
rect 58046 11506 58098 11518
rect 58046 11442 58098 11454
rect 6526 11394 6578 11406
rect 12350 11394 12402 11406
rect 5730 11342 5742 11394
rect 5794 11342 5806 11394
rect 7410 11342 7422 11394
rect 7474 11342 7486 11394
rect 7746 11342 7758 11394
rect 7810 11342 7822 11394
rect 10770 11342 10782 11394
rect 10834 11342 10846 11394
rect 6526 11330 6578 11342
rect 12350 11330 12402 11342
rect 13358 11394 13410 11406
rect 17054 11394 17106 11406
rect 21870 11394 21922 11406
rect 26574 11394 26626 11406
rect 16706 11342 16718 11394
rect 16770 11342 16782 11394
rect 17602 11342 17614 11394
rect 17666 11342 17678 11394
rect 17938 11342 17950 11394
rect 18002 11342 18014 11394
rect 19058 11342 19070 11394
rect 19122 11342 19134 11394
rect 19506 11342 19518 11394
rect 19570 11342 19582 11394
rect 20290 11342 20302 11394
rect 20354 11342 20366 11394
rect 22306 11342 22318 11394
rect 22370 11342 22382 11394
rect 25666 11342 25678 11394
rect 25730 11342 25742 11394
rect 13358 11330 13410 11342
rect 17054 11330 17106 11342
rect 21870 11330 21922 11342
rect 26574 11330 26626 11342
rect 26798 11394 26850 11406
rect 29150 11394 29202 11406
rect 32286 11394 32338 11406
rect 27346 11342 27358 11394
rect 27410 11342 27422 11394
rect 31378 11342 31390 11394
rect 31442 11342 31454 11394
rect 26798 11330 26850 11342
rect 29150 11330 29202 11342
rect 32286 11330 32338 11342
rect 33294 11394 33346 11406
rect 33294 11330 33346 11342
rect 33518 11394 33570 11406
rect 40350 11394 40402 11406
rect 41806 11394 41858 11406
rect 35074 11342 35086 11394
rect 35138 11342 35150 11394
rect 41234 11342 41246 11394
rect 41298 11342 41310 11394
rect 33518 11330 33570 11342
rect 40350 11330 40402 11342
rect 41806 11330 41858 11342
rect 42030 11394 42082 11406
rect 42030 11330 42082 11342
rect 42366 11394 42418 11406
rect 42366 11330 42418 11342
rect 43038 11394 43090 11406
rect 43038 11330 43090 11342
rect 43262 11394 43314 11406
rect 45390 11394 45442 11406
rect 44146 11342 44158 11394
rect 44210 11342 44222 11394
rect 43262 11330 43314 11342
rect 45390 11330 45442 11342
rect 46398 11394 46450 11406
rect 46398 11330 46450 11342
rect 47630 11394 47682 11406
rect 47630 11330 47682 11342
rect 47966 11394 48018 11406
rect 50878 11394 50930 11406
rect 48962 11342 48974 11394
rect 49026 11342 49038 11394
rect 49858 11342 49870 11394
rect 49922 11342 49934 11394
rect 47966 11330 48018 11342
rect 50878 11330 50930 11342
rect 51102 11394 51154 11406
rect 51762 11342 51774 11394
rect 51826 11342 51838 11394
rect 51102 11330 51154 11342
rect 4958 11282 5010 11294
rect 12686 11282 12738 11294
rect 16494 11282 16546 11294
rect 20750 11282 20802 11294
rect 25902 11282 25954 11294
rect 30382 11282 30434 11294
rect 40686 11282 40738 11294
rect 42702 11282 42754 11294
rect 3602 11230 3614 11282
rect 3666 11230 3678 11282
rect 5842 11230 5854 11282
rect 5906 11230 5918 11282
rect 10434 11230 10446 11282
rect 10498 11230 10510 11282
rect 15138 11230 15150 11282
rect 15202 11230 15214 11282
rect 18610 11230 18622 11282
rect 18674 11230 18686 11282
rect 18946 11230 18958 11282
rect 19010 11230 19022 11282
rect 22978 11230 22990 11282
rect 23042 11230 23054 11282
rect 27234 11230 27246 11282
rect 27298 11230 27310 11282
rect 34850 11230 34862 11282
rect 34914 11230 34926 11282
rect 39442 11230 39454 11282
rect 39506 11230 39518 11282
rect 41458 11230 41470 11282
rect 41522 11230 41534 11282
rect 4958 11218 5010 11230
rect 12686 11218 12738 11230
rect 16494 11218 16546 11230
rect 20750 11218 20802 11230
rect 25902 11218 25954 11230
rect 30382 11218 30434 11230
rect 40686 11218 40738 11230
rect 42702 11218 42754 11230
rect 44830 11282 44882 11294
rect 44830 11218 44882 11230
rect 45166 11282 45218 11294
rect 45166 11218 45218 11230
rect 45726 11282 45778 11294
rect 45726 11218 45778 11230
rect 45950 11282 46002 11294
rect 45950 11218 46002 11230
rect 47182 11282 47234 11294
rect 47182 11218 47234 11230
rect 47406 11282 47458 11294
rect 53118 11282 53170 11294
rect 49074 11230 49086 11282
rect 49138 11230 49150 11282
rect 54226 11230 54238 11282
rect 54290 11230 54302 11282
rect 47406 11218 47458 11230
rect 53118 11218 53170 11230
rect 20638 11170 20690 11182
rect 20638 11106 20690 11118
rect 21310 11170 21362 11182
rect 21310 11106 21362 11118
rect 26350 11170 26402 11182
rect 26350 11106 26402 11118
rect 26686 11170 26738 11182
rect 26686 11106 26738 11118
rect 32734 11170 32786 11182
rect 32734 11106 32786 11118
rect 33070 11170 33122 11182
rect 33070 11106 33122 11118
rect 33966 11170 34018 11182
rect 33966 11106 34018 11118
rect 36430 11170 36482 11182
rect 36430 11106 36482 11118
rect 40574 11170 40626 11182
rect 40574 11106 40626 11118
rect 41918 11170 41970 11182
rect 41918 11106 41970 11118
rect 44046 11170 44098 11182
rect 44046 11106 44098 11118
rect 47518 11170 47570 11182
rect 52670 11170 52722 11182
rect 48290 11118 48302 11170
rect 48354 11118 48366 11170
rect 51426 11118 51438 11170
rect 51490 11118 51502 11170
rect 47518 11106 47570 11118
rect 52670 11106 52722 11118
rect 52782 11170 52834 11182
rect 52782 11106 52834 11118
rect 52894 11170 52946 11182
rect 52894 11106 52946 11118
rect 1344 11002 62608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 62608 11002
rect 1344 10916 62608 10950
rect 4846 10834 4898 10846
rect 4846 10770 4898 10782
rect 5182 10834 5234 10846
rect 5182 10770 5234 10782
rect 5630 10834 5682 10846
rect 5630 10770 5682 10782
rect 6078 10834 6130 10846
rect 6078 10770 6130 10782
rect 6302 10834 6354 10846
rect 6302 10770 6354 10782
rect 7758 10834 7810 10846
rect 7758 10770 7810 10782
rect 8878 10834 8930 10846
rect 8878 10770 8930 10782
rect 12462 10834 12514 10846
rect 12462 10770 12514 10782
rect 13246 10834 13298 10846
rect 13246 10770 13298 10782
rect 13470 10834 13522 10846
rect 21534 10834 21586 10846
rect 21186 10782 21198 10834
rect 21250 10782 21262 10834
rect 13470 10770 13522 10782
rect 21534 10770 21586 10782
rect 21870 10834 21922 10846
rect 21870 10770 21922 10782
rect 22094 10834 22146 10846
rect 22094 10770 22146 10782
rect 24558 10834 24610 10846
rect 24558 10770 24610 10782
rect 25230 10834 25282 10846
rect 25230 10770 25282 10782
rect 25454 10834 25506 10846
rect 25454 10770 25506 10782
rect 26350 10834 26402 10846
rect 26350 10770 26402 10782
rect 33518 10834 33570 10846
rect 33518 10770 33570 10782
rect 36094 10834 36146 10846
rect 36094 10770 36146 10782
rect 36766 10834 36818 10846
rect 36766 10770 36818 10782
rect 39790 10834 39842 10846
rect 39790 10770 39842 10782
rect 42478 10834 42530 10846
rect 46510 10834 46562 10846
rect 45154 10782 45166 10834
rect 45218 10782 45230 10834
rect 42478 10770 42530 10782
rect 46510 10770 46562 10782
rect 48078 10834 48130 10846
rect 48078 10770 48130 10782
rect 56702 10834 56754 10846
rect 56702 10770 56754 10782
rect 57150 10834 57202 10846
rect 57150 10770 57202 10782
rect 5966 10722 6018 10734
rect 5966 10658 6018 10670
rect 7422 10722 7474 10734
rect 8542 10722 8594 10734
rect 22318 10722 22370 10734
rect 8306 10670 8318 10722
rect 8370 10670 8382 10722
rect 10994 10670 11006 10722
rect 11058 10670 11070 10722
rect 16370 10670 16382 10722
rect 16434 10670 16446 10722
rect 17602 10670 17614 10722
rect 17666 10670 17678 10722
rect 18050 10670 18062 10722
rect 18114 10670 18126 10722
rect 7422 10658 7474 10670
rect 8542 10658 8594 10670
rect 22318 10658 22370 10670
rect 23214 10722 23266 10734
rect 23214 10658 23266 10670
rect 24334 10722 24386 10734
rect 24334 10658 24386 10670
rect 26462 10722 26514 10734
rect 33182 10722 33234 10734
rect 41022 10722 41074 10734
rect 27346 10670 27358 10722
rect 27410 10670 27422 10722
rect 34626 10670 34638 10722
rect 34690 10670 34702 10722
rect 37986 10670 37998 10722
rect 38050 10670 38062 10722
rect 26462 10658 26514 10670
rect 33182 10658 33234 10670
rect 41022 10658 41074 10670
rect 41694 10722 41746 10734
rect 46734 10722 46786 10734
rect 43586 10670 43598 10722
rect 43650 10670 43662 10722
rect 41694 10658 41746 10670
rect 46734 10658 46786 10670
rect 47854 10722 47906 10734
rect 47854 10658 47906 10670
rect 48190 10722 48242 10734
rect 49298 10670 49310 10722
rect 49362 10670 49374 10722
rect 53106 10670 53118 10722
rect 53170 10670 53182 10722
rect 48190 10658 48242 10670
rect 6638 10610 6690 10622
rect 8990 10610 9042 10622
rect 11678 10610 11730 10622
rect 12798 10610 12850 10622
rect 6850 10558 6862 10610
rect 6914 10558 6926 10610
rect 7970 10558 7982 10610
rect 8034 10558 8046 10610
rect 9762 10558 9774 10610
rect 9826 10558 9838 10610
rect 10210 10558 10222 10610
rect 10274 10558 10286 10610
rect 10882 10558 10894 10610
rect 10946 10558 10958 10610
rect 11890 10558 11902 10610
rect 11954 10558 11966 10610
rect 12450 10558 12462 10610
rect 12514 10558 12526 10610
rect 6638 10546 6690 10558
rect 8990 10546 9042 10558
rect 11678 10546 11730 10558
rect 12798 10546 12850 10558
rect 13022 10610 13074 10622
rect 18286 10610 18338 10622
rect 15250 10558 15262 10610
rect 15314 10558 15326 10610
rect 15474 10558 15486 10610
rect 15538 10558 15550 10610
rect 16482 10558 16494 10610
rect 16546 10558 16558 10610
rect 13022 10546 13074 10558
rect 18286 10546 18338 10558
rect 18958 10610 19010 10622
rect 18958 10546 19010 10558
rect 19518 10610 19570 10622
rect 19518 10546 19570 10558
rect 20862 10610 20914 10622
rect 20862 10546 20914 10558
rect 23550 10610 23602 10622
rect 23550 10546 23602 10558
rect 23774 10610 23826 10622
rect 33406 10610 33458 10622
rect 25666 10558 25678 10610
rect 25730 10558 25742 10610
rect 26002 10558 26014 10610
rect 26066 10558 26078 10610
rect 27010 10558 27022 10610
rect 27074 10558 27086 10610
rect 28578 10558 28590 10610
rect 28642 10558 28654 10610
rect 29922 10558 29934 10610
rect 29986 10558 29998 10610
rect 30706 10558 30718 10610
rect 30770 10558 30782 10610
rect 31490 10558 31502 10610
rect 31554 10558 31566 10610
rect 23774 10546 23826 10558
rect 33406 10546 33458 10558
rect 33630 10610 33682 10622
rect 33630 10546 33682 10558
rect 33966 10610 34018 10622
rect 34974 10610 35026 10622
rect 42030 10610 42082 10622
rect 47742 10610 47794 10622
rect 50430 10610 50482 10622
rect 54126 10610 54178 10622
rect 34178 10558 34190 10610
rect 34242 10558 34254 10610
rect 35186 10558 35198 10610
rect 35250 10558 35262 10610
rect 35970 10558 35982 10610
rect 36034 10558 36046 10610
rect 41346 10558 41358 10610
rect 41410 10558 41422 10610
rect 42242 10558 42254 10610
rect 42306 10558 42318 10610
rect 46946 10558 46958 10610
rect 47010 10558 47022 10610
rect 47282 10558 47294 10610
rect 47346 10558 47358 10610
rect 48962 10558 48974 10610
rect 49026 10558 49038 10610
rect 50642 10558 50654 10610
rect 50706 10558 50718 10610
rect 52658 10558 52670 10610
rect 52722 10558 52734 10610
rect 54338 10558 54350 10610
rect 54402 10558 54414 10610
rect 33966 10546 34018 10558
rect 34974 10546 35026 10558
rect 42030 10546 42082 10558
rect 47742 10546 47794 10558
rect 50430 10546 50482 10558
rect 54126 10546 54178 10558
rect 13358 10498 13410 10510
rect 11218 10446 11230 10498
rect 11282 10446 11294 10498
rect 13358 10434 13410 10446
rect 13918 10498 13970 10510
rect 13918 10434 13970 10446
rect 16046 10498 16098 10510
rect 21982 10498 22034 10510
rect 39230 10498 39282 10510
rect 20402 10446 20414 10498
rect 20466 10446 20478 10498
rect 24658 10446 24670 10498
rect 24722 10446 24734 10498
rect 25442 10446 25454 10498
rect 25506 10446 25518 10498
rect 28242 10446 28254 10498
rect 28306 10446 28318 10498
rect 31378 10446 31390 10498
rect 31442 10446 31454 10498
rect 16046 10434 16098 10446
rect 21982 10434 22034 10446
rect 39230 10434 39282 10446
rect 40350 10498 40402 10510
rect 40350 10434 40402 10446
rect 46622 10498 46674 10510
rect 46622 10434 46674 10446
rect 14142 10386 14194 10398
rect 18622 10386 18674 10398
rect 7970 10334 7982 10386
rect 8034 10334 8046 10386
rect 12226 10334 12238 10386
rect 12290 10334 12302 10386
rect 14466 10334 14478 10386
rect 14530 10334 14542 10386
rect 14142 10322 14194 10334
rect 18622 10322 18674 10334
rect 19182 10386 19234 10398
rect 19182 10322 19234 10334
rect 22990 10386 23042 10398
rect 22990 10322 23042 10334
rect 23102 10386 23154 10398
rect 23102 10322 23154 10334
rect 31278 10386 31330 10398
rect 31278 10322 31330 10334
rect 39342 10386 39394 10398
rect 39342 10322 39394 10334
rect 40238 10386 40290 10398
rect 40238 10322 40290 10334
rect 41358 10386 41410 10398
rect 42242 10334 42254 10386
rect 42306 10334 42318 10386
rect 48850 10334 48862 10386
rect 48914 10334 48926 10386
rect 52546 10334 52558 10386
rect 52610 10334 52622 10386
rect 41358 10322 41410 10334
rect 1344 10218 62608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 62608 10218
rect 1344 10132 62608 10166
rect 21758 10050 21810 10062
rect 5618 9998 5630 10050
rect 5682 10047 5694 10050
rect 6290 10047 6302 10050
rect 5682 10001 6302 10047
rect 5682 9998 5694 10001
rect 6290 9998 6302 10001
rect 6354 9998 6366 10050
rect 19730 9998 19742 10050
rect 19794 9998 19806 10050
rect 21758 9986 21810 9998
rect 22878 10050 22930 10062
rect 38222 10050 38274 10062
rect 50430 10050 50482 10062
rect 31042 9998 31054 10050
rect 31106 10047 31118 10050
rect 31714 10047 31726 10050
rect 31106 10001 31726 10047
rect 31106 9998 31118 10001
rect 31714 9998 31726 10001
rect 31778 9998 31790 10050
rect 47394 9998 47406 10050
rect 47458 9998 47470 10050
rect 22878 9986 22930 9998
rect 38222 9986 38274 9998
rect 50430 9986 50482 9998
rect 6302 9938 6354 9950
rect 13806 9938 13858 9950
rect 7522 9886 7534 9938
rect 7586 9886 7598 9938
rect 6302 9874 6354 9886
rect 13806 9874 13858 9886
rect 16046 9938 16098 9950
rect 31390 9938 31442 9950
rect 19170 9886 19182 9938
rect 19234 9886 19246 9938
rect 23986 9886 23998 9938
rect 24050 9886 24062 9938
rect 24994 9886 25006 9938
rect 25058 9886 25070 9938
rect 26226 9886 26238 9938
rect 26290 9886 26302 9938
rect 28018 9886 28030 9938
rect 28082 9886 28094 9938
rect 30482 9886 30494 9938
rect 30546 9886 30558 9938
rect 16046 9874 16098 9886
rect 31390 9874 31442 9886
rect 34078 9938 34130 9950
rect 34078 9874 34130 9886
rect 37886 9938 37938 9950
rect 37886 9874 37938 9886
rect 38446 9938 38498 9950
rect 38446 9874 38498 9886
rect 55582 9938 55634 9950
rect 55582 9874 55634 9886
rect 56366 9938 56418 9950
rect 56366 9874 56418 9886
rect 5966 9826 6018 9838
rect 5966 9762 6018 9774
rect 7086 9826 7138 9838
rect 7086 9762 7138 9774
rect 8318 9826 8370 9838
rect 8318 9762 8370 9774
rect 8990 9826 9042 9838
rect 14030 9826 14082 9838
rect 9762 9774 9774 9826
rect 9826 9774 9838 9826
rect 10210 9774 10222 9826
rect 10274 9774 10286 9826
rect 12002 9774 12014 9826
rect 12066 9774 12078 9826
rect 8990 9762 9042 9774
rect 14030 9762 14082 9774
rect 14702 9826 14754 9838
rect 14702 9762 14754 9774
rect 15038 9826 15090 9838
rect 25566 9826 25618 9838
rect 31950 9826 32002 9838
rect 17042 9774 17054 9826
rect 17106 9774 17118 9826
rect 17938 9774 17950 9826
rect 18002 9774 18014 9826
rect 19282 9774 19294 9826
rect 19346 9774 19358 9826
rect 23202 9774 23214 9826
rect 23266 9774 23278 9826
rect 24210 9774 24222 9826
rect 24274 9774 24286 9826
rect 25106 9774 25118 9826
rect 25170 9774 25182 9826
rect 25890 9774 25902 9826
rect 25954 9774 25966 9826
rect 28130 9774 28142 9826
rect 28194 9774 28206 9826
rect 29362 9774 29374 9826
rect 29426 9774 29438 9826
rect 30258 9774 30270 9826
rect 30322 9774 30334 9826
rect 15038 9762 15090 9774
rect 25566 9762 25618 9774
rect 31950 9762 32002 9774
rect 33966 9826 34018 9838
rect 37214 9826 37266 9838
rect 34514 9774 34526 9826
rect 34578 9774 34590 9826
rect 35410 9774 35422 9826
rect 35474 9774 35486 9826
rect 33966 9762 34018 9774
rect 37214 9762 37266 9774
rect 37662 9826 37714 9838
rect 37662 9762 37714 9774
rect 38782 9826 38834 9838
rect 38782 9762 38834 9774
rect 40126 9826 40178 9838
rect 40126 9762 40178 9774
rect 40350 9826 40402 9838
rect 40350 9762 40402 9774
rect 41582 9826 41634 9838
rect 41582 9762 41634 9774
rect 42702 9826 42754 9838
rect 45166 9826 45218 9838
rect 43586 9774 43598 9826
rect 43650 9774 43662 9826
rect 44258 9774 44270 9826
rect 44322 9774 44334 9826
rect 42702 9762 42754 9774
rect 45166 9762 45218 9774
rect 45390 9826 45442 9838
rect 51998 9826 52050 9838
rect 46386 9774 46398 9826
rect 46450 9774 46462 9826
rect 47506 9774 47518 9826
rect 47570 9774 47582 9826
rect 48402 9774 48414 9826
rect 48466 9774 48478 9826
rect 45390 9762 45442 9774
rect 51998 9762 52050 9774
rect 52782 9826 52834 9838
rect 52782 9762 52834 9774
rect 15262 9714 15314 9726
rect 21422 9714 21474 9726
rect 23438 9714 23490 9726
rect 9650 9662 9662 9714
rect 9714 9662 9726 9714
rect 10546 9662 10558 9714
rect 10610 9662 10622 9714
rect 11666 9662 11678 9714
rect 11730 9662 11742 9714
rect 18162 9662 18174 9714
rect 18226 9662 18238 9714
rect 21970 9662 21982 9714
rect 22034 9662 22046 9714
rect 22530 9662 22542 9714
rect 22594 9662 22606 9714
rect 15262 9650 15314 9662
rect 21422 9650 21474 9662
rect 23438 9650 23490 9662
rect 29822 9714 29874 9726
rect 29822 9650 29874 9662
rect 29934 9714 29986 9726
rect 35982 9714 36034 9726
rect 32946 9662 32958 9714
rect 33010 9662 33022 9714
rect 33394 9662 33406 9714
rect 33458 9662 33470 9714
rect 34962 9662 34974 9714
rect 35026 9662 35038 9714
rect 29934 9650 29986 9662
rect 35982 9650 36034 9662
rect 39118 9714 39170 9726
rect 45726 9714 45778 9726
rect 41010 9662 41022 9714
rect 41074 9662 41086 9714
rect 41346 9662 41358 9714
rect 41410 9662 41422 9714
rect 43474 9662 43486 9714
rect 43538 9662 43550 9714
rect 48850 9662 48862 9714
rect 48914 9662 48926 9714
rect 50642 9662 50654 9714
rect 50706 9662 50718 9714
rect 51202 9662 51214 9714
rect 51266 9662 51278 9714
rect 51650 9662 51662 9714
rect 51714 9662 51726 9714
rect 54002 9662 54014 9714
rect 54066 9662 54078 9714
rect 39118 9650 39170 9662
rect 45726 9650 45778 9662
rect 6862 9602 6914 9614
rect 6862 9538 6914 9550
rect 8654 9602 8706 9614
rect 14814 9602 14866 9614
rect 14354 9550 14366 9602
rect 14418 9550 14430 9602
rect 8654 9538 8706 9550
rect 14814 9538 14866 9550
rect 15710 9602 15762 9614
rect 15710 9538 15762 9550
rect 15934 9602 15986 9614
rect 15934 9538 15986 9550
rect 16158 9602 16210 9614
rect 16158 9538 16210 9550
rect 16942 9602 16994 9614
rect 16942 9538 16994 9550
rect 22990 9602 23042 9614
rect 22990 9538 23042 9550
rect 32510 9602 32562 9614
rect 36094 9602 36146 9614
rect 35522 9550 35534 9602
rect 35586 9550 35598 9602
rect 32510 9538 32562 9550
rect 36094 9538 36146 9550
rect 36990 9602 37042 9614
rect 36990 9538 37042 9550
rect 37102 9602 37154 9614
rect 37102 9538 37154 9550
rect 39678 9602 39730 9614
rect 39678 9538 39730 9550
rect 39790 9602 39842 9614
rect 39790 9538 39842 9550
rect 39902 9602 39954 9614
rect 39902 9538 39954 9550
rect 41918 9602 41970 9614
rect 41918 9538 41970 9550
rect 42478 9602 42530 9614
rect 42478 9538 42530 9550
rect 42590 9602 42642 9614
rect 45838 9602 45890 9614
rect 44146 9550 44158 9602
rect 44210 9550 44222 9602
rect 44818 9550 44830 9602
rect 44882 9550 44894 9602
rect 42590 9538 42642 9550
rect 45838 9538 45890 9550
rect 46062 9602 46114 9614
rect 46062 9538 46114 9550
rect 50094 9602 50146 9614
rect 50094 9538 50146 9550
rect 55022 9602 55074 9614
rect 55022 9538 55074 9550
rect 55918 9602 55970 9614
rect 55918 9538 55970 9550
rect 1344 9434 62608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 62608 9434
rect 1344 9348 62608 9382
rect 9998 9266 10050 9278
rect 6738 9214 6750 9266
rect 6802 9214 6814 9266
rect 9998 9202 10050 9214
rect 13022 9266 13074 9278
rect 13022 9202 13074 9214
rect 13134 9266 13186 9278
rect 25342 9266 25394 9278
rect 24098 9214 24110 9266
rect 24162 9214 24174 9266
rect 13134 9202 13186 9214
rect 25342 9202 25394 9214
rect 25566 9266 25618 9278
rect 25566 9202 25618 9214
rect 26350 9266 26402 9278
rect 26350 9202 26402 9214
rect 27246 9266 27298 9278
rect 27246 9202 27298 9214
rect 28590 9266 28642 9278
rect 28590 9202 28642 9214
rect 28814 9266 28866 9278
rect 28814 9202 28866 9214
rect 30942 9266 30994 9278
rect 30942 9202 30994 9214
rect 31278 9266 31330 9278
rect 31278 9202 31330 9214
rect 31502 9266 31554 9278
rect 31502 9202 31554 9214
rect 31614 9266 31666 9278
rect 31614 9202 31666 9214
rect 31726 9266 31778 9278
rect 31726 9202 31778 9214
rect 41806 9266 41858 9278
rect 41806 9202 41858 9214
rect 42366 9266 42418 9278
rect 42366 9202 42418 9214
rect 43598 9266 43650 9278
rect 43598 9202 43650 9214
rect 46062 9266 46114 9278
rect 46062 9202 46114 9214
rect 52782 9266 52834 9278
rect 52782 9202 52834 9214
rect 54126 9266 54178 9278
rect 54126 9202 54178 9214
rect 54574 9266 54626 9278
rect 54574 9202 54626 9214
rect 12910 9154 12962 9166
rect 17726 9154 17778 9166
rect 23662 9154 23714 9166
rect 8866 9102 8878 9154
rect 8930 9102 8942 9154
rect 11778 9102 11790 9154
rect 11842 9102 11854 9154
rect 15138 9102 15150 9154
rect 15202 9102 15214 9154
rect 16370 9102 16382 9154
rect 16434 9102 16446 9154
rect 19058 9102 19070 9154
rect 19122 9102 19134 9154
rect 12910 9090 12962 9102
rect 17726 9090 17778 9102
rect 23662 9090 23714 9102
rect 25230 9154 25282 9166
rect 29486 9154 29538 9166
rect 26898 9102 26910 9154
rect 26962 9102 26974 9154
rect 25230 9090 25282 9102
rect 29486 9090 29538 9102
rect 29710 9154 29762 9166
rect 29710 9090 29762 9102
rect 32398 9154 32450 9166
rect 34750 9154 34802 9166
rect 35646 9154 35698 9166
rect 33842 9102 33854 9154
rect 33906 9102 33918 9154
rect 35522 9102 35534 9154
rect 35586 9102 35598 9154
rect 32398 9090 32450 9102
rect 34750 9090 34802 9102
rect 35646 9090 35698 9102
rect 35758 9154 35810 9166
rect 40350 9154 40402 9166
rect 37874 9102 37886 9154
rect 37938 9102 37950 9154
rect 35758 9090 35810 9102
rect 40350 9090 40402 9102
rect 43150 9154 43202 9166
rect 48190 9154 48242 9166
rect 45490 9102 45502 9154
rect 45554 9102 45566 9154
rect 43150 9090 43202 9102
rect 48190 9090 48242 9102
rect 51438 9154 51490 9166
rect 51438 9090 51490 9102
rect 7310 9042 7362 9054
rect 7310 8978 7362 8990
rect 8094 9042 8146 9054
rect 13582 9042 13634 9054
rect 8754 8990 8766 9042
rect 8818 8990 8830 9042
rect 8094 8978 8146 8990
rect 13582 8978 13634 8990
rect 14142 9042 14194 9054
rect 17278 9042 17330 9054
rect 20974 9042 21026 9054
rect 14466 8990 14478 9042
rect 14530 8990 14542 9042
rect 15922 8990 15934 9042
rect 15986 8990 15998 9042
rect 19730 8990 19742 9042
rect 19794 8990 19806 9042
rect 14142 8978 14194 8990
rect 17278 8978 17330 8990
rect 20974 8978 21026 8990
rect 21086 9042 21138 9054
rect 23214 9042 23266 9054
rect 21634 8990 21646 9042
rect 21698 8990 21710 9042
rect 21086 8978 21138 8990
rect 23214 8978 23266 8990
rect 23438 9042 23490 9054
rect 26574 9042 26626 9054
rect 25890 8990 25902 9042
rect 25954 8990 25966 9042
rect 26114 8990 26126 9042
rect 26178 8990 26190 9042
rect 23438 8978 23490 8990
rect 26574 8978 26626 8990
rect 27694 9042 27746 9054
rect 27694 8978 27746 8990
rect 28030 9042 28082 9054
rect 28030 8978 28082 8990
rect 28366 9042 28418 9054
rect 28366 8978 28418 8990
rect 28702 9042 28754 9054
rect 28702 8978 28754 8990
rect 29262 9042 29314 9054
rect 29262 8978 29314 8990
rect 32286 9042 32338 9054
rect 32286 8978 32338 8990
rect 32622 9042 32674 9054
rect 34862 9042 34914 9054
rect 33394 8990 33406 9042
rect 33458 8990 33470 9042
rect 33954 8990 33966 9042
rect 34018 8990 34030 9042
rect 32622 8978 32674 8990
rect 34862 8978 34914 8990
rect 35982 9042 36034 9054
rect 38558 9042 38610 9054
rect 36530 8990 36542 9042
rect 36594 8990 36606 9042
rect 37762 8990 37774 9042
rect 37826 8990 37838 9042
rect 35982 8978 36034 8990
rect 38558 8978 38610 8990
rect 38894 9042 38946 9054
rect 38894 8978 38946 8990
rect 39118 9042 39170 9054
rect 39118 8978 39170 8990
rect 40126 9042 40178 9054
rect 40126 8978 40178 8990
rect 41022 9042 41074 9054
rect 41022 8978 41074 8990
rect 41470 9042 41522 9054
rect 41470 8978 41522 8990
rect 41694 9042 41746 9054
rect 42702 9042 42754 9054
rect 46286 9042 46338 9054
rect 42354 8990 42366 9042
rect 42418 8990 42430 9042
rect 42914 8990 42926 9042
rect 42978 8990 42990 9042
rect 44146 8990 44158 9042
rect 44210 8990 44222 9042
rect 44482 8990 44494 9042
rect 44546 8990 44558 9042
rect 45602 8990 45614 9042
rect 45666 8990 45678 9042
rect 41694 8978 41746 8990
rect 42702 8978 42754 8990
rect 46286 8978 46338 8990
rect 46734 9042 46786 9054
rect 48738 8990 48750 9042
rect 48802 8990 48814 9042
rect 49410 8990 49422 9042
rect 49474 8990 49486 9042
rect 51650 8990 51662 9042
rect 51714 8990 51726 9042
rect 52658 8990 52670 9042
rect 52722 8990 52734 9042
rect 46734 8978 46786 8990
rect 7086 8930 7138 8942
rect 7086 8866 7138 8878
rect 10446 8930 10498 8942
rect 23326 8930 23378 8942
rect 18834 8878 18846 8930
rect 18898 8878 18910 8930
rect 21746 8878 21758 8930
rect 21810 8878 21822 8930
rect 10446 8866 10498 8878
rect 23326 8866 23378 8878
rect 24670 8930 24722 8942
rect 28142 8930 28194 8942
rect 30270 8930 30322 8942
rect 35870 8930 35922 8942
rect 39006 8930 39058 8942
rect 26226 8878 26238 8930
rect 26290 8878 26302 8930
rect 29810 8878 29822 8930
rect 29874 8878 29886 8930
rect 33618 8878 33630 8930
rect 33682 8878 33694 8930
rect 36866 8878 36878 8930
rect 36930 8878 36942 8930
rect 24670 8866 24722 8878
rect 28142 8866 28194 8878
rect 30270 8866 30322 8878
rect 35870 8866 35922 8878
rect 39006 8866 39058 8878
rect 39566 8930 39618 8942
rect 39566 8866 39618 8878
rect 44942 8930 44994 8942
rect 49646 8930 49698 8942
rect 47842 8878 47854 8930
rect 47906 8878 47918 8930
rect 44942 8866 44994 8878
rect 49646 8866 49698 8878
rect 53678 8930 53730 8942
rect 53678 8866 53730 8878
rect 7758 8818 7810 8830
rect 24446 8818 24498 8830
rect 18722 8766 18734 8818
rect 18786 8766 18798 8818
rect 7758 8754 7810 8766
rect 24446 8754 24498 8766
rect 30046 8818 30098 8830
rect 30046 8754 30098 8766
rect 34750 8818 34802 8830
rect 39790 8818 39842 8830
rect 36978 8766 36990 8818
rect 37042 8766 37054 8818
rect 34750 8754 34802 8766
rect 39790 8754 39842 8766
rect 40238 8818 40290 8830
rect 40238 8754 40290 8766
rect 40910 8818 40962 8830
rect 47954 8766 47966 8818
rect 48018 8766 48030 8818
rect 40910 8754 40962 8766
rect 1344 8650 62608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 62608 8650
rect 1344 8564 62608 8598
rect 18162 8430 18174 8482
rect 18226 8430 18238 8482
rect 47730 8430 47742 8482
rect 47794 8430 47806 8482
rect 8318 8370 8370 8382
rect 8318 8306 8370 8318
rect 20302 8370 20354 8382
rect 51438 8370 51490 8382
rect 22082 8318 22094 8370
rect 22146 8318 22158 8370
rect 24210 8318 24222 8370
rect 24274 8318 24286 8370
rect 29922 8318 29934 8370
rect 29986 8318 29998 8370
rect 32050 8318 32062 8370
rect 32114 8318 32126 8370
rect 37202 8318 37214 8370
rect 37266 8318 37278 8370
rect 37986 8318 37998 8370
rect 38050 8318 38062 8370
rect 39890 8318 39902 8370
rect 39954 8318 39966 8370
rect 43138 8318 43150 8370
rect 43202 8318 43214 8370
rect 20302 8306 20354 8318
rect 51438 8306 51490 8318
rect 51998 8370 52050 8382
rect 51998 8306 52050 8318
rect 52894 8370 52946 8382
rect 52894 8306 52946 8318
rect 53342 8370 53394 8382
rect 53342 8306 53394 8318
rect 53790 8370 53842 8382
rect 53790 8306 53842 8318
rect 7758 8258 7810 8270
rect 7758 8194 7810 8206
rect 8206 8258 8258 8270
rect 8206 8194 8258 8206
rect 11006 8258 11058 8270
rect 11006 8194 11058 8206
rect 12462 8258 12514 8270
rect 12462 8194 12514 8206
rect 12798 8258 12850 8270
rect 19854 8258 19906 8270
rect 16258 8206 16270 8258
rect 16322 8206 16334 8258
rect 17378 8206 17390 8258
rect 17442 8206 17454 8258
rect 19282 8206 19294 8258
rect 19346 8206 19358 8258
rect 12798 8194 12850 8206
rect 19854 8194 19906 8206
rect 20078 8258 20130 8270
rect 20078 8194 20130 8206
rect 20414 8258 20466 8270
rect 24782 8258 24834 8270
rect 21410 8206 21422 8258
rect 21474 8206 21486 8258
rect 20414 8194 20466 8206
rect 24782 8194 24834 8206
rect 27134 8258 27186 8270
rect 27134 8194 27186 8206
rect 27358 8258 27410 8270
rect 27358 8194 27410 8206
rect 28590 8258 28642 8270
rect 33294 8258 33346 8270
rect 29138 8206 29150 8258
rect 29202 8206 29214 8258
rect 28590 8194 28642 8206
rect 33294 8194 33346 8206
rect 33966 8258 34018 8270
rect 33966 8194 34018 8206
rect 34414 8258 34466 8270
rect 34414 8194 34466 8206
rect 35982 8258 36034 8270
rect 35982 8194 36034 8206
rect 36990 8258 37042 8270
rect 46510 8258 46562 8270
rect 37314 8206 37326 8258
rect 37378 8206 37390 8258
rect 38098 8206 38110 8258
rect 38162 8206 38174 8258
rect 38994 8206 39006 8258
rect 39058 8206 39070 8258
rect 40226 8206 40238 8258
rect 40290 8206 40302 8258
rect 42354 8206 42366 8258
rect 42418 8206 42430 8258
rect 43586 8206 43598 8258
rect 43650 8206 43662 8258
rect 45042 8206 45054 8258
rect 45106 8206 45118 8258
rect 46946 8206 46958 8258
rect 47010 8206 47022 8258
rect 48514 8206 48526 8258
rect 48578 8206 48590 8258
rect 48850 8206 48862 8258
rect 48914 8206 48926 8258
rect 36990 8194 37042 8206
rect 46510 8194 46562 8206
rect 49086 8202 49138 8214
rect 8430 8146 8482 8158
rect 34638 8146 34690 8158
rect 41022 8146 41074 8158
rect 9090 8094 9102 8146
rect 9154 8094 9166 8146
rect 11778 8094 11790 8146
rect 11842 8094 11854 8146
rect 12226 8094 12238 8146
rect 12290 8094 12302 8146
rect 18610 8094 18622 8146
rect 18674 8094 18686 8146
rect 32610 8094 32622 8146
rect 32674 8094 32686 8146
rect 32946 8094 32958 8146
rect 33010 8094 33022 8146
rect 35410 8094 35422 8146
rect 35474 8094 35486 8146
rect 35746 8094 35758 8146
rect 35810 8094 35822 8146
rect 39106 8094 39118 8146
rect 39170 8094 39182 8146
rect 39778 8094 39790 8146
rect 39842 8094 39854 8146
rect 42018 8094 42030 8146
rect 42082 8094 42094 8146
rect 45378 8094 45390 8146
rect 45442 8094 45454 8146
rect 49086 8138 49138 8150
rect 8430 8082 8482 8094
rect 34638 8082 34690 8094
rect 41022 8082 41074 8094
rect 15262 8034 15314 8046
rect 14130 7982 14142 8034
rect 14194 7982 14206 8034
rect 15262 7970 15314 7982
rect 15934 8034 15986 8046
rect 28366 8034 28418 8046
rect 26114 7982 26126 8034
rect 26178 7982 26190 8034
rect 27682 7982 27694 8034
rect 27746 7982 27758 8034
rect 15934 7970 15986 7982
rect 28366 7970 28418 7982
rect 28478 8034 28530 8046
rect 28478 7970 28530 7982
rect 33630 8034 33682 8046
rect 33630 7970 33682 7982
rect 34302 8034 34354 8046
rect 34302 7970 34354 7982
rect 36318 8034 36370 8046
rect 36318 7970 36370 7982
rect 41358 8034 41410 8046
rect 41358 7970 41410 7982
rect 49198 8034 49250 8046
rect 49198 7970 49250 7982
rect 49310 8034 49362 8046
rect 54126 8034 54178 8046
rect 50306 7982 50318 8034
rect 50370 7982 50382 8034
rect 49310 7970 49362 7982
rect 54126 7970 54178 7982
rect 1344 7866 62608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 62608 7866
rect 1344 7780 62608 7814
rect 8318 7698 8370 7710
rect 8318 7634 8370 7646
rect 8542 7698 8594 7710
rect 8542 7634 8594 7646
rect 9998 7698 10050 7710
rect 9998 7634 10050 7646
rect 16046 7698 16098 7710
rect 16046 7634 16098 7646
rect 16718 7698 16770 7710
rect 16718 7634 16770 7646
rect 20414 7698 20466 7710
rect 20414 7634 20466 7646
rect 20638 7698 20690 7710
rect 31166 7698 31218 7710
rect 28018 7646 28030 7698
rect 28082 7646 28094 7698
rect 30034 7646 30046 7698
rect 30098 7646 30110 7698
rect 20638 7634 20690 7646
rect 31166 7634 31218 7646
rect 41358 7698 41410 7710
rect 41358 7634 41410 7646
rect 41470 7698 41522 7710
rect 41470 7634 41522 7646
rect 42366 7698 42418 7710
rect 42366 7634 42418 7646
rect 43710 7698 43762 7710
rect 43710 7634 43762 7646
rect 44382 7698 44434 7710
rect 44382 7634 44434 7646
rect 44606 7698 44658 7710
rect 44606 7634 44658 7646
rect 45166 7698 45218 7710
rect 45166 7634 45218 7646
rect 46734 7698 46786 7710
rect 48078 7698 48130 7710
rect 47170 7646 47182 7698
rect 47234 7646 47246 7698
rect 46734 7634 46786 7646
rect 48078 7634 48130 7646
rect 51662 7698 51714 7710
rect 51662 7634 51714 7646
rect 52110 7698 52162 7710
rect 52110 7634 52162 7646
rect 8206 7586 8258 7598
rect 16606 7586 16658 7598
rect 20302 7586 20354 7598
rect 28478 7586 28530 7598
rect 10882 7534 10894 7586
rect 10946 7534 10958 7586
rect 13458 7534 13470 7586
rect 13522 7534 13534 7586
rect 18722 7534 18734 7586
rect 18786 7534 18798 7586
rect 20066 7534 20078 7586
rect 20130 7534 20142 7586
rect 25666 7534 25678 7586
rect 25730 7534 25742 7586
rect 8206 7522 8258 7534
rect 16606 7522 16658 7534
rect 20302 7522 20354 7534
rect 28478 7522 28530 7534
rect 28814 7586 28866 7598
rect 28814 7522 28866 7534
rect 29150 7586 29202 7598
rect 30830 7586 30882 7598
rect 39230 7586 39282 7598
rect 29922 7534 29934 7586
rect 29986 7534 29998 7586
rect 33170 7534 33182 7586
rect 33234 7534 33246 7586
rect 29150 7522 29202 7534
rect 30830 7522 30882 7534
rect 39230 7522 39282 7534
rect 39342 7586 39394 7598
rect 39342 7522 39394 7534
rect 43374 7586 43426 7598
rect 43374 7522 43426 7534
rect 43486 7586 43538 7598
rect 43486 7522 43538 7534
rect 44158 7586 44210 7598
rect 44158 7522 44210 7534
rect 44494 7586 44546 7598
rect 45826 7534 45838 7586
rect 45890 7534 45902 7586
rect 49970 7534 49982 7586
rect 50034 7534 50046 7586
rect 44494 7522 44546 7534
rect 22430 7474 22482 7486
rect 29374 7474 29426 7486
rect 12674 7422 12686 7474
rect 12738 7422 12750 7474
rect 15922 7422 15934 7474
rect 15986 7422 15998 7474
rect 21634 7422 21646 7474
rect 21698 7422 21710 7474
rect 22866 7422 22878 7474
rect 22930 7422 22942 7474
rect 27794 7422 27806 7474
rect 27858 7422 27870 7474
rect 22430 7410 22482 7422
rect 29374 7410 29426 7422
rect 29710 7474 29762 7486
rect 31054 7474 31106 7486
rect 30482 7422 30494 7474
rect 30546 7422 30558 7474
rect 29710 7410 29762 7422
rect 31054 7410 31106 7422
rect 31502 7474 31554 7486
rect 31502 7410 31554 7422
rect 32510 7474 32562 7486
rect 36318 7474 36370 7486
rect 33506 7422 33518 7474
rect 33570 7422 33582 7474
rect 34066 7422 34078 7474
rect 34130 7422 34142 7474
rect 34514 7422 34526 7474
rect 34578 7422 34590 7474
rect 35522 7422 35534 7474
rect 35586 7422 35598 7474
rect 32510 7410 32562 7422
rect 36318 7410 36370 7422
rect 38110 7474 38162 7486
rect 39566 7474 39618 7486
rect 38770 7422 38782 7474
rect 38834 7422 38846 7474
rect 38110 7410 38162 7422
rect 39566 7410 39618 7422
rect 40798 7474 40850 7486
rect 40798 7410 40850 7422
rect 41246 7474 41298 7486
rect 46398 7474 46450 7486
rect 42914 7422 42926 7474
rect 42978 7422 42990 7474
rect 45602 7422 45614 7474
rect 45666 7422 45678 7474
rect 47394 7422 47406 7474
rect 47458 7422 47470 7474
rect 41246 7410 41298 7422
rect 46398 7410 46450 7422
rect 28926 7362 28978 7374
rect 40350 7362 40402 7374
rect 48190 7362 48242 7374
rect 15586 7310 15598 7362
rect 15650 7310 15662 7362
rect 20290 7310 20302 7362
rect 20354 7310 20366 7362
rect 23202 7310 23214 7362
rect 23266 7310 23278 7362
rect 32050 7310 32062 7362
rect 32114 7310 32126 7362
rect 33170 7310 33182 7362
rect 33234 7310 33246 7362
rect 35410 7310 35422 7362
rect 35474 7310 35486 7362
rect 41906 7310 41918 7362
rect 41970 7310 41982 7362
rect 43362 7310 43374 7362
rect 43426 7310 43438 7362
rect 28926 7298 28978 7310
rect 40350 7298 40402 7310
rect 48190 7298 48242 7310
rect 48862 7362 48914 7374
rect 48862 7298 48914 7310
rect 51102 7362 51154 7374
rect 51102 7298 51154 7310
rect 52446 7362 52498 7374
rect 52446 7298 52498 7310
rect 52894 7362 52946 7374
rect 52894 7298 52946 7310
rect 12238 7250 12290 7262
rect 12238 7186 12290 7198
rect 16718 7250 16770 7262
rect 16718 7186 16770 7198
rect 17502 7250 17554 7262
rect 27470 7250 27522 7262
rect 39790 7250 39842 7262
rect 21074 7198 21086 7250
rect 21138 7198 21150 7250
rect 30258 7198 30270 7250
rect 30322 7198 30334 7250
rect 17502 7186 17554 7198
rect 27470 7186 27522 7198
rect 39790 7186 39842 7198
rect 40126 7250 40178 7262
rect 40126 7186 40178 7198
rect 1344 7082 62608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 62608 7082
rect 1344 6996 62608 7030
rect 10558 6914 10610 6926
rect 10558 6850 10610 6862
rect 23102 6914 23154 6926
rect 23102 6850 23154 6862
rect 26462 6914 26514 6926
rect 26462 6850 26514 6862
rect 26798 6914 26850 6926
rect 31614 6914 31666 6926
rect 42590 6914 42642 6926
rect 30034 6862 30046 6914
rect 30098 6862 30110 6914
rect 33282 6862 33294 6914
rect 33346 6862 33358 6914
rect 26798 6850 26850 6862
rect 31614 6850 31666 6862
rect 42590 6850 42642 6862
rect 45390 6914 45442 6926
rect 45390 6850 45442 6862
rect 10894 6802 10946 6814
rect 28478 6802 28530 6814
rect 45054 6802 45106 6814
rect 20514 6750 20526 6802
rect 20578 6750 20590 6802
rect 22194 6750 22206 6802
rect 22258 6750 22270 6802
rect 32162 6750 32174 6802
rect 32226 6750 32238 6802
rect 33618 6750 33630 6802
rect 33682 6750 33694 6802
rect 35746 6750 35758 6802
rect 35810 6750 35822 6802
rect 10894 6738 10946 6750
rect 28478 6738 28530 6750
rect 45054 6738 45106 6750
rect 45838 6802 45890 6814
rect 49522 6750 49534 6802
rect 49586 6750 49598 6802
rect 45838 6738 45890 6750
rect 9550 6690 9602 6702
rect 9550 6626 9602 6638
rect 9662 6690 9714 6702
rect 9662 6626 9714 6638
rect 9774 6690 9826 6702
rect 9774 6626 9826 6638
rect 10110 6690 10162 6702
rect 12462 6690 12514 6702
rect 11666 6638 11678 6690
rect 11730 6638 11742 6690
rect 10110 6626 10162 6638
rect 12462 6626 12514 6638
rect 13022 6690 13074 6702
rect 13022 6626 13074 6638
rect 13470 6690 13522 6702
rect 13470 6626 13522 6638
rect 14702 6690 14754 6702
rect 14702 6626 14754 6638
rect 15822 6690 15874 6702
rect 15822 6626 15874 6638
rect 16270 6690 16322 6702
rect 16270 6626 16322 6638
rect 16606 6690 16658 6702
rect 16606 6626 16658 6638
rect 16942 6690 16994 6702
rect 21646 6690 21698 6702
rect 20178 6638 20190 6690
rect 20242 6638 20254 6690
rect 16942 6626 16994 6638
rect 21646 6626 21698 6638
rect 24334 6690 24386 6702
rect 24334 6626 24386 6638
rect 24670 6690 24722 6702
rect 29822 6690 29874 6702
rect 32622 6690 32674 6702
rect 45726 6690 45778 6702
rect 27234 6638 27246 6690
rect 27298 6638 27310 6690
rect 30034 6638 30046 6690
rect 30098 6638 30110 6690
rect 33506 6638 33518 6690
rect 33570 6638 33582 6690
rect 34290 6638 34302 6690
rect 34354 6638 34366 6690
rect 37538 6638 37550 6690
rect 37602 6638 37614 6690
rect 43250 6638 43262 6690
rect 43314 6638 43326 6690
rect 44258 6638 44270 6690
rect 44322 6638 44334 6690
rect 24670 6626 24722 6638
rect 29822 6626 29874 6638
rect 32622 6626 32674 6638
rect 45726 6626 45778 6638
rect 45950 6690 46002 6702
rect 45950 6626 46002 6638
rect 47518 6690 47570 6702
rect 47518 6626 47570 6638
rect 48414 6690 48466 6702
rect 48414 6626 48466 6638
rect 49086 6690 49138 6702
rect 49086 6626 49138 6638
rect 50318 6690 50370 6702
rect 50318 6626 50370 6638
rect 50766 6690 50818 6702
rect 50766 6626 50818 6638
rect 51214 6690 51266 6702
rect 51214 6626 51266 6638
rect 51662 6690 51714 6702
rect 51662 6626 51714 6638
rect 13806 6578 13858 6590
rect 11554 6526 11566 6578
rect 11618 6526 11630 6578
rect 13806 6514 13858 6526
rect 14366 6578 14418 6590
rect 14366 6514 14418 6526
rect 15374 6578 15426 6590
rect 19630 6578 19682 6590
rect 18498 6526 18510 6578
rect 18562 6526 18574 6578
rect 15374 6514 15426 6526
rect 19630 6514 19682 6526
rect 21310 6578 21362 6590
rect 21310 6514 21362 6526
rect 21982 6578 22034 6590
rect 21982 6514 22034 6526
rect 23102 6578 23154 6590
rect 23102 6514 23154 6526
rect 23214 6578 23266 6590
rect 23214 6514 23266 6526
rect 25006 6578 25058 6590
rect 25006 6514 25058 6526
rect 25342 6578 25394 6590
rect 25342 6514 25394 6526
rect 25678 6578 25730 6590
rect 25678 6514 25730 6526
rect 26014 6578 26066 6590
rect 28254 6578 28306 6590
rect 27570 6526 27582 6578
rect 27634 6526 27646 6578
rect 26014 6514 26066 6526
rect 28254 6514 28306 6526
rect 29486 6578 29538 6590
rect 29486 6514 29538 6526
rect 29598 6578 29650 6590
rect 31726 6578 31778 6590
rect 35198 6578 35250 6590
rect 30930 6526 30942 6578
rect 30994 6526 31006 6578
rect 34514 6526 34526 6578
rect 34578 6526 34590 6578
rect 29598 6514 29650 6526
rect 31726 6514 31778 6526
rect 35198 6514 35250 6526
rect 35310 6578 35362 6590
rect 36430 6578 36482 6590
rect 42702 6578 42754 6590
rect 44830 6578 44882 6590
rect 35410 6526 35422 6578
rect 35474 6526 35486 6578
rect 39218 6526 39230 6578
rect 39282 6526 39294 6578
rect 41794 6526 41806 6578
rect 41858 6526 41870 6578
rect 44146 6526 44158 6578
rect 44210 6526 44222 6578
rect 35310 6514 35362 6526
rect 36430 6514 36482 6526
rect 42702 6514 42754 6526
rect 44830 6514 44882 6526
rect 46174 6578 46226 6590
rect 48638 6578 48690 6590
rect 47842 6526 47854 6578
rect 47906 6526 47918 6578
rect 46174 6514 46226 6526
rect 48638 6514 48690 6526
rect 48750 6578 48802 6590
rect 49970 6526 49982 6578
rect 50034 6526 50046 6578
rect 48750 6514 48802 6526
rect 16718 6466 16770 6478
rect 16718 6402 16770 6414
rect 17502 6466 17554 6478
rect 17502 6402 17554 6414
rect 23774 6466 23826 6478
rect 23774 6402 23826 6414
rect 25230 6466 25282 6478
rect 25230 6402 25282 6414
rect 28366 6466 28418 6478
rect 28366 6402 28418 6414
rect 31278 6466 31330 6478
rect 31278 6402 31330 6414
rect 34974 6466 35026 6478
rect 34974 6402 35026 6414
rect 36318 6466 36370 6478
rect 36318 6402 36370 6414
rect 40014 6466 40066 6478
rect 47070 6466 47122 6478
rect 43250 6414 43262 6466
rect 43314 6414 43326 6466
rect 40014 6402 40066 6414
rect 47070 6402 47122 6414
rect 47294 6466 47346 6478
rect 47294 6402 47346 6414
rect 47406 6466 47458 6478
rect 47406 6402 47458 6414
rect 48190 6466 48242 6478
rect 48190 6402 48242 6414
rect 52110 6466 52162 6478
rect 52110 6402 52162 6414
rect 1344 6298 62608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 62608 6298
rect 1344 6212 62608 6246
rect 12462 6130 12514 6142
rect 12462 6066 12514 6078
rect 13246 6130 13298 6142
rect 13246 6066 13298 6078
rect 13470 6130 13522 6142
rect 13470 6066 13522 6078
rect 14478 6130 14530 6142
rect 14478 6066 14530 6078
rect 14926 6130 14978 6142
rect 14926 6066 14978 6078
rect 15374 6130 15426 6142
rect 15374 6066 15426 6078
rect 15822 6130 15874 6142
rect 15822 6066 15874 6078
rect 16830 6130 16882 6142
rect 16830 6066 16882 6078
rect 17502 6130 17554 6142
rect 20414 6130 20466 6142
rect 18834 6078 18846 6130
rect 18898 6078 18910 6130
rect 17502 6066 17554 6078
rect 20414 6066 20466 6078
rect 20974 6130 21026 6142
rect 20974 6066 21026 6078
rect 21422 6130 21474 6142
rect 21422 6066 21474 6078
rect 21982 6130 22034 6142
rect 21982 6066 22034 6078
rect 22990 6130 23042 6142
rect 22990 6066 23042 6078
rect 23438 6130 23490 6142
rect 23438 6066 23490 6078
rect 24334 6130 24386 6142
rect 24334 6066 24386 6078
rect 24782 6130 24834 6142
rect 24782 6066 24834 6078
rect 25454 6130 25506 6142
rect 29934 6130 29986 6142
rect 35422 6130 35474 6142
rect 26338 6078 26350 6130
rect 26402 6078 26414 6130
rect 31602 6078 31614 6130
rect 31666 6078 31678 6130
rect 25454 6066 25506 6078
rect 29934 6066 29986 6078
rect 35422 6066 35474 6078
rect 39566 6130 39618 6142
rect 39566 6066 39618 6078
rect 39790 6130 39842 6142
rect 44942 6130 44994 6142
rect 47182 6130 47234 6142
rect 42466 6078 42478 6130
rect 42530 6078 42542 6130
rect 45266 6078 45278 6130
rect 45330 6078 45342 6130
rect 39790 6066 39842 6078
rect 44942 6066 44994 6078
rect 47182 6066 47234 6078
rect 47630 6130 47682 6142
rect 47630 6066 47682 6078
rect 48862 6130 48914 6142
rect 48862 6066 48914 6078
rect 49086 6130 49138 6142
rect 49086 6066 49138 6078
rect 49422 6130 49474 6142
rect 49422 6066 49474 6078
rect 49982 6130 50034 6142
rect 49982 6066 50034 6078
rect 50318 6130 50370 6142
rect 50318 6066 50370 6078
rect 13806 6018 13858 6030
rect 31054 6018 31106 6030
rect 28130 5966 28142 6018
rect 28194 5966 28206 6018
rect 13806 5954 13858 5966
rect 31054 5954 31106 5966
rect 34078 6018 34130 6030
rect 34078 5954 34130 5966
rect 35086 6018 35138 6030
rect 35086 5954 35138 5966
rect 35198 6018 35250 6030
rect 35198 5954 35250 5966
rect 41582 6018 41634 6030
rect 46958 6018 47010 6030
rect 43250 5966 43262 6018
rect 43314 5966 43326 6018
rect 41582 5954 41634 5966
rect 46958 5954 47010 5966
rect 47966 6018 48018 6030
rect 47966 5954 48018 5966
rect 48078 6018 48130 6030
rect 48078 5954 48130 5966
rect 48750 6018 48802 6030
rect 48750 5954 48802 5966
rect 19854 5906 19906 5918
rect 19854 5842 19906 5854
rect 22430 5906 22482 5918
rect 22430 5842 22482 5854
rect 27470 5906 27522 5918
rect 28814 5906 28866 5918
rect 28018 5854 28030 5906
rect 28082 5854 28094 5906
rect 27470 5842 27522 5854
rect 28814 5842 28866 5854
rect 30158 5906 30210 5918
rect 30158 5842 30210 5854
rect 31278 5906 31330 5918
rect 31278 5842 31330 5854
rect 32510 5906 32562 5918
rect 32510 5842 32562 5854
rect 33070 5906 33122 5918
rect 38446 5906 38498 5918
rect 33282 5854 33294 5906
rect 33346 5854 33358 5906
rect 34290 5854 34302 5906
rect 34354 5854 34366 5906
rect 35634 5854 35646 5906
rect 35698 5854 35710 5906
rect 33070 5842 33122 5854
rect 38446 5842 38498 5854
rect 38782 5906 38834 5918
rect 41918 5906 41970 5918
rect 40114 5854 40126 5906
rect 40178 5854 40190 5906
rect 41346 5854 41358 5906
rect 41410 5854 41422 5906
rect 38782 5842 38834 5854
rect 41918 5842 41970 5854
rect 42142 5906 42194 5918
rect 42142 5842 42194 5854
rect 45614 5906 45666 5918
rect 45614 5842 45666 5854
rect 45838 5906 45890 5918
rect 45838 5842 45890 5854
rect 46174 5906 46226 5918
rect 46174 5842 46226 5854
rect 46846 5906 46898 5918
rect 46846 5842 46898 5854
rect 16382 5794 16434 5806
rect 16382 5730 16434 5742
rect 29150 5794 29202 5806
rect 39678 5794 39730 5806
rect 50766 5794 50818 5806
rect 32050 5742 32062 5794
rect 32114 5742 32126 5794
rect 34514 5742 34526 5794
rect 34578 5742 34590 5794
rect 36082 5742 36094 5794
rect 36146 5742 36158 5794
rect 38210 5742 38222 5794
rect 38274 5742 38286 5794
rect 46386 5742 46398 5794
rect 46450 5742 46462 5794
rect 29150 5730 29202 5742
rect 39678 5730 39730 5742
rect 50766 5730 50818 5742
rect 30382 5682 30434 5694
rect 22418 5630 22430 5682
rect 22482 5679 22494 5682
rect 23314 5679 23326 5682
rect 22482 5633 23326 5679
rect 22482 5630 22494 5633
rect 23314 5630 23326 5633
rect 23378 5630 23390 5682
rect 24098 5630 24110 5682
rect 24162 5679 24174 5682
rect 24770 5679 24782 5682
rect 24162 5633 24782 5679
rect 24162 5630 24174 5633
rect 24770 5630 24782 5633
rect 24834 5630 24846 5682
rect 30706 5630 30718 5682
rect 30770 5630 30782 5682
rect 49634 5630 49646 5682
rect 49698 5679 49710 5682
rect 50194 5679 50206 5682
rect 49698 5633 50206 5679
rect 49698 5630 49710 5633
rect 50194 5630 50206 5633
rect 50258 5630 50270 5682
rect 30382 5618 30434 5630
rect 1344 5514 62608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 62608 5514
rect 1344 5428 62608 5462
rect 31390 5346 31442 5358
rect 24098 5294 24110 5346
rect 24162 5343 24174 5346
rect 25106 5343 25118 5346
rect 24162 5297 25118 5343
rect 24162 5294 24174 5297
rect 25106 5294 25118 5297
rect 25170 5294 25182 5346
rect 25666 5294 25678 5346
rect 25730 5343 25742 5346
rect 26786 5343 26798 5346
rect 25730 5297 26798 5343
rect 25730 5294 25742 5297
rect 26786 5294 26798 5297
rect 26850 5294 26862 5346
rect 31390 5282 31442 5294
rect 31726 5346 31778 5358
rect 31726 5282 31778 5294
rect 35646 5346 35698 5358
rect 35646 5282 35698 5294
rect 35982 5346 36034 5358
rect 35982 5282 36034 5294
rect 40574 5346 40626 5358
rect 40574 5282 40626 5294
rect 45726 5346 45778 5358
rect 45726 5282 45778 5294
rect 46062 5346 46114 5358
rect 46062 5282 46114 5294
rect 13806 5234 13858 5246
rect 13806 5170 13858 5182
rect 16046 5234 16098 5246
rect 16046 5170 16098 5182
rect 16382 5234 16434 5246
rect 16382 5170 16434 5182
rect 18846 5234 18898 5246
rect 18846 5170 18898 5182
rect 19406 5234 19458 5246
rect 19406 5170 19458 5182
rect 19966 5234 20018 5246
rect 19966 5170 20018 5182
rect 20302 5234 20354 5246
rect 20302 5170 20354 5182
rect 20862 5234 20914 5246
rect 20862 5170 20914 5182
rect 21870 5234 21922 5246
rect 21870 5170 21922 5182
rect 22430 5234 22482 5246
rect 22430 5170 22482 5182
rect 22990 5234 23042 5246
rect 22990 5170 23042 5182
rect 23662 5234 23714 5246
rect 23662 5170 23714 5182
rect 24110 5234 24162 5246
rect 24110 5170 24162 5182
rect 24670 5234 24722 5246
rect 24670 5170 24722 5182
rect 25006 5234 25058 5246
rect 25006 5170 25058 5182
rect 25678 5234 25730 5246
rect 25678 5170 25730 5182
rect 26574 5234 26626 5246
rect 26574 5170 26626 5182
rect 27134 5234 27186 5246
rect 27134 5170 27186 5182
rect 31614 5234 31666 5246
rect 43038 5234 43090 5246
rect 36978 5182 36990 5234
rect 37042 5182 37054 5234
rect 39106 5182 39118 5234
rect 39170 5182 39182 5234
rect 47506 5182 47518 5234
rect 47570 5182 47582 5234
rect 49634 5182 49646 5234
rect 49698 5182 49710 5234
rect 31614 5170 31666 5182
rect 43038 5170 43090 5182
rect 15486 5122 15538 5134
rect 15486 5058 15538 5070
rect 16942 5122 16994 5134
rect 16942 5058 16994 5070
rect 27694 5122 27746 5134
rect 43374 5122 43426 5134
rect 50206 5122 50258 5134
rect 28242 5070 28254 5122
rect 28306 5070 28318 5122
rect 32050 5070 32062 5122
rect 32114 5070 32126 5122
rect 33058 5070 33070 5122
rect 33122 5070 33134 5122
rect 33954 5070 33966 5122
rect 34018 5070 34030 5122
rect 34962 5070 34974 5122
rect 35026 5070 35038 5122
rect 39890 5070 39902 5122
rect 39954 5070 39966 5122
rect 43810 5070 43822 5122
rect 43874 5070 43886 5122
rect 45042 5070 45054 5122
rect 45106 5070 45118 5122
rect 46834 5070 46846 5122
rect 46898 5070 46910 5122
rect 27694 5058 27746 5070
rect 43374 5058 43426 5070
rect 50206 5058 50258 5070
rect 28030 5010 28082 5022
rect 27346 4958 27358 5010
rect 27410 4958 27422 5010
rect 29586 4958 29598 5010
rect 29650 4958 29662 5010
rect 32162 4958 32174 5010
rect 32226 4958 32238 5010
rect 34850 4958 34862 5010
rect 34914 4958 34926 5010
rect 42018 4958 42030 5010
rect 42082 4958 42094 5010
rect 44146 4958 44158 5010
rect 44210 4958 44222 5010
rect 44930 4958 44942 5010
rect 44994 4958 45006 5010
rect 28030 4946 28082 4958
rect 21534 4898 21586 4910
rect 21534 4834 21586 4846
rect 26126 4898 26178 4910
rect 26126 4834 26178 4846
rect 1344 4730 62608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 62608 4730
rect 1344 4644 62608 4678
rect 21086 4562 21138 4574
rect 21086 4498 21138 4510
rect 21534 4562 21586 4574
rect 21534 4498 21586 4510
rect 21982 4562 22034 4574
rect 21982 4498 22034 4510
rect 22766 4562 22818 4574
rect 22766 4498 22818 4510
rect 23214 4562 23266 4574
rect 23214 4498 23266 4510
rect 23662 4562 23714 4574
rect 23662 4498 23714 4510
rect 24110 4562 24162 4574
rect 24110 4498 24162 4510
rect 24670 4562 24722 4574
rect 24670 4498 24722 4510
rect 25454 4562 25506 4574
rect 25454 4498 25506 4510
rect 25902 4562 25954 4574
rect 25902 4498 25954 4510
rect 26686 4562 26738 4574
rect 26686 4498 26738 4510
rect 27022 4562 27074 4574
rect 27022 4498 27074 4510
rect 28478 4562 28530 4574
rect 28478 4498 28530 4510
rect 28926 4562 28978 4574
rect 28926 4498 28978 4510
rect 29262 4562 29314 4574
rect 29262 4498 29314 4510
rect 31390 4562 31442 4574
rect 31390 4498 31442 4510
rect 33966 4562 34018 4574
rect 33966 4498 34018 4510
rect 36878 4562 36930 4574
rect 36878 4498 36930 4510
rect 41022 4562 41074 4574
rect 47630 4562 47682 4574
rect 42130 4510 42142 4562
rect 42194 4510 42206 4562
rect 41022 4498 41074 4510
rect 47630 4498 47682 4510
rect 48974 4562 49026 4574
rect 48974 4498 49026 4510
rect 47294 4450 47346 4462
rect 30146 4398 30158 4450
rect 30210 4398 30222 4450
rect 33058 4398 33070 4450
rect 33122 4398 33134 4450
rect 35970 4398 35982 4450
rect 36034 4398 36046 4450
rect 45714 4398 45726 4450
rect 45778 4398 45790 4450
rect 47294 4386 47346 4398
rect 48078 4450 48130 4462
rect 48078 4386 48130 4398
rect 27918 4338 27970 4350
rect 27918 4274 27970 4286
rect 31950 4338 32002 4350
rect 33406 4338 33458 4350
rect 46734 4338 46786 4350
rect 32386 4286 32398 4338
rect 32450 4286 32462 4338
rect 40226 4286 40238 4338
rect 40290 4286 40302 4338
rect 43810 4286 43822 4338
rect 43874 4286 43886 4338
rect 31950 4274 32002 4286
rect 33406 4274 33458 4286
rect 46734 4274 46786 4286
rect 27582 4226 27634 4238
rect 49310 4226 49362 4238
rect 37314 4174 37326 4226
rect 37378 4174 37390 4226
rect 38210 4174 38222 4226
rect 38274 4174 38286 4226
rect 27582 4162 27634 4174
rect 49310 4162 49362 4174
rect 27570 4062 27582 4114
rect 27634 4111 27646 4114
rect 28466 4111 28478 4114
rect 27634 4065 28478 4111
rect 27634 4062 27646 4065
rect 28466 4062 28478 4065
rect 28530 4062 28542 4114
rect 1344 3946 62608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 62608 3946
rect 1344 3860 62608 3894
rect 36094 3778 36146 3790
rect 36094 3714 36146 3726
rect 38334 3778 38386 3790
rect 45938 3726 45950 3778
rect 46002 3775 46014 3778
rect 46946 3775 46958 3778
rect 46002 3729 46958 3775
rect 46002 3726 46014 3729
rect 46946 3726 46958 3729
rect 47010 3726 47022 3778
rect 38334 3714 38386 3726
rect 23550 3666 23602 3678
rect 23550 3602 23602 3614
rect 24110 3666 24162 3678
rect 24110 3602 24162 3614
rect 24782 3666 24834 3678
rect 24782 3602 24834 3614
rect 25230 3666 25282 3678
rect 25230 3602 25282 3614
rect 26126 3666 26178 3678
rect 26126 3602 26178 3614
rect 27470 3666 27522 3678
rect 27470 3602 27522 3614
rect 27918 3666 27970 3678
rect 27918 3602 27970 3614
rect 28926 3666 28978 3678
rect 28926 3602 28978 3614
rect 29598 3666 29650 3678
rect 29598 3602 29650 3614
rect 31054 3666 31106 3678
rect 31054 3602 31106 3614
rect 33518 3666 33570 3678
rect 33518 3602 33570 3614
rect 39006 3666 39058 3678
rect 43822 3666 43874 3678
rect 40562 3614 40574 3666
rect 40626 3614 40638 3666
rect 42690 3614 42702 3666
rect 42754 3614 42766 3666
rect 39006 3602 39058 3614
rect 43822 3602 43874 3614
rect 45166 3666 45218 3678
rect 45166 3602 45218 3614
rect 45502 3666 45554 3678
rect 45502 3602 45554 3614
rect 46062 3666 46114 3678
rect 46062 3602 46114 3614
rect 46510 3666 46562 3678
rect 46510 3602 46562 3614
rect 46958 3666 47010 3678
rect 46958 3602 47010 3614
rect 47966 3666 48018 3678
rect 47966 3602 48018 3614
rect 48526 3666 48578 3678
rect 48526 3602 48578 3614
rect 25678 3554 25730 3566
rect 33406 3554 33458 3566
rect 30034 3502 30046 3554
rect 30098 3502 30110 3554
rect 31378 3502 31390 3554
rect 31442 3502 31454 3554
rect 33058 3502 33070 3554
rect 33122 3502 33134 3554
rect 25678 3490 25730 3502
rect 33406 3490 33458 3502
rect 33630 3554 33682 3566
rect 33630 3490 33682 3502
rect 33966 3554 34018 3566
rect 33966 3490 34018 3502
rect 34974 3554 35026 3566
rect 34974 3490 35026 3502
rect 38446 3554 38498 3566
rect 44270 3554 44322 3566
rect 39890 3502 39902 3554
rect 39954 3502 39966 3554
rect 38446 3490 38498 3502
rect 44270 3490 44322 3502
rect 47518 3554 47570 3566
rect 47518 3490 47570 3502
rect 26574 3442 26626 3454
rect 26574 3378 26626 3390
rect 27022 3442 27074 3454
rect 27022 3378 27074 3390
rect 29822 3442 29874 3454
rect 29822 3378 29874 3390
rect 31614 3442 31666 3454
rect 31614 3378 31666 3390
rect 32398 3442 32450 3454
rect 34638 3442 34690 3454
rect 32722 3390 32734 3442
rect 32786 3390 32798 3442
rect 34290 3390 34302 3442
rect 34354 3390 34366 3442
rect 32398 3378 32450 3390
rect 34638 3378 34690 3390
rect 35534 3442 35586 3454
rect 38334 3442 38386 3454
rect 37202 3390 37214 3442
rect 37266 3390 37278 3442
rect 35534 3378 35586 3390
rect 38334 3378 38386 3390
rect 44606 3442 44658 3454
rect 44606 3378 44658 3390
rect 7646 3330 7698 3342
rect 7646 3266 7698 3278
rect 1344 3162 62608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 62608 3162
rect 1344 3076 62608 3110
<< via1 >>
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 17950 60174 18002 60226
rect 48974 60174 49026 60226
rect 27582 60062 27634 60114
rect 15374 59950 15426 60002
rect 16942 59950 16994 60002
rect 28590 59950 28642 60002
rect 33966 59950 34018 60002
rect 34974 59950 35026 60002
rect 47966 59950 48018 60002
rect 13582 59838 13634 59890
rect 13806 59838 13858 59890
rect 19966 59838 20018 59890
rect 20862 59838 20914 59890
rect 23214 59838 23266 59890
rect 23774 59838 23826 59890
rect 23886 59838 23938 59890
rect 27358 59838 27410 59890
rect 31166 59838 31218 59890
rect 33070 59838 33122 59890
rect 38558 59838 38610 59890
rect 14142 59726 14194 59778
rect 14478 59726 14530 59778
rect 14814 59726 14866 59778
rect 15374 59726 15426 59778
rect 15934 59726 15986 59778
rect 16158 59726 16210 59778
rect 16270 59726 16322 59778
rect 16382 59726 16434 59778
rect 20078 59726 20130 59778
rect 20302 59726 20354 59778
rect 20974 59726 21026 59778
rect 21198 59726 21250 59778
rect 22094 59726 22146 59778
rect 24110 59726 24162 59778
rect 25006 59726 25058 59778
rect 26350 59726 26402 59778
rect 28366 59726 28418 59778
rect 29822 59726 29874 59778
rect 32174 59726 32226 59778
rect 32286 59726 32338 59778
rect 32398 59726 32450 59778
rect 32622 59726 32674 59778
rect 33182 59726 33234 59778
rect 33742 59726 33794 59778
rect 34638 59726 34690 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 14030 59390 14082 59442
rect 16158 59390 16210 59442
rect 22094 59390 22146 59442
rect 27470 59390 27522 59442
rect 30046 59390 30098 59442
rect 49758 59390 49810 59442
rect 14926 59278 14978 59330
rect 17950 59278 18002 59330
rect 24334 59278 24386 59330
rect 30830 59278 30882 59330
rect 33742 59278 33794 59330
rect 34190 59278 34242 59330
rect 34750 59278 34802 59330
rect 62190 59278 62242 59330
rect 20526 59166 20578 59218
rect 24558 59166 24610 59218
rect 25566 59166 25618 59218
rect 26462 59166 26514 59218
rect 35086 59166 35138 59218
rect 48750 59166 48802 59218
rect 16942 59054 16994 59106
rect 23774 59054 23826 59106
rect 29598 59054 29650 59106
rect 35534 59054 35586 59106
rect 36094 59054 36146 59106
rect 19406 58942 19458 58994
rect 23438 58942 23490 58994
rect 26126 58942 26178 58994
rect 32622 58942 32674 58994
rect 33182 58942 33234 58994
rect 33518 58942 33570 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 13470 58606 13522 58658
rect 13806 58606 13858 58658
rect 24894 58606 24946 58658
rect 29486 58606 29538 58658
rect 33742 58606 33794 58658
rect 20414 58494 20466 58546
rect 21982 58494 22034 58546
rect 52110 58494 52162 58546
rect 52782 58494 52834 58546
rect 17950 58382 18002 58434
rect 18510 58382 18562 58434
rect 19182 58382 19234 58434
rect 19630 58382 19682 58434
rect 22542 58382 22594 58434
rect 22878 58382 22930 58434
rect 24110 58382 24162 58434
rect 24782 58382 24834 58434
rect 25006 58382 25058 58434
rect 27022 58382 27074 58434
rect 27806 58382 27858 58434
rect 29598 58382 29650 58434
rect 31166 58382 31218 58434
rect 31278 58382 31330 58434
rect 51326 58382 51378 58434
rect 14030 58270 14082 58322
rect 14702 58270 14754 58322
rect 27694 58270 27746 58322
rect 30158 58270 30210 58322
rect 50766 58270 50818 58322
rect 16494 58158 16546 58210
rect 17166 58158 17218 58210
rect 17838 58158 17890 58210
rect 21310 58158 21362 58210
rect 21646 58158 21698 58210
rect 26686 58158 26738 58210
rect 28254 58158 28306 58210
rect 28590 58158 28642 58210
rect 35198 58158 35250 58210
rect 36430 58158 36482 58210
rect 37102 58158 37154 58210
rect 40798 58158 40850 58210
rect 41134 58158 41186 58210
rect 44382 58158 44434 58210
rect 45166 58158 45218 58210
rect 45614 58158 45666 58210
rect 46062 58158 46114 58210
rect 47630 58158 47682 58210
rect 48078 58158 48130 58210
rect 48526 58158 48578 58210
rect 48974 58158 49026 58210
rect 49422 58158 49474 58210
rect 49870 58158 49922 58210
rect 50206 58158 50258 58210
rect 51662 58158 51714 58210
rect 53230 58158 53282 58210
rect 54462 58158 54514 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 14030 57822 14082 57874
rect 14478 57822 14530 57874
rect 14590 57822 14642 57874
rect 24558 57822 24610 57874
rect 24670 57822 24722 57874
rect 40014 57822 40066 57874
rect 42254 57822 42306 57874
rect 43710 57822 43762 57874
rect 47518 57822 47570 57874
rect 48190 57822 48242 57874
rect 49198 57822 49250 57874
rect 14702 57710 14754 57762
rect 15710 57710 15762 57762
rect 16158 57710 16210 57762
rect 19406 57710 19458 57762
rect 24334 57710 24386 57762
rect 24446 57710 24498 57762
rect 33630 57710 33682 57762
rect 35198 57710 35250 57762
rect 36430 57710 36482 57762
rect 44718 57710 44770 57762
rect 49758 57710 49810 57762
rect 51886 57710 51938 57762
rect 52110 57710 52162 57762
rect 56814 57710 56866 57762
rect 14366 57598 14418 57650
rect 15038 57598 15090 57650
rect 16382 57598 16434 57650
rect 18846 57598 18898 57650
rect 19182 57598 19234 57650
rect 19630 57598 19682 57650
rect 19966 57598 20018 57650
rect 21198 57598 21250 57650
rect 21870 57598 21922 57650
rect 22094 57598 22146 57650
rect 23886 57598 23938 57650
rect 25678 57598 25730 57650
rect 26014 57598 26066 57650
rect 28142 57598 28194 57650
rect 29262 57598 29314 57650
rect 29598 57598 29650 57650
rect 30158 57598 30210 57650
rect 31166 57598 31218 57650
rect 32398 57598 32450 57650
rect 33742 57598 33794 57650
rect 34302 57598 34354 57650
rect 35534 57598 35586 57650
rect 47966 57598 48018 57650
rect 49982 57598 50034 57650
rect 51438 57598 51490 57650
rect 52334 57598 52386 57650
rect 52558 57598 52610 57650
rect 52894 57598 52946 57650
rect 53118 57598 53170 57650
rect 53566 57598 53618 57650
rect 53790 57598 53842 57650
rect 54014 57598 54066 57650
rect 55806 57598 55858 57650
rect 12686 57486 12738 57538
rect 13134 57486 13186 57538
rect 13582 57486 13634 57538
rect 18174 57486 18226 57538
rect 19294 57486 19346 57538
rect 26126 57486 26178 57538
rect 28478 57486 28530 57538
rect 29822 57486 29874 57538
rect 31726 57486 31778 57538
rect 36094 57486 36146 57538
rect 36878 57486 36930 57538
rect 37326 57486 37378 57538
rect 37774 57486 37826 57538
rect 41246 57486 41298 57538
rect 41806 57486 41858 57538
rect 46510 57486 46562 57538
rect 47070 57486 47122 57538
rect 50654 57486 50706 57538
rect 50990 57486 51042 57538
rect 52782 57486 52834 57538
rect 53678 57486 53730 57538
rect 55022 57486 55074 57538
rect 55470 57486 55522 57538
rect 16718 57374 16770 57426
rect 17614 57374 17666 57426
rect 17950 57374 18002 57426
rect 23214 57374 23266 57426
rect 34638 57374 34690 57426
rect 45838 57374 45890 57426
rect 46174 57374 46226 57426
rect 46734 57374 46786 57426
rect 51774 57374 51826 57426
rect 54462 57374 54514 57426
rect 54798 57374 54850 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 15262 57038 15314 57090
rect 15598 57038 15650 57090
rect 17166 57038 17218 57090
rect 25678 57038 25730 57090
rect 32174 57038 32226 57090
rect 32510 57038 32562 57090
rect 37214 57038 37266 57090
rect 38558 57038 38610 57090
rect 51438 57038 51490 57090
rect 55022 57038 55074 57090
rect 12126 56926 12178 56978
rect 14030 56926 14082 56978
rect 15038 56926 15090 56978
rect 19406 56926 19458 56978
rect 21310 56926 21362 56978
rect 26462 56926 26514 56978
rect 31166 56926 31218 56978
rect 32734 56926 32786 56978
rect 33406 56926 33458 56978
rect 38558 56926 38610 56978
rect 39566 56926 39618 56978
rect 41358 56926 41410 56978
rect 42702 56926 42754 56978
rect 44942 56926 44994 56978
rect 56366 56926 56418 56978
rect 57822 56926 57874 56978
rect 13022 56814 13074 56866
rect 13582 56814 13634 56866
rect 16046 56814 16098 56866
rect 16830 56814 16882 56866
rect 18510 56814 18562 56866
rect 19518 56814 19570 56866
rect 20526 56814 20578 56866
rect 20750 56814 20802 56866
rect 22094 56814 22146 56866
rect 22766 56814 22818 56866
rect 24110 56814 24162 56866
rect 26686 56814 26738 56866
rect 27582 56814 27634 56866
rect 29598 56814 29650 56866
rect 30382 56814 30434 56866
rect 30606 56814 30658 56866
rect 40686 56814 40738 56866
rect 40910 56814 40962 56866
rect 41470 56814 41522 56866
rect 42590 56814 42642 56866
rect 55694 56814 55746 56866
rect 57262 56814 57314 56866
rect 14366 56702 14418 56754
rect 14702 56702 14754 56754
rect 16270 56702 16322 56754
rect 17614 56702 17666 56754
rect 18174 56702 18226 56754
rect 18734 56702 18786 56754
rect 19742 56702 19794 56754
rect 21422 56702 21474 56754
rect 21982 56702 22034 56754
rect 23998 56702 24050 56754
rect 24558 56702 24610 56754
rect 28030 56702 28082 56754
rect 29262 56702 29314 56754
rect 29934 56702 29986 56754
rect 31278 56702 31330 56754
rect 31390 56702 31442 56754
rect 31502 56702 31554 56754
rect 33070 56702 33122 56754
rect 33742 56702 33794 56754
rect 35086 56702 35138 56754
rect 37102 56702 37154 56754
rect 40462 56702 40514 56754
rect 42254 56702 42306 56754
rect 45838 56702 45890 56754
rect 46510 56702 46562 56754
rect 47630 56702 47682 56754
rect 53790 56702 53842 56754
rect 55470 56702 55522 56754
rect 57038 56702 57090 56754
rect 58270 56702 58322 56754
rect 11678 56590 11730 56642
rect 12574 56590 12626 56642
rect 17726 56590 17778 56642
rect 17950 56590 18002 56642
rect 18286 56590 18338 56642
rect 23102 56590 23154 56642
rect 24334 56590 24386 56642
rect 24446 56590 24498 56642
rect 31054 56590 31106 56642
rect 33294 56590 33346 56642
rect 33854 56590 33906 56642
rect 33966 56590 34018 56642
rect 36206 56590 36258 56642
rect 37662 56590 37714 56642
rect 37998 56590 38050 56642
rect 38894 56590 38946 56642
rect 40126 56590 40178 56642
rect 40798 56590 40850 56642
rect 43486 56590 43538 56642
rect 44046 56590 44098 56642
rect 45502 56590 45554 56642
rect 46174 56590 46226 56642
rect 48974 56590 49026 56642
rect 50094 56590 50146 56642
rect 52222 56590 52274 56642
rect 52894 56590 52946 56642
rect 56030 56590 56082 56642
rect 56478 56590 56530 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 15598 56254 15650 56306
rect 21198 56254 21250 56306
rect 23662 56254 23714 56306
rect 30382 56254 30434 56306
rect 31390 56254 31442 56306
rect 32062 56254 32114 56306
rect 32398 56254 32450 56306
rect 38446 56254 38498 56306
rect 38558 56254 38610 56306
rect 46734 56254 46786 56306
rect 48078 56254 48130 56306
rect 48862 56254 48914 56306
rect 51662 56254 51714 56306
rect 55358 56254 55410 56306
rect 58382 56254 58434 56306
rect 59278 56254 59330 56306
rect 16158 56142 16210 56194
rect 16606 56142 16658 56194
rect 21870 56142 21922 56194
rect 22990 56142 23042 56194
rect 23550 56142 23602 56194
rect 24334 56142 24386 56194
rect 25566 56142 25618 56194
rect 27022 56142 27074 56194
rect 27470 56142 27522 56194
rect 28142 56142 28194 56194
rect 28814 56142 28866 56194
rect 29150 56142 29202 56194
rect 30494 56142 30546 56194
rect 31614 56142 31666 56194
rect 32174 56142 32226 56194
rect 34638 56142 34690 56194
rect 42926 56142 42978 56194
rect 45278 56142 45330 56194
rect 45614 56142 45666 56194
rect 47070 56142 47122 56194
rect 49870 56142 49922 56194
rect 55582 56142 55634 56194
rect 57822 56142 57874 56194
rect 15038 56030 15090 56082
rect 15934 56030 15986 56082
rect 17502 56030 17554 56082
rect 18510 56030 18562 56082
rect 19742 56030 19794 56082
rect 20190 56030 20242 56082
rect 20638 56030 20690 56082
rect 21086 56030 21138 56082
rect 22094 56030 22146 56082
rect 22430 56030 22482 56082
rect 22766 56030 22818 56082
rect 23438 56030 23490 56082
rect 25230 56030 25282 56082
rect 25790 56030 25842 56082
rect 25902 56030 25954 56082
rect 27582 56030 27634 56082
rect 27918 56030 27970 56082
rect 29374 56030 29426 56082
rect 29598 56030 29650 56082
rect 29934 56030 29986 56082
rect 30830 56030 30882 56082
rect 31278 56030 31330 56082
rect 31950 56030 32002 56082
rect 33182 56030 33234 56082
rect 33630 56030 33682 56082
rect 33854 56030 33906 56082
rect 35422 56030 35474 56082
rect 36206 56030 36258 56082
rect 37102 56030 37154 56082
rect 37886 56030 37938 56082
rect 38334 56030 38386 56082
rect 45950 56030 46002 56082
rect 48190 56030 48242 56082
rect 49758 56030 49810 56082
rect 50542 56030 50594 56082
rect 54910 56030 54962 56082
rect 55134 56030 55186 56082
rect 57038 56030 57090 56082
rect 57710 56030 57762 56082
rect 58270 56030 58322 56082
rect 11230 55918 11282 55970
rect 11678 55918 11730 55970
rect 12126 55918 12178 55970
rect 12574 55918 12626 55970
rect 13022 55918 13074 55970
rect 13470 55918 13522 55970
rect 13806 55918 13858 55970
rect 14366 55918 14418 55970
rect 14702 55918 14754 55970
rect 18174 55918 18226 55970
rect 33406 55918 33458 55970
rect 34638 55918 34690 55970
rect 37662 55918 37714 55970
rect 39006 55918 39058 55970
rect 39454 55918 39506 55970
rect 40126 55918 40178 55970
rect 41022 55918 41074 55970
rect 41470 55918 41522 55970
rect 42254 55918 42306 55970
rect 47630 55918 47682 55970
rect 54238 55918 54290 55970
rect 55358 55918 55410 55970
rect 56142 55918 56194 55970
rect 13022 55806 13074 55858
rect 14366 55806 14418 55858
rect 23102 55806 23154 55858
rect 27470 55806 27522 55858
rect 30382 55806 30434 55858
rect 31166 55806 31218 55858
rect 33070 55806 33122 55858
rect 44830 55806 44882 55858
rect 46286 55806 46338 55858
rect 49198 55806 49250 55858
rect 50430 55806 50482 55858
rect 53118 55806 53170 55858
rect 56702 55806 56754 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 20638 55470 20690 55522
rect 31054 55470 31106 55522
rect 35310 55470 35362 55522
rect 41022 55470 41074 55522
rect 55806 55470 55858 55522
rect 15486 55358 15538 55410
rect 18398 55358 18450 55410
rect 23774 55358 23826 55410
rect 25342 55358 25394 55410
rect 29598 55358 29650 55410
rect 30158 55358 30210 55410
rect 32734 55358 32786 55410
rect 38894 55358 38946 55410
rect 42926 55358 42978 55410
rect 46174 55358 46226 55410
rect 47742 55358 47794 55410
rect 23438 55246 23490 55298
rect 24222 55246 24274 55298
rect 24782 55246 24834 55298
rect 25230 55246 25282 55298
rect 25678 55246 25730 55298
rect 26574 55246 26626 55298
rect 27134 55246 27186 55298
rect 27694 55246 27746 55298
rect 28478 55246 28530 55298
rect 29262 55246 29314 55298
rect 29486 55246 29538 55298
rect 29822 55246 29874 55298
rect 30046 55246 30098 55298
rect 30718 55246 30770 55298
rect 31390 55246 31442 55298
rect 32174 55246 32226 55298
rect 32622 55246 32674 55298
rect 35646 55246 35698 55298
rect 36990 55246 37042 55298
rect 39006 55246 39058 55298
rect 39678 55246 39730 55298
rect 40574 55246 40626 55298
rect 42590 55246 42642 55298
rect 43374 55246 43426 55298
rect 45726 55246 45778 55298
rect 47966 55246 48018 55298
rect 48750 55246 48802 55298
rect 49310 55246 49362 55298
rect 50318 55246 50370 55298
rect 52670 55246 52722 55298
rect 53230 55246 53282 55298
rect 53902 55246 53954 55298
rect 55582 55246 55634 55298
rect 56702 55246 56754 55298
rect 58158 55246 58210 55298
rect 1710 55134 1762 55186
rect 14142 55134 14194 55186
rect 16494 55134 16546 55186
rect 19182 55134 19234 55186
rect 25566 55134 25618 55186
rect 26686 55134 26738 55186
rect 27806 55134 27858 55186
rect 30270 55134 30322 55186
rect 31950 55134 32002 55186
rect 33406 55134 33458 55186
rect 37326 55134 37378 55186
rect 42814 55134 42866 55186
rect 42926 55134 42978 55186
rect 45502 55134 45554 55186
rect 46510 55134 46562 55186
rect 48414 55134 48466 55186
rect 54126 55134 54178 55186
rect 55470 55134 55522 55186
rect 58718 55134 58770 55186
rect 58942 55134 58994 55186
rect 59278 55134 59330 55186
rect 59614 55134 59666 55186
rect 61070 55134 61122 55186
rect 2046 55022 2098 55074
rect 2494 55022 2546 55074
rect 9998 55022 10050 55074
rect 10558 55022 10610 55074
rect 11006 55022 11058 55074
rect 11454 55022 11506 55074
rect 11902 55022 11954 55074
rect 12350 55022 12402 55074
rect 13022 55022 13074 55074
rect 21982 55022 22034 55074
rect 23102 55022 23154 55074
rect 26910 55022 26962 55074
rect 28254 55022 28306 55074
rect 35870 55022 35922 55074
rect 36318 55022 36370 55074
rect 41918 55022 41970 55074
rect 42254 55022 42306 55074
rect 43934 55022 43986 55074
rect 44270 55022 44322 55074
rect 44942 55022 44994 55074
rect 47182 55022 47234 55074
rect 47406 55022 47458 55074
rect 51214 55022 51266 55074
rect 51662 55022 51714 55074
rect 51886 55022 51938 55074
rect 51998 55022 52050 55074
rect 52110 55022 52162 55074
rect 53566 55022 53618 55074
rect 58382 55022 58434 55074
rect 58494 55022 58546 55074
rect 60734 55022 60786 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 12686 54686 12738 54738
rect 13246 54686 13298 54738
rect 14590 54686 14642 54738
rect 15038 54686 15090 54738
rect 20862 54686 20914 54738
rect 29486 54686 29538 54738
rect 36318 54686 36370 54738
rect 37774 54686 37826 54738
rect 39342 54686 39394 54738
rect 44718 54686 44770 54738
rect 47070 54686 47122 54738
rect 48750 54686 48802 54738
rect 59390 54686 59442 54738
rect 13806 54574 13858 54626
rect 15934 54574 15986 54626
rect 16718 54574 16770 54626
rect 17390 54574 17442 54626
rect 17614 54574 17666 54626
rect 18510 54574 18562 54626
rect 20302 54574 20354 54626
rect 20974 54574 21026 54626
rect 21534 54574 21586 54626
rect 21870 54574 21922 54626
rect 22542 54574 22594 54626
rect 23886 54574 23938 54626
rect 24558 54574 24610 54626
rect 28478 54574 28530 54626
rect 30942 54574 30994 54626
rect 31390 54574 31442 54626
rect 32174 54574 32226 54626
rect 32510 54574 32562 54626
rect 37214 54574 37266 54626
rect 38446 54574 38498 54626
rect 45614 54574 45666 54626
rect 47406 54574 47458 54626
rect 47630 54574 47682 54626
rect 49870 54574 49922 54626
rect 52110 54574 52162 54626
rect 52782 54574 52834 54626
rect 53230 54574 53282 54626
rect 55918 54574 55970 54626
rect 12462 54462 12514 54514
rect 12798 54462 12850 54514
rect 13134 54462 13186 54514
rect 13694 54462 13746 54514
rect 14254 54462 14306 54514
rect 15374 54462 15426 54514
rect 16158 54462 16210 54514
rect 16830 54462 16882 54514
rect 17950 54462 18002 54514
rect 18622 54462 18674 54514
rect 18958 54462 19010 54514
rect 19518 54462 19570 54514
rect 20190 54462 20242 54514
rect 21646 54462 21698 54514
rect 22094 54462 22146 54514
rect 23438 54462 23490 54514
rect 24334 54462 24386 54514
rect 28030 54462 28082 54514
rect 28702 54462 28754 54514
rect 29262 54462 29314 54514
rect 29486 54462 29538 54514
rect 29710 54462 29762 54514
rect 30158 54462 30210 54514
rect 30606 54462 30658 54514
rect 31278 54462 31330 54514
rect 33182 54462 33234 54514
rect 36654 54462 36706 54514
rect 36878 54462 36930 54514
rect 37438 54462 37490 54514
rect 38110 54462 38162 54514
rect 41358 54462 41410 54514
rect 45054 54462 45106 54514
rect 45726 54462 45778 54514
rect 46286 54462 46338 54514
rect 46622 54462 46674 54514
rect 46958 54462 47010 54514
rect 50430 54462 50482 54514
rect 51662 54462 51714 54514
rect 53454 54462 53506 54514
rect 53790 54462 53842 54514
rect 54462 54462 54514 54514
rect 54686 54462 54738 54514
rect 56590 54462 56642 54514
rect 9662 54350 9714 54402
rect 10222 54350 10274 54402
rect 10670 54350 10722 54402
rect 11006 54350 11058 54402
rect 11790 54350 11842 54402
rect 12126 54350 12178 54402
rect 17502 54350 17554 54402
rect 17838 54350 17890 54402
rect 19854 54350 19906 54402
rect 21310 54350 21362 54402
rect 25230 54350 25282 54402
rect 27358 54350 27410 54402
rect 33854 54350 33906 54402
rect 35982 54350 36034 54402
rect 38894 54350 38946 54402
rect 39790 54350 39842 54402
rect 40238 54350 40290 54402
rect 41134 54350 41186 54402
rect 42142 54350 42194 54402
rect 44270 54350 44322 54402
rect 47518 54350 47570 54402
rect 48190 54350 48242 54402
rect 49310 54350 49362 54402
rect 55694 54350 55746 54402
rect 60510 54350 60562 54402
rect 61070 54350 61122 54402
rect 61518 54350 61570 54402
rect 61854 54350 61906 54402
rect 12238 54238 12290 54290
rect 13246 54238 13298 54290
rect 13806 54238 13858 54290
rect 16718 54238 16770 54290
rect 22990 54238 23042 54290
rect 24670 54238 24722 54290
rect 38782 54238 38834 54290
rect 39342 54238 39394 54290
rect 46846 54238 46898 54290
rect 48078 54238 48130 54290
rect 49086 54238 49138 54290
rect 54350 54238 54402 54290
rect 56702 54238 56754 54290
rect 57934 54238 57986 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 10670 53902 10722 53954
rect 13806 53902 13858 53954
rect 16270 53902 16322 53954
rect 23998 53902 24050 53954
rect 27694 53902 27746 53954
rect 30158 53902 30210 53954
rect 30382 53902 30434 53954
rect 30830 53902 30882 53954
rect 31278 53902 31330 53954
rect 44942 53902 44994 53954
rect 52894 53902 52946 53954
rect 56926 53902 56978 53954
rect 57710 53902 57762 53954
rect 11678 53790 11730 53842
rect 18846 53790 18898 53842
rect 20750 53790 20802 53842
rect 21982 53790 22034 53842
rect 22206 53790 22258 53842
rect 25118 53790 25170 53842
rect 31502 53790 31554 53842
rect 31838 53790 31890 53842
rect 45390 53790 45442 53842
rect 51102 53790 51154 53842
rect 58158 53790 58210 53842
rect 61294 53790 61346 53842
rect 10110 53678 10162 53730
rect 10894 53678 10946 53730
rect 12910 53678 12962 53730
rect 13694 53678 13746 53730
rect 14142 53678 14194 53730
rect 14814 53678 14866 53730
rect 15150 53678 15202 53730
rect 15486 53678 15538 53730
rect 15710 53678 15762 53730
rect 16046 53678 16098 53730
rect 16270 53678 16322 53730
rect 17278 53678 17330 53730
rect 18174 53678 18226 53730
rect 18734 53678 18786 53730
rect 19070 53678 19122 53730
rect 19854 53678 19906 53730
rect 21534 53678 21586 53730
rect 22318 53678 22370 53730
rect 24782 53678 24834 53730
rect 25454 53678 25506 53730
rect 26686 53678 26738 53730
rect 27246 53678 27298 53730
rect 27470 53678 27522 53730
rect 27918 53678 27970 53730
rect 29262 53678 29314 53730
rect 30718 53678 30770 53730
rect 31950 53678 32002 53730
rect 36094 53678 36146 53730
rect 36206 53678 36258 53730
rect 39454 53678 39506 53730
rect 40014 53678 40066 53730
rect 43262 53678 43314 53730
rect 43710 53678 43762 53730
rect 44270 53678 44322 53730
rect 45614 53678 45666 53730
rect 48862 53678 48914 53730
rect 49086 53678 49138 53730
rect 49534 53678 49586 53730
rect 49758 53678 49810 53730
rect 50990 53678 51042 53730
rect 51998 53678 52050 53730
rect 53678 53678 53730 53730
rect 55134 53678 55186 53730
rect 55582 53678 55634 53730
rect 55918 53678 55970 53730
rect 58046 53678 58098 53730
rect 58382 53678 58434 53730
rect 59054 53678 59106 53730
rect 9662 53566 9714 53618
rect 11454 53566 11506 53618
rect 12350 53566 12402 53618
rect 12574 53566 12626 53618
rect 16830 53566 16882 53618
rect 17166 53566 17218 53618
rect 17838 53566 17890 53618
rect 28478 53566 28530 53618
rect 28590 53566 28642 53618
rect 30942 53566 30994 53618
rect 32398 53566 32450 53618
rect 34302 53566 34354 53618
rect 37662 53566 37714 53618
rect 40910 53566 40962 53618
rect 41246 53566 41298 53618
rect 41582 53566 41634 53618
rect 44046 53566 44098 53618
rect 44830 53566 44882 53618
rect 45054 53566 45106 53618
rect 46510 53566 46562 53618
rect 50094 53566 50146 53618
rect 51214 53566 51266 53618
rect 51662 53566 51714 53618
rect 52670 53566 52722 53618
rect 8654 53454 8706 53506
rect 9102 53454 9154 53506
rect 10558 53454 10610 53506
rect 11790 53454 11842 53506
rect 13582 53454 13634 53506
rect 14478 53454 14530 53506
rect 15262 53454 15314 53506
rect 15822 53454 15874 53506
rect 16942 53454 16994 53506
rect 18510 53454 18562 53506
rect 19294 53454 19346 53506
rect 20190 53454 20242 53506
rect 27582 53454 27634 53506
rect 28254 53454 28306 53506
rect 29710 53454 29762 53506
rect 31726 53454 31778 53506
rect 32510 53454 32562 53506
rect 32846 53454 32898 53506
rect 33182 53454 33234 53506
rect 35422 53454 35474 53506
rect 38782 53454 38834 53506
rect 39230 53454 39282 53506
rect 40686 53454 40738 53506
rect 41918 53454 41970 53506
rect 42366 53454 42418 53506
rect 43038 53454 43090 53506
rect 43934 53454 43986 53506
rect 48302 53454 48354 53506
rect 48974 53454 49026 53506
rect 53230 53454 53282 53506
rect 59614 53454 59666 53506
rect 60734 53454 60786 53506
rect 61854 53454 61906 53506
rect 62190 53454 62242 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 9102 53118 9154 53170
rect 9886 53118 9938 53170
rect 19966 53118 20018 53170
rect 25342 53118 25394 53170
rect 25790 53118 25842 53170
rect 25902 53118 25954 53170
rect 27022 53118 27074 53170
rect 28142 53118 28194 53170
rect 29262 53118 29314 53170
rect 29710 53118 29762 53170
rect 45502 53118 45554 53170
rect 46398 53118 46450 53170
rect 53566 53118 53618 53170
rect 53790 53118 53842 53170
rect 60734 53118 60786 53170
rect 15038 53006 15090 53058
rect 16606 53006 16658 53058
rect 17838 53006 17890 53058
rect 18734 53006 18786 53058
rect 22206 53006 22258 53058
rect 25230 53006 25282 53058
rect 26686 53006 26738 53058
rect 32398 53006 32450 53058
rect 39006 53006 39058 53058
rect 39342 53006 39394 53058
rect 40910 53006 40962 53058
rect 42702 53006 42754 53058
rect 45278 53006 45330 53058
rect 46510 53006 46562 53058
rect 46734 53006 46786 53058
rect 47966 53006 48018 53058
rect 49982 53006 50034 53058
rect 53902 53006 53954 53058
rect 55022 53006 55074 53058
rect 57486 53006 57538 53058
rect 58830 53006 58882 53058
rect 7758 52894 7810 52946
rect 14366 52894 14418 52946
rect 15150 52894 15202 52946
rect 15598 52894 15650 52946
rect 15822 52894 15874 52946
rect 16382 52894 16434 52946
rect 20414 52894 20466 52946
rect 20638 52894 20690 52946
rect 21086 52894 21138 52946
rect 21534 52894 21586 52946
rect 23214 52894 23266 52946
rect 25566 52894 25618 52946
rect 26014 52894 26066 52946
rect 26462 52894 26514 52946
rect 30494 52894 30546 52946
rect 31278 52894 31330 52946
rect 32174 52894 32226 52946
rect 32510 52894 32562 52946
rect 33294 52894 33346 52946
rect 33518 52894 33570 52946
rect 33966 52894 34018 52946
rect 34526 52894 34578 52946
rect 35086 52894 35138 52946
rect 40126 52894 40178 52946
rect 41134 52894 41186 52946
rect 45054 52894 45106 52946
rect 45838 52894 45890 52946
rect 46062 52894 46114 52946
rect 47518 52894 47570 52946
rect 47742 52894 47794 52946
rect 48190 52894 48242 52946
rect 49198 52894 49250 52946
rect 49422 52894 49474 52946
rect 49870 52894 49922 52946
rect 50990 52894 51042 52946
rect 51326 52894 51378 52946
rect 51550 52894 51602 52946
rect 51998 52894 52050 52946
rect 52558 52894 52610 52946
rect 54238 52894 54290 52946
rect 54798 52894 54850 52946
rect 56814 52894 56866 52946
rect 57822 52894 57874 52946
rect 59054 52894 59106 52946
rect 59614 52894 59666 52946
rect 8094 52782 8146 52834
rect 8542 52782 8594 52834
rect 10446 52782 10498 52834
rect 10894 52782 10946 52834
rect 11230 52782 11282 52834
rect 11566 52782 11618 52834
rect 13694 52782 13746 52834
rect 17502 52782 17554 52834
rect 20526 52782 20578 52834
rect 23326 52782 23378 52834
rect 30158 52782 30210 52834
rect 31502 52782 31554 52834
rect 33406 52782 33458 52834
rect 34750 52782 34802 52834
rect 35870 52782 35922 52834
rect 37998 52782 38050 52834
rect 40014 52782 40066 52834
rect 41694 52782 41746 52834
rect 44270 52782 44322 52834
rect 44606 52782 44658 52834
rect 47854 52782 47906 52834
rect 50206 52782 50258 52834
rect 51102 52782 51154 52834
rect 52110 52782 52162 52834
rect 52446 52782 52498 52834
rect 54350 52782 54402 52834
rect 56590 52782 56642 52834
rect 58382 52782 58434 52834
rect 58942 52782 58994 52834
rect 60286 52782 60338 52834
rect 61294 52782 61346 52834
rect 61966 52782 62018 52834
rect 10110 52670 10162 52722
rect 11342 52670 11394 52722
rect 15150 52670 15202 52722
rect 21422 52670 21474 52722
rect 31614 52670 31666 52722
rect 34190 52670 34242 52722
rect 38446 52670 38498 52722
rect 38782 52670 38834 52722
rect 43822 52670 43874 52722
rect 45614 52670 45666 52722
rect 55582 52670 55634 52722
rect 55918 52670 55970 52722
rect 57150 52670 57202 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 7870 52334 7922 52386
rect 8318 52334 8370 52386
rect 23102 52334 23154 52386
rect 37102 52334 37154 52386
rect 50094 52334 50146 52386
rect 6862 52222 6914 52274
rect 8318 52222 8370 52274
rect 9102 52222 9154 52274
rect 9550 52222 9602 52274
rect 14366 52222 14418 52274
rect 15262 52222 15314 52274
rect 15710 52222 15762 52274
rect 17614 52222 17666 52274
rect 19742 52222 19794 52274
rect 22206 52222 22258 52274
rect 23326 52222 23378 52274
rect 23998 52222 24050 52274
rect 28254 52222 28306 52274
rect 32734 52222 32786 52274
rect 43150 52222 43202 52274
rect 44270 52222 44322 52274
rect 45390 52222 45442 52274
rect 47294 52222 47346 52274
rect 55694 52222 55746 52274
rect 58270 52222 58322 52274
rect 60734 52222 60786 52274
rect 61070 52222 61122 52274
rect 61518 52222 61570 52274
rect 7422 52110 7474 52162
rect 10110 52110 10162 52162
rect 13694 52110 13746 52162
rect 13806 52110 13858 52162
rect 15150 52110 15202 52162
rect 15822 52110 15874 52162
rect 16046 52110 16098 52162
rect 20526 52110 20578 52162
rect 21198 52110 21250 52162
rect 21870 52110 21922 52162
rect 23662 52110 23714 52162
rect 24334 52110 24386 52162
rect 25342 52110 25394 52162
rect 29934 52110 29986 52162
rect 32174 52110 32226 52162
rect 32510 52110 32562 52162
rect 32846 52110 32898 52162
rect 34862 52110 34914 52162
rect 35086 52110 35138 52162
rect 35422 52110 35474 52162
rect 35758 52110 35810 52162
rect 36206 52110 36258 52162
rect 36990 52110 37042 52162
rect 40350 52110 40402 52162
rect 43710 52110 43762 52162
rect 45166 52110 45218 52162
rect 45726 52110 45778 52162
rect 45950 52110 46002 52162
rect 46734 52110 46786 52162
rect 48302 52110 48354 52162
rect 48862 52110 48914 52162
rect 49982 52110 50034 52162
rect 51886 52110 51938 52162
rect 52558 52110 52610 52162
rect 52782 52110 52834 52162
rect 52894 52110 52946 52162
rect 53118 52110 53170 52162
rect 53454 52110 53506 52162
rect 53902 52110 53954 52162
rect 54798 52110 54850 52162
rect 55470 52110 55522 52162
rect 57710 52110 57762 52162
rect 58830 52110 58882 52162
rect 59614 52110 59666 52162
rect 11678 51998 11730 52050
rect 12574 51998 12626 52050
rect 12910 51998 12962 52050
rect 14478 51998 14530 52050
rect 17278 51998 17330 52050
rect 21534 51998 21586 52050
rect 24222 51998 24274 52050
rect 24558 51998 24610 52050
rect 24782 51998 24834 52050
rect 26126 51998 26178 52050
rect 29150 51998 29202 52050
rect 30270 51998 30322 52050
rect 30382 51998 30434 52050
rect 30606 51998 30658 52050
rect 31838 51998 31890 52050
rect 34638 51998 34690 52050
rect 38446 51998 38498 52050
rect 41022 51998 41074 52050
rect 43486 51998 43538 52050
rect 48078 51998 48130 52050
rect 51550 51998 51602 52050
rect 54126 51998 54178 52050
rect 7870 51886 7922 51938
rect 8766 51886 8818 51938
rect 10446 51886 10498 51938
rect 14254 51886 14306 51938
rect 16942 51886 16994 51938
rect 21422 51886 21474 51938
rect 29262 51886 29314 51938
rect 30494 51886 30546 51938
rect 35422 51886 35474 51938
rect 39790 51886 39842 51938
rect 44830 51886 44882 51938
rect 46286 51886 46338 51938
rect 47742 51886 47794 51938
rect 53678 51886 53730 51938
rect 58830 51886 58882 51938
rect 60062 51886 60114 51938
rect 61966 51886 62018 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 4846 51550 4898 51602
rect 5854 51550 5906 51602
rect 7198 51550 7250 51602
rect 8206 51550 8258 51602
rect 8654 51550 8706 51602
rect 10222 51550 10274 51602
rect 13470 51550 13522 51602
rect 17502 51550 17554 51602
rect 18958 51550 19010 51602
rect 20078 51550 20130 51602
rect 23438 51550 23490 51602
rect 25230 51550 25282 51602
rect 26350 51550 26402 51602
rect 26574 51550 26626 51602
rect 27806 51550 27858 51602
rect 28926 51550 28978 51602
rect 29374 51550 29426 51602
rect 29598 51550 29650 51602
rect 32398 51550 32450 51602
rect 39790 51550 39842 51602
rect 40238 51550 40290 51602
rect 43150 51550 43202 51602
rect 44718 51550 44770 51602
rect 44942 51550 44994 51602
rect 45838 51550 45890 51602
rect 47742 51550 47794 51602
rect 61294 51550 61346 51602
rect 17390 51438 17442 51490
rect 18286 51438 18338 51490
rect 21534 51438 21586 51490
rect 24558 51438 24610 51490
rect 30270 51438 30322 51490
rect 31614 51438 31666 51490
rect 33966 51438 34018 51490
rect 36766 51438 36818 51490
rect 38110 51438 38162 51490
rect 38334 51438 38386 51490
rect 39454 51438 39506 51490
rect 41918 51438 41970 51490
rect 44606 51438 44658 51490
rect 53342 51438 53394 51490
rect 60846 51438 60898 51490
rect 13358 51326 13410 51378
rect 13694 51326 13746 51378
rect 14030 51326 14082 51378
rect 17950 51326 18002 51378
rect 18846 51326 18898 51378
rect 22990 51326 23042 51378
rect 23774 51326 23826 51378
rect 24446 51326 24498 51378
rect 25454 51326 25506 51378
rect 26686 51326 26738 51378
rect 26798 51326 26850 51378
rect 29822 51326 29874 51378
rect 31278 51326 31330 51378
rect 32062 51326 32114 51378
rect 32174 51326 32226 51378
rect 32510 51326 32562 51378
rect 33518 51326 33570 51378
rect 34974 51326 35026 51378
rect 36430 51326 36482 51378
rect 37102 51326 37154 51378
rect 38670 51326 38722 51378
rect 43822 51326 43874 51378
rect 49198 51326 49250 51378
rect 53566 51326 53618 51378
rect 54350 51326 54402 51378
rect 54574 51326 54626 51378
rect 57038 51326 57090 51378
rect 2942 51214 2994 51266
rect 4174 51214 4226 51266
rect 6414 51214 6466 51266
rect 6862 51214 6914 51266
rect 7646 51214 7698 51266
rect 9102 51214 9154 51266
rect 12686 51214 12738 51266
rect 12910 51214 12962 51266
rect 14702 51214 14754 51266
rect 16830 51214 16882 51266
rect 22654 51214 22706 51266
rect 29710 51214 29762 51266
rect 41022 51214 41074 51266
rect 44270 51214 44322 51266
rect 48974 51214 49026 51266
rect 49982 51214 50034 51266
rect 52110 51214 52162 51266
rect 56702 51214 56754 51266
rect 57822 51214 57874 51266
rect 59950 51214 60002 51266
rect 60398 51214 60450 51266
rect 61742 51214 61794 51266
rect 62190 51214 62242 51266
rect 12126 51102 12178 51154
rect 17502 51102 17554 51154
rect 30606 51102 30658 51154
rect 33630 51102 33682 51154
rect 37102 51102 37154 51154
rect 39006 51102 39058 51154
rect 55022 51102 55074 51154
rect 60398 51102 60450 51154
rect 61966 51102 62018 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 3614 50766 3666 50818
rect 4510 50766 4562 50818
rect 22542 50766 22594 50818
rect 22878 50766 22930 50818
rect 24334 50766 24386 50818
rect 34526 50766 34578 50818
rect 36094 50766 36146 50818
rect 47630 50766 47682 50818
rect 49422 50766 49474 50818
rect 50878 50766 50930 50818
rect 60510 50766 60562 50818
rect 61294 50766 61346 50818
rect 6190 50654 6242 50706
rect 7870 50654 7922 50706
rect 15822 50654 15874 50706
rect 31390 50654 31442 50706
rect 33518 50654 33570 50706
rect 34750 50654 34802 50706
rect 36318 50654 36370 50706
rect 39790 50654 39842 50706
rect 40350 50654 40402 50706
rect 41694 50654 41746 50706
rect 46398 50654 46450 50706
rect 47518 50654 47570 50706
rect 49758 50654 49810 50706
rect 53230 50654 53282 50706
rect 59950 50654 60002 50706
rect 60622 50654 60674 50706
rect 61518 50654 61570 50706
rect 61966 50654 62018 50706
rect 5182 50542 5234 50594
rect 7086 50542 7138 50594
rect 9326 50542 9378 50594
rect 9886 50542 9938 50594
rect 10110 50542 10162 50594
rect 13022 50542 13074 50594
rect 13806 50542 13858 50594
rect 14366 50542 14418 50594
rect 15150 50542 15202 50594
rect 15486 50542 15538 50594
rect 15934 50542 15986 50594
rect 20526 50542 20578 50594
rect 21870 50542 21922 50594
rect 23326 50542 23378 50594
rect 24446 50542 24498 50594
rect 25790 50542 25842 50594
rect 26238 50542 26290 50594
rect 28030 50542 28082 50594
rect 28590 50542 28642 50594
rect 29710 50542 29762 50594
rect 30606 50542 30658 50594
rect 30942 50542 30994 50594
rect 33406 50542 33458 50594
rect 34638 50542 34690 50594
rect 35086 50542 35138 50594
rect 35310 50542 35362 50594
rect 40014 50542 40066 50594
rect 41246 50542 41298 50594
rect 42478 50542 42530 50594
rect 42702 50542 42754 50594
rect 43262 50542 43314 50594
rect 43710 50542 43762 50594
rect 44270 50542 44322 50594
rect 45950 50542 46002 50594
rect 47182 50542 47234 50594
rect 48078 50542 48130 50594
rect 48526 50542 48578 50594
rect 49198 50542 49250 50594
rect 50318 50542 50370 50594
rect 50654 50542 50706 50594
rect 50990 50542 51042 50594
rect 51438 50542 51490 50594
rect 51662 50542 51714 50594
rect 53006 50542 53058 50594
rect 54238 50542 54290 50594
rect 55246 50542 55298 50594
rect 55694 50542 55746 50594
rect 58046 50542 58098 50594
rect 58718 50542 58770 50594
rect 59390 50542 59442 50594
rect 3614 50430 3666 50482
rect 4398 50430 4450 50482
rect 6638 50430 6690 50482
rect 8430 50430 8482 50482
rect 8654 50430 8706 50482
rect 8766 50430 8818 50482
rect 8990 50430 9042 50482
rect 9550 50430 9602 50482
rect 11230 50430 11282 50482
rect 13582 50430 13634 50482
rect 15262 50430 15314 50482
rect 15710 50430 15762 50482
rect 16158 50430 16210 50482
rect 18734 50430 18786 50482
rect 20638 50430 20690 50482
rect 20750 50430 20802 50482
rect 21758 50430 21810 50482
rect 25006 50430 25058 50482
rect 29374 50430 29426 50482
rect 37326 50430 37378 50482
rect 40798 50430 40850 50482
rect 41022 50430 41074 50482
rect 43038 50430 43090 50482
rect 45054 50430 45106 50482
rect 45838 50430 45890 50482
rect 48414 50430 48466 50482
rect 49758 50430 49810 50482
rect 49982 50430 50034 50482
rect 51886 50430 51938 50482
rect 56926 50430 56978 50482
rect 58494 50430 58546 50482
rect 59166 50430 59218 50482
rect 61182 50430 61234 50482
rect 1934 50318 1986 50370
rect 2382 50318 2434 50370
rect 2830 50318 2882 50370
rect 4062 50318 4114 50370
rect 7534 50318 7586 50370
rect 10446 50318 10498 50370
rect 14702 50318 14754 50370
rect 16830 50318 16882 50370
rect 19966 50318 20018 50370
rect 20302 50318 20354 50370
rect 23662 50318 23714 50370
rect 35758 50318 35810 50370
rect 39118 50318 39170 50370
rect 41134 50318 41186 50370
rect 42142 50318 42194 50370
rect 45166 50318 45218 50370
rect 50430 50318 50482 50370
rect 51550 50318 51602 50370
rect 57822 50318 57874 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 3054 49982 3106 50034
rect 5966 49982 6018 50034
rect 6414 49982 6466 50034
rect 6750 49982 6802 50034
rect 7310 49982 7362 50034
rect 8094 49982 8146 50034
rect 10222 49982 10274 50034
rect 11566 49982 11618 50034
rect 16718 49982 16770 50034
rect 25678 49982 25730 50034
rect 27134 49982 27186 50034
rect 30718 49982 30770 50034
rect 30830 49982 30882 50034
rect 31278 49982 31330 50034
rect 33406 49982 33458 50034
rect 38446 49982 38498 50034
rect 49758 49982 49810 50034
rect 51214 49982 51266 50034
rect 51438 49982 51490 50034
rect 54798 49982 54850 50034
rect 56590 49982 56642 50034
rect 61854 49982 61906 50034
rect 2382 49870 2434 49922
rect 3390 49870 3442 49922
rect 12686 49870 12738 49922
rect 16382 49870 16434 49922
rect 16494 49870 16546 49922
rect 16606 49870 16658 49922
rect 18398 49870 18450 49922
rect 21422 49870 21474 49922
rect 22430 49870 22482 49922
rect 30270 49870 30322 49922
rect 30494 49870 30546 49922
rect 30606 49870 30658 49922
rect 31950 49870 32002 49922
rect 32398 49870 32450 49922
rect 33070 49870 33122 49922
rect 33182 49870 33234 49922
rect 33742 49870 33794 49922
rect 36654 49870 36706 49922
rect 38894 49870 38946 49922
rect 40350 49870 40402 49922
rect 48862 49870 48914 49922
rect 51662 49870 51714 49922
rect 51774 49870 51826 49922
rect 52894 49870 52946 49922
rect 55694 49870 55746 49922
rect 2718 49758 2770 49810
rect 8430 49758 8482 49810
rect 8654 49758 8706 49810
rect 9102 49758 9154 49810
rect 12462 49758 12514 49810
rect 13246 49758 13298 49810
rect 13918 49758 13970 49810
rect 14366 49758 14418 49810
rect 14590 49758 14642 49810
rect 15710 49758 15762 49810
rect 16830 49758 16882 49810
rect 19518 49758 19570 49810
rect 20302 49758 20354 49810
rect 21758 49758 21810 49810
rect 22766 49758 22818 49810
rect 24110 49758 24162 49810
rect 25230 49758 25282 49810
rect 25566 49758 25618 49810
rect 25790 49758 25842 49810
rect 31614 49758 31666 49810
rect 34190 49758 34242 49810
rect 34750 49758 34802 49810
rect 35534 49758 35586 49810
rect 39902 49758 39954 49810
rect 41022 49758 41074 49810
rect 42142 49758 42194 49810
rect 42814 49758 42866 49810
rect 43598 49758 43650 49810
rect 44830 49758 44882 49810
rect 45726 49758 45778 49810
rect 47406 49758 47458 49810
rect 47742 49758 47794 49810
rect 49198 49758 49250 49810
rect 49646 49758 49698 49810
rect 50430 49758 50482 49810
rect 50766 49758 50818 49810
rect 50990 49758 51042 49810
rect 54238 49758 54290 49810
rect 55806 49758 55858 49810
rect 56926 49758 56978 49810
rect 57150 49758 57202 49810
rect 58046 49758 58098 49810
rect 58270 49758 58322 49810
rect 58718 49758 58770 49810
rect 58942 49758 58994 49810
rect 59838 49758 59890 49810
rect 61294 49758 61346 49810
rect 1822 49646 1874 49698
rect 3950 49646 4002 49698
rect 4510 49646 4562 49698
rect 4958 49646 5010 49698
rect 5518 49646 5570 49698
rect 7758 49646 7810 49698
rect 8878 49646 8930 49698
rect 14478 49646 14530 49698
rect 15486 49646 15538 49698
rect 24670 49646 24722 49698
rect 29822 49646 29874 49698
rect 45502 49646 45554 49698
rect 57486 49646 57538 49698
rect 58494 49646 58546 49698
rect 59390 49646 59442 49698
rect 60286 49646 60338 49698
rect 60846 49646 60898 49698
rect 1822 49534 1874 49586
rect 2158 49534 2210 49586
rect 13582 49534 13634 49586
rect 19966 49534 20018 49586
rect 29038 49534 29090 49586
rect 38782 49534 38834 49586
rect 39342 49534 39394 49586
rect 39678 49534 39730 49586
rect 44158 49534 44210 49586
rect 50878 49534 50930 49586
rect 55134 49534 55186 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 11006 49198 11058 49250
rect 21310 49198 21362 49250
rect 21758 49198 21810 49250
rect 30942 49198 30994 49250
rect 34974 49198 35026 49250
rect 42702 49198 42754 49250
rect 48078 49198 48130 49250
rect 51438 49198 51490 49250
rect 54574 49198 54626 49250
rect 4510 49086 4562 49138
rect 5630 49086 5682 49138
rect 6862 49086 6914 49138
rect 10110 49086 10162 49138
rect 10446 49086 10498 49138
rect 11342 49086 11394 49138
rect 21422 49086 21474 49138
rect 27694 49086 27746 49138
rect 32622 49086 32674 49138
rect 35870 49086 35922 49138
rect 37102 49086 37154 49138
rect 44046 49086 44098 49138
rect 45950 49086 46002 49138
rect 47070 49086 47122 49138
rect 49310 49086 49362 49138
rect 52782 49086 52834 49138
rect 58382 49086 58434 49138
rect 59278 49086 59330 49138
rect 59950 49086 60002 49138
rect 60510 49086 60562 49138
rect 2494 48974 2546 49026
rect 4062 48974 4114 49026
rect 4734 48974 4786 49026
rect 5854 48974 5906 49026
rect 7198 48974 7250 49026
rect 10670 48974 10722 49026
rect 11678 48974 11730 49026
rect 12126 48974 12178 49026
rect 14142 48974 14194 49026
rect 14366 48974 14418 49026
rect 15598 48974 15650 49026
rect 17614 48974 17666 49026
rect 18510 48974 18562 49026
rect 19742 48974 19794 49026
rect 20078 48974 20130 49026
rect 22094 48974 22146 49026
rect 22766 48974 22818 49026
rect 24110 48974 24162 49026
rect 24446 48974 24498 49026
rect 28254 48974 28306 49026
rect 29598 48974 29650 49026
rect 30046 48974 30098 49026
rect 31502 48974 31554 49026
rect 32286 48974 32338 49026
rect 34302 48974 34354 49026
rect 35646 48974 35698 49026
rect 36206 48974 36258 49026
rect 36878 48974 36930 49026
rect 37438 48974 37490 49026
rect 38110 48974 38162 49026
rect 38558 48974 38610 49026
rect 39342 48974 39394 49026
rect 40574 48974 40626 49026
rect 42366 48974 42418 49026
rect 43486 48974 43538 49026
rect 46958 48974 47010 49026
rect 47182 48974 47234 49026
rect 48974 48974 49026 49026
rect 49870 48974 49922 49026
rect 50206 48974 50258 49026
rect 50766 48974 50818 49026
rect 52894 48974 52946 49026
rect 53790 48974 53842 49026
rect 58158 48974 58210 49026
rect 59054 48974 59106 49026
rect 59614 48974 59666 49026
rect 60734 48974 60786 49026
rect 61630 48974 61682 49026
rect 2046 48862 2098 48914
rect 2718 48862 2770 48914
rect 3502 48862 3554 48914
rect 7982 48862 8034 48914
rect 11566 48862 11618 48914
rect 12910 48862 12962 48914
rect 14814 48862 14866 48914
rect 15262 48862 15314 48914
rect 16942 48862 16994 48914
rect 17950 48862 18002 48914
rect 20638 48862 20690 48914
rect 22318 48862 22370 48914
rect 24558 48862 24610 48914
rect 26686 48862 26738 48914
rect 28030 48862 28082 48914
rect 30942 48862 30994 48914
rect 34414 48862 34466 48914
rect 36094 48862 36146 48914
rect 37326 48862 37378 48914
rect 39454 48862 39506 48914
rect 41134 48862 41186 48914
rect 43262 48862 43314 48914
rect 45278 48862 45330 48914
rect 45726 48862 45778 48914
rect 47742 48862 47794 48914
rect 48190 48862 48242 48914
rect 48750 48862 48802 48914
rect 50654 48862 50706 48914
rect 54014 48862 54066 48914
rect 56814 48862 56866 48914
rect 1710 48750 1762 48802
rect 3166 48750 3218 48802
rect 4174 48750 4226 48802
rect 5070 48750 5122 48802
rect 6190 48750 6242 48802
rect 11902 48750 11954 48802
rect 12574 48750 12626 48802
rect 13806 48750 13858 48802
rect 15934 48750 15986 48802
rect 25454 48750 25506 48802
rect 28590 48750 28642 48802
rect 35310 48750 35362 48802
rect 37886 48750 37938 48802
rect 38894 48750 38946 48802
rect 44942 48750 44994 48802
rect 47966 48750 48018 48802
rect 51774 48750 51826 48802
rect 54910 48750 54962 48802
rect 55470 48750 55522 48802
rect 57822 48750 57874 48802
rect 58718 48750 58770 48802
rect 61070 48750 61122 48802
rect 61742 48750 61794 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 1710 48414 1762 48466
rect 4174 48414 4226 48466
rect 4958 48414 5010 48466
rect 8094 48414 8146 48466
rect 8766 48414 8818 48466
rect 12798 48414 12850 48466
rect 23326 48414 23378 48466
rect 24334 48414 24386 48466
rect 27246 48414 27298 48466
rect 31614 48414 31666 48466
rect 36542 48414 36594 48466
rect 37662 48414 37714 48466
rect 40126 48414 40178 48466
rect 54350 48414 54402 48466
rect 56702 48414 56754 48466
rect 3054 48302 3106 48354
rect 4622 48302 4674 48354
rect 5742 48302 5794 48354
rect 10670 48302 10722 48354
rect 13134 48302 13186 48354
rect 22206 48302 22258 48354
rect 30046 48302 30098 48354
rect 30606 48302 30658 48354
rect 31054 48302 31106 48354
rect 33182 48302 33234 48354
rect 33742 48302 33794 48354
rect 35310 48302 35362 48354
rect 35758 48302 35810 48354
rect 36654 48302 36706 48354
rect 36766 48302 36818 48354
rect 40014 48302 40066 48354
rect 41582 48302 41634 48354
rect 44158 48302 44210 48354
rect 47742 48302 47794 48354
rect 49982 48302 50034 48354
rect 50878 48302 50930 48354
rect 52446 48302 52498 48354
rect 59614 48302 59666 48354
rect 62078 48302 62130 48354
rect 1934 48190 1986 48242
rect 5294 48190 5346 48242
rect 6302 48190 6354 48242
rect 6750 48190 6802 48242
rect 8318 48190 8370 48242
rect 8990 48190 9042 48242
rect 13582 48190 13634 48242
rect 14702 48190 14754 48242
rect 15374 48190 15426 48242
rect 16606 48190 16658 48242
rect 18062 48190 18114 48242
rect 18286 48190 18338 48242
rect 20078 48190 20130 48242
rect 20526 48190 20578 48242
rect 23774 48190 23826 48242
rect 23998 48190 24050 48242
rect 28590 48190 28642 48242
rect 29038 48190 29090 48242
rect 29822 48190 29874 48242
rect 31278 48190 31330 48242
rect 33070 48190 33122 48242
rect 34302 48190 34354 48242
rect 34862 48190 34914 48242
rect 36094 48190 36146 48242
rect 36430 48190 36482 48242
rect 37214 48190 37266 48242
rect 37438 48190 37490 48242
rect 37774 48190 37826 48242
rect 38110 48190 38162 48242
rect 39566 48190 39618 48242
rect 40350 48190 40402 48242
rect 41134 48190 41186 48242
rect 42030 48190 42082 48242
rect 42590 48190 42642 48242
rect 44606 48190 44658 48242
rect 45502 48190 45554 48242
rect 47070 48190 47122 48242
rect 47630 48190 47682 48242
rect 49422 48190 49474 48242
rect 50654 48190 50706 48242
rect 51214 48190 51266 48242
rect 51438 48190 51490 48242
rect 51774 48190 51826 48242
rect 54574 48190 54626 48242
rect 54798 48190 54850 48242
rect 55246 48190 55298 48242
rect 55470 48190 55522 48242
rect 57150 48190 57202 48242
rect 57710 48190 57762 48242
rect 57934 48190 57986 48242
rect 58270 48190 58322 48242
rect 58494 48190 58546 48242
rect 58942 48190 58994 48242
rect 61854 48190 61906 48242
rect 8878 48078 8930 48130
rect 9550 48078 9602 48130
rect 9774 48078 9826 48130
rect 21086 48078 21138 48130
rect 25342 48078 25394 48130
rect 32622 48078 32674 48130
rect 33854 48078 33906 48130
rect 38446 48078 38498 48130
rect 38782 48078 38834 48130
rect 39230 48078 39282 48130
rect 40014 48078 40066 48130
rect 41470 48078 41522 48130
rect 43038 48078 43090 48130
rect 45614 48078 45666 48130
rect 48078 48078 48130 48130
rect 48862 48078 48914 48130
rect 49870 48078 49922 48130
rect 51326 48078 51378 48130
rect 54686 48078 54738 48130
rect 57822 48078 57874 48130
rect 58382 48078 58434 48130
rect 12462 47966 12514 48018
rect 16718 47966 16770 48018
rect 25902 47966 25954 48018
rect 28926 47966 28978 48018
rect 46286 47966 46338 48018
rect 56030 47966 56082 48018
rect 57374 47966 57426 48018
rect 61518 47966 61570 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 8542 47630 8594 47682
rect 24110 47630 24162 47682
rect 26574 47630 26626 47682
rect 30942 47630 30994 47682
rect 33630 47630 33682 47682
rect 35646 47630 35698 47682
rect 41582 47630 41634 47682
rect 46062 47630 46114 47682
rect 51774 47630 51826 47682
rect 53566 47630 53618 47682
rect 59278 47630 59330 47682
rect 61966 47630 62018 47682
rect 4622 47518 4674 47570
rect 9214 47518 9266 47570
rect 16158 47518 16210 47570
rect 19854 47518 19906 47570
rect 22542 47518 22594 47570
rect 23662 47518 23714 47570
rect 27806 47518 27858 47570
rect 37998 47518 38050 47570
rect 43038 47518 43090 47570
rect 51326 47518 51378 47570
rect 53118 47518 53170 47570
rect 53678 47518 53730 47570
rect 60958 47518 61010 47570
rect 1710 47406 1762 47458
rect 9326 47406 9378 47458
rect 10334 47406 10386 47458
rect 10558 47406 10610 47458
rect 11230 47406 11282 47458
rect 12014 47406 12066 47458
rect 12686 47406 12738 47458
rect 14030 47406 14082 47458
rect 14254 47406 14306 47458
rect 15486 47406 15538 47458
rect 16046 47406 16098 47458
rect 16494 47406 16546 47458
rect 17502 47406 17554 47458
rect 19966 47406 20018 47458
rect 20302 47406 20354 47458
rect 21310 47406 21362 47458
rect 24446 47406 24498 47458
rect 25790 47406 25842 47458
rect 29374 47406 29426 47458
rect 30606 47406 30658 47458
rect 31502 47406 31554 47458
rect 33294 47406 33346 47458
rect 34302 47406 34354 47458
rect 35086 47406 35138 47458
rect 35310 47406 35362 47458
rect 35870 47406 35922 47458
rect 37662 47406 37714 47458
rect 41806 47406 41858 47458
rect 43822 47406 43874 47458
rect 45838 47406 45890 47458
rect 47518 47406 47570 47458
rect 48862 47406 48914 47458
rect 49534 47406 49586 47458
rect 51438 47406 51490 47458
rect 52110 47406 52162 47458
rect 55022 47406 55074 47458
rect 55470 47406 55522 47458
rect 56366 47406 56418 47458
rect 56814 47406 56866 47458
rect 57598 47406 57650 47458
rect 58494 47406 58546 47458
rect 58942 47406 58994 47458
rect 59726 47406 59778 47458
rect 60622 47406 60674 47458
rect 60734 47406 60786 47458
rect 2494 47294 2546 47346
rect 4958 47294 5010 47346
rect 6526 47294 6578 47346
rect 9214 47294 9266 47346
rect 12798 47294 12850 47346
rect 13582 47294 13634 47346
rect 14702 47294 14754 47346
rect 15374 47294 15426 47346
rect 16270 47294 16322 47346
rect 16606 47294 16658 47346
rect 18062 47294 18114 47346
rect 21422 47294 21474 47346
rect 21982 47294 22034 47346
rect 23326 47294 23378 47346
rect 24782 47294 24834 47346
rect 25006 47294 25058 47346
rect 26014 47294 26066 47346
rect 26910 47294 26962 47346
rect 28142 47294 28194 47346
rect 28254 47294 28306 47346
rect 28366 47294 28418 47346
rect 28590 47294 28642 47346
rect 31950 47294 32002 47346
rect 33070 47294 33122 47346
rect 34078 47294 34130 47346
rect 37214 47294 37266 47346
rect 39118 47294 39170 47346
rect 42590 47294 42642 47346
rect 42702 47294 42754 47346
rect 43374 47294 43426 47346
rect 43486 47294 43538 47346
rect 43598 47294 43650 47346
rect 46174 47294 46226 47346
rect 49982 47294 50034 47346
rect 50094 47294 50146 47346
rect 50206 47294 50258 47346
rect 50878 47294 50930 47346
rect 51102 47294 51154 47346
rect 55806 47294 55858 47346
rect 56926 47294 56978 47346
rect 62190 47294 62242 47346
rect 5070 47182 5122 47234
rect 10894 47182 10946 47234
rect 11118 47182 11170 47234
rect 11902 47182 11954 47234
rect 13470 47182 13522 47234
rect 22990 47182 23042 47234
rect 27582 47182 27634 47234
rect 35422 47182 35474 47234
rect 36318 47182 36370 47234
rect 40574 47182 40626 47234
rect 42366 47182 42418 47234
rect 44270 47182 44322 47234
rect 44830 47182 44882 47234
rect 45166 47182 45218 47234
rect 50318 47182 50370 47234
rect 51214 47182 51266 47234
rect 51886 47182 51938 47234
rect 52670 47182 52722 47234
rect 57934 47182 57986 47234
rect 60622 47182 60674 47234
rect 61630 47182 61682 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 5294 46846 5346 46898
rect 8542 46846 8594 46898
rect 12798 46846 12850 46898
rect 13022 46846 13074 46898
rect 13134 46846 13186 46898
rect 13246 46846 13298 46898
rect 18622 46846 18674 46898
rect 27470 46846 27522 46898
rect 38222 46846 38274 46898
rect 42254 46846 42306 46898
rect 43822 46846 43874 46898
rect 44046 46846 44098 46898
rect 45726 46846 45778 46898
rect 45838 46846 45890 46898
rect 45950 46846 46002 46898
rect 46398 46846 46450 46898
rect 49310 46846 49362 46898
rect 50430 46846 50482 46898
rect 53342 46846 53394 46898
rect 53678 46846 53730 46898
rect 2270 46734 2322 46786
rect 3614 46734 3666 46786
rect 3950 46734 4002 46786
rect 6638 46734 6690 46786
rect 6862 46734 6914 46786
rect 8430 46734 8482 46786
rect 10446 46734 10498 46786
rect 10670 46734 10722 46786
rect 10782 46734 10834 46786
rect 11790 46734 11842 46786
rect 14478 46734 14530 46786
rect 15374 46734 15426 46786
rect 15934 46734 15986 46786
rect 17726 46734 17778 46786
rect 17950 46734 18002 46786
rect 19742 46734 19794 46786
rect 22878 46734 22930 46786
rect 23998 46734 24050 46786
rect 24558 46734 24610 46786
rect 25566 46734 25618 46786
rect 28814 46734 28866 46786
rect 31614 46734 31666 46786
rect 32174 46734 32226 46786
rect 32510 46734 32562 46786
rect 33406 46734 33458 46786
rect 33854 46734 33906 46786
rect 40910 46734 40962 46786
rect 42814 46734 42866 46786
rect 43374 46734 43426 46786
rect 45390 46734 45442 46786
rect 45614 46734 45666 46786
rect 47518 46734 47570 46786
rect 48078 46734 48130 46786
rect 48190 46734 48242 46786
rect 49422 46734 49474 46786
rect 49870 46734 49922 46786
rect 51550 46734 51602 46786
rect 53902 46734 53954 46786
rect 54462 46734 54514 46786
rect 56702 46734 56754 46786
rect 56814 46734 56866 46786
rect 57486 46734 57538 46786
rect 2494 46622 2546 46674
rect 2718 46622 2770 46674
rect 3838 46622 3890 46674
rect 6078 46622 6130 46674
rect 7310 46622 7362 46674
rect 8318 46622 8370 46674
rect 9550 46622 9602 46674
rect 9774 46622 9826 46674
rect 13806 46622 13858 46674
rect 14702 46622 14754 46674
rect 16158 46622 16210 46674
rect 19294 46622 19346 46674
rect 21086 46622 21138 46674
rect 22766 46622 22818 46674
rect 22990 46622 23042 46674
rect 23326 46622 23378 46674
rect 23774 46622 23826 46674
rect 24334 46622 24386 46674
rect 27806 46622 27858 46674
rect 28590 46622 28642 46674
rect 29710 46622 29762 46674
rect 29934 46622 29986 46674
rect 31390 46622 31442 46674
rect 33630 46622 33682 46674
rect 34190 46622 34242 46674
rect 40014 46622 40066 46674
rect 42590 46622 42642 46674
rect 44382 46622 44434 46674
rect 44830 46622 44882 46674
rect 46734 46622 46786 46674
rect 47294 46622 47346 46674
rect 48974 46622 49026 46674
rect 50542 46622 50594 46674
rect 54798 46622 54850 46674
rect 55246 46622 55298 46674
rect 55694 46622 55746 46674
rect 58158 46622 58210 46674
rect 59054 46622 59106 46674
rect 60286 46622 60338 46674
rect 61518 46622 61570 46674
rect 61966 46622 62018 46674
rect 62190 46622 62242 46674
rect 1934 46510 1986 46562
rect 2606 46510 2658 46562
rect 4510 46510 4562 46562
rect 4846 46510 4898 46562
rect 6302 46510 6354 46562
rect 8766 46510 8818 46562
rect 14030 46510 14082 46562
rect 16270 46510 16322 46562
rect 16494 46510 16546 46562
rect 16830 46510 16882 46562
rect 18286 46510 18338 46562
rect 21310 46510 21362 46562
rect 24670 46510 24722 46562
rect 28142 46510 28194 46562
rect 33742 46510 33794 46562
rect 34974 46510 35026 46562
rect 37102 46510 37154 46562
rect 43934 46510 43986 46562
rect 54350 46510 54402 46562
rect 57262 46510 57314 46562
rect 61294 46510 61346 46562
rect 61742 46510 61794 46562
rect 3166 46398 3218 46450
rect 3390 46398 3442 46450
rect 8990 46398 9042 46450
rect 10110 46398 10162 46450
rect 11006 46398 11058 46450
rect 11230 46398 11282 46450
rect 12014 46398 12066 46450
rect 12350 46398 12402 46450
rect 21422 46398 21474 46450
rect 41134 46398 41186 46450
rect 41470 46398 41522 46450
rect 48078 46398 48130 46450
rect 53566 46398 53618 46450
rect 56702 46398 56754 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 7422 46062 7474 46114
rect 9774 46062 9826 46114
rect 9998 46062 10050 46114
rect 11790 46062 11842 46114
rect 18174 46062 18226 46114
rect 24782 46062 24834 46114
rect 28254 46062 28306 46114
rect 28590 46062 28642 46114
rect 37102 46062 37154 46114
rect 39678 46062 39730 46114
rect 46062 46062 46114 46114
rect 55694 46062 55746 46114
rect 5742 45950 5794 46002
rect 8654 45950 8706 46002
rect 11342 45950 11394 46002
rect 18958 45950 19010 46002
rect 20078 45950 20130 46002
rect 24222 45950 24274 46002
rect 28030 45950 28082 46002
rect 29598 45950 29650 46002
rect 30382 45950 30434 46002
rect 31278 45950 31330 46002
rect 44270 45950 44322 46002
rect 44942 45950 44994 46002
rect 47966 45950 48018 46002
rect 51550 45950 51602 46002
rect 55470 45950 55522 46002
rect 60622 45950 60674 46002
rect 5182 45838 5234 45890
rect 6078 45838 6130 45890
rect 8542 45838 8594 45890
rect 9214 45838 9266 45890
rect 10446 45838 10498 45890
rect 11230 45838 11282 45890
rect 11790 45838 11842 45890
rect 12350 45838 12402 45890
rect 13470 45838 13522 45890
rect 14366 45838 14418 45890
rect 15150 45838 15202 45890
rect 18622 45838 18674 45890
rect 18846 45838 18898 45890
rect 19742 45838 19794 45890
rect 21422 45838 21474 45890
rect 24558 45838 24610 45890
rect 25790 45838 25842 45890
rect 26014 45838 26066 45890
rect 26350 45838 26402 45890
rect 26798 45838 26850 45890
rect 27022 45838 27074 45890
rect 27470 45838 27522 45890
rect 29150 45838 29202 45890
rect 29486 45838 29538 45890
rect 29710 45838 29762 45890
rect 31166 45838 31218 45890
rect 35534 45838 35586 45890
rect 40238 45838 40290 45890
rect 41358 45838 41410 45890
rect 46846 45838 46898 45890
rect 47854 45838 47906 45890
rect 50094 45838 50146 45890
rect 50542 45838 50594 45890
rect 51326 45838 51378 45890
rect 53118 45838 53170 45890
rect 55582 45838 55634 45890
rect 56478 45838 56530 45890
rect 60510 45838 60562 45890
rect 61294 45838 61346 45890
rect 61966 45838 62018 45890
rect 62190 45838 62242 45890
rect 3054 45726 3106 45778
rect 4510 45726 4562 45778
rect 4734 45726 4786 45778
rect 6750 45726 6802 45778
rect 7198 45726 7250 45778
rect 8654 45726 8706 45778
rect 10558 45726 10610 45778
rect 11454 45726 11506 45778
rect 12910 45726 12962 45778
rect 14254 45726 14306 45778
rect 16718 45726 16770 45778
rect 22094 45726 22146 45778
rect 25118 45726 25170 45778
rect 25342 45726 25394 45778
rect 26574 45726 26626 45778
rect 30942 45726 30994 45778
rect 33966 45726 34018 45778
rect 34862 45726 34914 45778
rect 35198 45726 35250 45778
rect 38222 45726 38274 45778
rect 40350 45726 40402 45778
rect 42142 45726 42194 45778
rect 45390 45726 45442 45778
rect 46622 45726 46674 45778
rect 49758 45726 49810 45778
rect 53342 45726 53394 45778
rect 53902 45726 53954 45778
rect 57038 45726 57090 45778
rect 58718 45726 58770 45778
rect 60846 45726 60898 45778
rect 1822 45614 1874 45666
rect 4286 45614 4338 45666
rect 4846 45614 4898 45666
rect 7758 45614 7810 45666
rect 9662 45614 9714 45666
rect 20862 45614 20914 45666
rect 24558 45614 24610 45666
rect 26014 45614 26066 45666
rect 26686 45614 26738 45666
rect 27582 45614 27634 45666
rect 27806 45614 27858 45666
rect 31390 45614 31442 45666
rect 32398 45614 32450 45666
rect 33518 45614 33570 45666
rect 34302 45614 34354 45666
rect 35870 45614 35922 45666
rect 36542 45614 36594 45666
rect 39342 45614 39394 45666
rect 41134 45614 41186 45666
rect 50878 45614 50930 45666
rect 51886 45614 51938 45666
rect 52782 45614 52834 45666
rect 59838 45614 59890 45666
rect 60734 45614 60786 45666
rect 61630 45614 61682 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 4174 45278 4226 45330
rect 7086 45278 7138 45330
rect 7310 45278 7362 45330
rect 8542 45278 8594 45330
rect 10670 45278 10722 45330
rect 11230 45278 11282 45330
rect 12798 45278 12850 45330
rect 17390 45278 17442 45330
rect 17614 45278 17666 45330
rect 26350 45278 26402 45330
rect 35198 45278 35250 45330
rect 40238 45278 40290 45330
rect 40910 45278 40962 45330
rect 45726 45278 45778 45330
rect 46846 45278 46898 45330
rect 53790 45278 53842 45330
rect 2606 45166 2658 45218
rect 3166 45166 3218 45218
rect 6638 45166 6690 45218
rect 7422 45166 7474 45218
rect 8206 45166 8258 45218
rect 10558 45166 10610 45218
rect 10782 45166 10834 45218
rect 12238 45166 12290 45218
rect 17726 45166 17778 45218
rect 21758 45166 21810 45218
rect 23886 45166 23938 45218
rect 24110 45166 24162 45218
rect 28142 45166 28194 45218
rect 35646 45166 35698 45218
rect 36542 45166 36594 45218
rect 41694 45166 41746 45218
rect 43262 45166 43314 45218
rect 43822 45166 43874 45218
rect 43934 45166 43986 45218
rect 47630 45166 47682 45218
rect 48862 45166 48914 45218
rect 49982 45166 50034 45218
rect 53678 45166 53730 45218
rect 55918 45166 55970 45218
rect 56926 45166 56978 45218
rect 61630 45166 61682 45218
rect 2382 45054 2434 45106
rect 3054 45054 3106 45106
rect 5294 45054 5346 45106
rect 6302 45054 6354 45106
rect 7870 45054 7922 45106
rect 8430 45054 8482 45106
rect 8766 45054 8818 45106
rect 9550 45054 9602 45106
rect 11566 45054 11618 45106
rect 12350 45054 12402 45106
rect 13022 45054 13074 45106
rect 13582 45054 13634 45106
rect 14702 45054 14754 45106
rect 15374 45054 15426 45106
rect 16270 45054 16322 45106
rect 18062 45054 18114 45106
rect 20190 45054 20242 45106
rect 20638 45054 20690 45106
rect 21086 45054 21138 45106
rect 22878 45054 22930 45106
rect 23214 45054 23266 45106
rect 23438 45054 23490 45106
rect 23998 45054 24050 45106
rect 24670 45054 24722 45106
rect 26014 45054 26066 45106
rect 29262 45054 29314 45106
rect 33406 45054 33458 45106
rect 33742 45054 33794 45106
rect 37214 45054 37266 45106
rect 38110 45054 38162 45106
rect 39230 45054 39282 45106
rect 41134 45054 41186 45106
rect 42142 45054 42194 45106
rect 43038 45054 43090 45106
rect 43710 45054 43762 45106
rect 44494 45054 44546 45106
rect 47182 45054 47234 45106
rect 47742 45054 47794 45106
rect 48974 45054 49026 45106
rect 50318 45054 50370 45106
rect 51214 45054 51266 45106
rect 53342 45054 53394 45106
rect 54014 45054 54066 45106
rect 54798 45054 54850 45106
rect 55582 45054 55634 45106
rect 60174 45054 60226 45106
rect 60734 45054 60786 45106
rect 61182 45054 61234 45106
rect 2046 44942 2098 44994
rect 4846 44942 4898 44994
rect 5742 44942 5794 44994
rect 6526 44942 6578 44994
rect 7310 44942 7362 44994
rect 9998 44942 10050 44994
rect 17726 44942 17778 44994
rect 18622 44942 18674 44994
rect 22654 44942 22706 44994
rect 25678 44942 25730 44994
rect 30046 44942 30098 44994
rect 32174 44942 32226 44994
rect 33966 44942 34018 44994
rect 34638 44942 34690 44994
rect 34862 44942 34914 44994
rect 39678 44942 39730 44994
rect 43150 44942 43202 44994
rect 47406 44942 47458 44994
rect 51438 44942 51490 44994
rect 53230 44942 53282 44994
rect 55246 44942 55298 44994
rect 55918 44942 55970 44994
rect 62190 44942 62242 44994
rect 3838 44830 3890 44882
rect 16718 44830 16770 44882
rect 20302 44830 20354 44882
rect 22766 44830 22818 44882
rect 24446 44830 24498 44882
rect 33294 44830 33346 44882
rect 34302 44830 34354 44882
rect 38334 44830 38386 44882
rect 39902 44830 39954 44882
rect 44270 44830 44322 44882
rect 48862 44830 48914 44882
rect 50654 44830 50706 44882
rect 58830 44830 58882 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 2718 44494 2770 44546
rect 29262 44494 29314 44546
rect 29710 44494 29762 44546
rect 32846 44494 32898 44546
rect 36318 44494 36370 44546
rect 41358 44494 41410 44546
rect 42590 44494 42642 44546
rect 42702 44494 42754 44546
rect 43374 44494 43426 44546
rect 43934 44494 43986 44546
rect 51774 44494 51826 44546
rect 54462 44494 54514 44546
rect 59838 44494 59890 44546
rect 60622 44494 60674 44546
rect 60958 44494 61010 44546
rect 3502 44382 3554 44434
rect 4622 44382 4674 44434
rect 5742 44382 5794 44434
rect 8654 44382 8706 44434
rect 10334 44382 10386 44434
rect 12238 44382 12290 44434
rect 16718 44382 16770 44434
rect 23998 44382 24050 44434
rect 24558 44382 24610 44434
rect 26798 44382 26850 44434
rect 28030 44382 28082 44434
rect 29262 44382 29314 44434
rect 29710 44382 29762 44434
rect 30158 44382 30210 44434
rect 34414 44382 34466 44434
rect 37886 44382 37938 44434
rect 39342 44382 39394 44434
rect 40126 44382 40178 44434
rect 41022 44382 41074 44434
rect 46174 44382 46226 44434
rect 53230 44382 53282 44434
rect 1822 44270 1874 44322
rect 3390 44270 3442 44322
rect 3614 44270 3666 44322
rect 4286 44270 4338 44322
rect 4398 44270 4450 44322
rect 4734 44270 4786 44322
rect 6078 44270 6130 44322
rect 6862 44270 6914 44322
rect 7198 44270 7250 44322
rect 7646 44270 7698 44322
rect 8318 44270 8370 44322
rect 10894 44270 10946 44322
rect 12126 44270 12178 44322
rect 13806 44270 13858 44322
rect 18062 44270 18114 44322
rect 18958 44270 19010 44322
rect 20526 44270 20578 44322
rect 21758 44270 21810 44322
rect 21982 44270 22034 44322
rect 22318 44270 22370 44322
rect 23102 44270 23154 44322
rect 23662 44270 23714 44322
rect 24894 44270 24946 44322
rect 25678 44270 25730 44322
rect 34302 44270 34354 44322
rect 34974 44270 35026 44322
rect 36206 44270 36258 44322
rect 37102 44270 37154 44322
rect 37774 44270 37826 44322
rect 38670 44270 38722 44322
rect 43150 44270 43202 44322
rect 43822 44270 43874 44322
rect 44718 44270 44770 44322
rect 44942 44270 44994 44322
rect 45166 44270 45218 44322
rect 46958 44270 47010 44322
rect 47406 44270 47458 44322
rect 48302 44270 48354 44322
rect 48638 44270 48690 44322
rect 49198 44270 49250 44322
rect 50430 44270 50482 44322
rect 50990 44270 51042 44322
rect 52670 44270 52722 44322
rect 54126 44270 54178 44322
rect 55358 44270 55410 44322
rect 56142 44270 56194 44322
rect 2046 44158 2098 44210
rect 2382 44158 2434 44210
rect 2606 44158 2658 44210
rect 3054 44158 3106 44210
rect 4174 44158 4226 44210
rect 5966 44158 6018 44210
rect 11790 44158 11842 44210
rect 12350 44158 12402 44210
rect 14590 44158 14642 44210
rect 17166 44158 17218 44210
rect 18846 44158 18898 44210
rect 20638 44158 20690 44210
rect 23998 44158 24050 44210
rect 25902 44158 25954 44210
rect 26238 44158 26290 44210
rect 27694 44158 27746 44210
rect 27806 44158 27858 44210
rect 31054 44158 31106 44210
rect 37326 44158 37378 44210
rect 37438 44158 37490 44210
rect 39118 44158 39170 44210
rect 40462 44158 40514 44210
rect 41582 44158 41634 44210
rect 42142 44158 42194 44210
rect 42814 44158 42866 44210
rect 45390 44158 45442 44210
rect 49646 44158 49698 44210
rect 50654 44158 50706 44210
rect 51998 44158 52050 44210
rect 53118 44158 53170 44210
rect 56814 44158 56866 44210
rect 61182 44158 61234 44210
rect 61518 44158 61570 44210
rect 3166 44046 3218 44098
rect 12910 44046 12962 44098
rect 17054 44046 17106 44098
rect 17502 44046 17554 44098
rect 22094 44046 22146 44098
rect 22542 44046 22594 44098
rect 27918 44046 27970 44098
rect 28142 44046 28194 44098
rect 28702 44046 28754 44098
rect 38334 44046 38386 44098
rect 48750 44046 48802 44098
rect 53230 44046 53282 44098
rect 53454 44046 53506 44098
rect 58718 44046 58770 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 3950 43710 4002 43762
rect 10222 43710 10274 43762
rect 12014 43710 12066 43762
rect 14590 43710 14642 43762
rect 14814 43710 14866 43762
rect 18958 43710 19010 43762
rect 27022 43710 27074 43762
rect 29598 43710 29650 43762
rect 30382 43710 30434 43762
rect 31502 43710 31554 43762
rect 33406 43710 33458 43762
rect 37998 43710 38050 43762
rect 42254 43710 42306 43762
rect 54350 43710 54402 43762
rect 2158 43598 2210 43650
rect 4286 43598 4338 43650
rect 5182 43598 5234 43650
rect 6302 43598 6354 43650
rect 8318 43598 8370 43650
rect 8878 43598 8930 43650
rect 9662 43598 9714 43650
rect 10110 43598 10162 43650
rect 11230 43598 11282 43650
rect 11342 43598 11394 43650
rect 12910 43598 12962 43650
rect 14702 43598 14754 43650
rect 15374 43598 15426 43650
rect 15598 43598 15650 43650
rect 16158 43598 16210 43650
rect 16830 43598 16882 43650
rect 21646 43598 21698 43650
rect 23662 43598 23714 43650
rect 25454 43598 25506 43650
rect 26462 43598 26514 43650
rect 26910 43598 26962 43650
rect 27470 43598 27522 43650
rect 28254 43598 28306 43650
rect 31614 43598 31666 43650
rect 32174 43598 32226 43650
rect 33070 43598 33122 43650
rect 34078 43598 34130 43650
rect 36990 43598 37042 43650
rect 37774 43598 37826 43650
rect 37886 43598 37938 43650
rect 40910 43598 40962 43650
rect 41358 43598 41410 43650
rect 41806 43598 41858 43650
rect 43822 43598 43874 43650
rect 45278 43598 45330 43650
rect 47966 43598 48018 43650
rect 49310 43598 49362 43650
rect 54238 43598 54290 43650
rect 55582 43598 55634 43650
rect 55806 43598 55858 43650
rect 56702 43598 56754 43650
rect 57822 43598 57874 43650
rect 4174 43486 4226 43538
rect 4510 43486 4562 43538
rect 4734 43486 4786 43538
rect 5518 43486 5570 43538
rect 5966 43486 6018 43538
rect 6974 43486 7026 43538
rect 7982 43486 8034 43538
rect 8990 43486 9042 43538
rect 9550 43486 9602 43538
rect 11006 43486 11058 43538
rect 11678 43486 11730 43538
rect 12238 43486 12290 43538
rect 12462 43486 12514 43538
rect 13694 43486 13746 43538
rect 14142 43486 14194 43538
rect 15262 43486 15314 43538
rect 15934 43486 15986 43538
rect 16606 43486 16658 43538
rect 17726 43486 17778 43538
rect 18622 43486 18674 43538
rect 19518 43486 19570 43538
rect 20638 43486 20690 43538
rect 23550 43486 23602 43538
rect 24110 43486 24162 43538
rect 25342 43486 25394 43538
rect 26126 43486 26178 43538
rect 27694 43486 27746 43538
rect 28590 43486 28642 43538
rect 29374 43486 29426 43538
rect 29710 43486 29762 43538
rect 29934 43486 29986 43538
rect 30270 43486 30322 43538
rect 30606 43486 30658 43538
rect 31054 43486 31106 43538
rect 32398 43486 32450 43538
rect 34190 43486 34242 43538
rect 34862 43486 34914 43538
rect 35310 43486 35362 43538
rect 36654 43486 36706 43538
rect 37326 43486 37378 43538
rect 38110 43486 38162 43538
rect 38558 43486 38610 43538
rect 39566 43486 39618 43538
rect 40238 43486 40290 43538
rect 41134 43486 41186 43538
rect 41694 43486 41746 43538
rect 42926 43486 42978 43538
rect 44158 43486 44210 43538
rect 44270 43486 44322 43538
rect 44382 43486 44434 43538
rect 47518 43486 47570 43538
rect 48190 43486 48242 43538
rect 49758 43486 49810 43538
rect 50878 43486 50930 43538
rect 52670 43486 52722 43538
rect 52894 43486 52946 43538
rect 53902 43486 53954 43538
rect 55022 43486 55074 43538
rect 55246 43486 55298 43538
rect 55918 43486 55970 43538
rect 56478 43486 56530 43538
rect 56814 43486 56866 43538
rect 59614 43486 59666 43538
rect 7422 43374 7474 43426
rect 8094 43374 8146 43426
rect 12798 43374 12850 43426
rect 13470 43374 13522 43426
rect 17950 43374 18002 43426
rect 18398 43374 18450 43426
rect 19294 43374 19346 43426
rect 19854 43374 19906 43426
rect 20302 43374 20354 43426
rect 24558 43374 24610 43426
rect 28366 43374 28418 43426
rect 40014 43374 40066 43426
rect 42590 43374 42642 43426
rect 43934 43374 43986 43426
rect 47182 43374 47234 43426
rect 48078 43374 48130 43426
rect 48862 43374 48914 43426
rect 50094 43374 50146 43426
rect 8878 43262 8930 43314
rect 12014 43262 12066 43314
rect 23102 43262 23154 43314
rect 23662 43262 23714 43314
rect 30830 43262 30882 43314
rect 31390 43262 31442 43314
rect 39118 43262 39170 43314
rect 41470 43262 41522 43314
rect 59166 43262 59218 43314
rect 61966 43262 62018 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 2494 42926 2546 42978
rect 4174 42926 4226 42978
rect 14702 42926 14754 42978
rect 29262 42926 29314 42978
rect 30046 42926 30098 42978
rect 34750 42926 34802 42978
rect 39902 42926 39954 42978
rect 41022 42926 41074 42978
rect 44270 42926 44322 42978
rect 46062 42926 46114 42978
rect 50878 42926 50930 42978
rect 51214 42926 51266 42978
rect 52782 42926 52834 42978
rect 56366 42926 56418 42978
rect 60622 42926 60674 42978
rect 3278 42814 3330 42866
rect 4622 42814 4674 42866
rect 8654 42814 8706 42866
rect 12462 42814 12514 42866
rect 21534 42814 21586 42866
rect 22654 42814 22706 42866
rect 23886 42814 23938 42866
rect 28142 42814 28194 42866
rect 29822 42814 29874 42866
rect 31726 42814 31778 42866
rect 32510 42814 32562 42866
rect 44158 42814 44210 42866
rect 56478 42814 56530 42866
rect 1822 42702 1874 42754
rect 3726 42702 3778 42754
rect 5630 42702 5682 42754
rect 5966 42702 6018 42754
rect 6638 42702 6690 42754
rect 7086 42702 7138 42754
rect 7646 42702 7698 42754
rect 8318 42702 8370 42754
rect 10558 42702 10610 42754
rect 12798 42702 12850 42754
rect 14254 42702 14306 42754
rect 14590 42702 14642 42754
rect 14814 42702 14866 42754
rect 15150 42702 15202 42754
rect 15374 42702 15426 42754
rect 23102 42702 23154 42754
rect 24110 42702 24162 42754
rect 24894 42702 24946 42754
rect 25230 42702 25282 42754
rect 25678 42702 25730 42754
rect 29486 42702 29538 42754
rect 30494 42702 30546 42754
rect 30718 42702 30770 42754
rect 30942 42702 30994 42754
rect 31166 42702 31218 42754
rect 31502 42702 31554 42754
rect 31838 42702 31890 42754
rect 32062 42702 32114 42754
rect 33182 42702 33234 42754
rect 34302 42702 34354 42754
rect 35086 42702 35138 42754
rect 37662 42702 37714 42754
rect 38894 42702 38946 42754
rect 40238 42702 40290 42754
rect 40798 42702 40850 42754
rect 41358 42702 41410 42754
rect 41694 42702 41746 42754
rect 42814 42702 42866 42754
rect 43598 42702 43650 42754
rect 45278 42702 45330 42754
rect 45726 42702 45778 42754
rect 46734 42702 46786 42754
rect 47854 42702 47906 42754
rect 51774 42702 51826 42754
rect 52894 42702 52946 42754
rect 54574 42702 54626 42754
rect 55918 42702 55970 42754
rect 57262 42702 57314 42754
rect 58158 42702 58210 42754
rect 58942 42702 58994 42754
rect 59726 42702 59778 42754
rect 60958 42702 61010 42754
rect 61406 42702 61458 42754
rect 2158 42590 2210 42642
rect 2830 42590 2882 42642
rect 3166 42590 3218 42642
rect 3502 42590 3554 42642
rect 4062 42590 4114 42642
rect 5742 42590 5794 42642
rect 6302 42590 6354 42642
rect 10334 42590 10386 42642
rect 12350 42590 12402 42642
rect 12686 42590 12738 42642
rect 13694 42590 13746 42642
rect 16270 42590 16322 42642
rect 19070 42590 19122 42642
rect 23438 42590 23490 42642
rect 26238 42590 26290 42642
rect 27246 42590 27298 42642
rect 27358 42590 27410 42642
rect 32622 42590 32674 42642
rect 35310 42590 35362 42642
rect 35646 42590 35698 42642
rect 37774 42590 37826 42642
rect 43486 42590 43538 42642
rect 45054 42590 45106 42642
rect 51998 42590 52050 42642
rect 53230 42590 53282 42642
rect 61630 42590 61682 42642
rect 2606 42478 2658 42530
rect 5070 42478 5122 42530
rect 7198 42478 7250 42530
rect 12126 42478 12178 42530
rect 17950 42478 18002 42530
rect 20302 42478 20354 42530
rect 21982 42478 22034 42530
rect 25230 42478 25282 42530
rect 26910 42478 26962 42530
rect 27022 42478 27074 42530
rect 27134 42478 27186 42530
rect 28030 42478 28082 42530
rect 28254 42478 28306 42530
rect 28478 42478 28530 42530
rect 30158 42478 30210 42530
rect 31278 42478 31330 42530
rect 33406 42478 33458 42530
rect 33742 42478 33794 42530
rect 36542 42478 36594 42530
rect 42478 42478 42530 42530
rect 46510 42478 46562 42530
rect 49422 42478 49474 42530
rect 58606 42478 58658 42530
rect 59502 42478 59554 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 3390 42142 3442 42194
rect 5182 42142 5234 42194
rect 12014 42142 12066 42194
rect 12798 42142 12850 42194
rect 14702 42142 14754 42194
rect 15486 42142 15538 42194
rect 16606 42142 16658 42194
rect 18398 42142 18450 42194
rect 26126 42142 26178 42194
rect 35198 42142 35250 42194
rect 41918 42142 41970 42194
rect 42590 42142 42642 42194
rect 44382 42142 44434 42194
rect 45166 42142 45218 42194
rect 46398 42142 46450 42194
rect 48190 42142 48242 42194
rect 53454 42142 53506 42194
rect 54910 42142 54962 42194
rect 57822 42142 57874 42194
rect 3278 42030 3330 42082
rect 3950 42030 4002 42082
rect 6638 42030 6690 42082
rect 6750 42030 6802 42082
rect 6974 42030 7026 42082
rect 7870 42030 7922 42082
rect 7982 42030 8034 42082
rect 8094 42030 8146 42082
rect 10782 42030 10834 42082
rect 12686 42030 12738 42082
rect 13246 42030 13298 42082
rect 14926 42030 14978 42082
rect 15038 42030 15090 42082
rect 18286 42030 18338 42082
rect 19182 42030 19234 42082
rect 20526 42030 20578 42082
rect 21422 42030 21474 42082
rect 26350 42030 26402 42082
rect 26910 42030 26962 42082
rect 27806 42030 27858 42082
rect 27918 42030 27970 42082
rect 31278 42030 31330 42082
rect 33406 42030 33458 42082
rect 36766 42030 36818 42082
rect 41134 42030 41186 42082
rect 42926 42030 42978 42082
rect 49422 42030 49474 42082
rect 51998 42030 52050 42082
rect 54014 42030 54066 42082
rect 58046 42030 58098 42082
rect 2942 41918 2994 41970
rect 3614 41918 3666 41970
rect 3838 41918 3890 41970
rect 6302 41918 6354 41970
rect 7310 41918 7362 41970
rect 8318 41918 8370 41970
rect 8654 41918 8706 41970
rect 12574 41918 12626 41970
rect 13918 41918 13970 41970
rect 14142 41918 14194 41970
rect 14478 41918 14530 41970
rect 15374 41918 15426 41970
rect 15598 41918 15650 41970
rect 16158 41918 16210 41970
rect 16830 41918 16882 41970
rect 17278 41918 17330 41970
rect 17502 41918 17554 41970
rect 17614 41918 17666 41970
rect 17950 41918 18002 41970
rect 19294 41918 19346 41970
rect 20078 41918 20130 41970
rect 20750 41918 20802 41970
rect 21646 41918 21698 41970
rect 22430 41918 22482 41970
rect 22766 41918 22818 41970
rect 23214 41918 23266 41970
rect 23438 41918 23490 41970
rect 24670 41918 24722 41970
rect 25790 41918 25842 41970
rect 26014 41918 26066 41970
rect 26574 41918 26626 41970
rect 27134 41918 27186 41970
rect 28142 41918 28194 41970
rect 29038 41918 29090 41970
rect 30046 41918 30098 41970
rect 30270 41918 30322 41970
rect 30606 41918 30658 41970
rect 31054 41918 31106 41970
rect 37774 41918 37826 41970
rect 39678 41918 39730 41970
rect 40462 41918 40514 41970
rect 40910 41918 40962 41970
rect 42030 41918 42082 41970
rect 42254 41918 42306 41970
rect 42702 41918 42754 41970
rect 43262 41918 43314 41970
rect 43710 41918 43762 41970
rect 44158 41918 44210 41970
rect 45390 41918 45442 41970
rect 45838 41918 45890 41970
rect 46734 41918 46786 41970
rect 47854 41918 47906 41970
rect 53902 41918 53954 41970
rect 54798 41918 54850 41970
rect 55358 41918 55410 41970
rect 55918 41918 55970 41970
rect 57038 41918 57090 41970
rect 58158 41918 58210 41970
rect 58830 41918 58882 41970
rect 62078 41918 62130 41970
rect 2158 41806 2210 41858
rect 2606 41806 2658 41858
rect 7534 41806 7586 41858
rect 9774 41806 9826 41858
rect 14366 41806 14418 41858
rect 24334 41806 24386 41858
rect 25342 41806 25394 41858
rect 29486 41806 29538 41858
rect 30158 41806 30210 41858
rect 31838 41806 31890 41858
rect 35646 41806 35698 41858
rect 38334 41806 38386 41858
rect 39790 41806 39842 41858
rect 44494 41806 44546 41858
rect 46062 41806 46114 41858
rect 47630 41806 47682 41858
rect 50542 41806 50594 41858
rect 51102 41806 51154 41858
rect 57374 41806 57426 41858
rect 59502 41806 59554 41858
rect 61630 41806 61682 41858
rect 3950 41694 4002 41746
rect 8766 41694 8818 41746
rect 9662 41694 9714 41746
rect 15934 41694 15986 41746
rect 16494 41694 16546 41746
rect 18398 41694 18450 41746
rect 19742 41694 19794 41746
rect 22094 41694 22146 41746
rect 32174 41694 32226 41746
rect 39566 41694 39618 41746
rect 46958 41694 47010 41746
rect 47294 41694 47346 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 8654 41358 8706 41410
rect 12014 41358 12066 41410
rect 22990 41358 23042 41410
rect 34078 41358 34130 41410
rect 35534 41358 35586 41410
rect 38110 41358 38162 41410
rect 38782 41358 38834 41410
rect 39118 41358 39170 41410
rect 40798 41358 40850 41410
rect 44382 41358 44434 41410
rect 53678 41358 53730 41410
rect 54238 41358 54290 41410
rect 54462 41358 54514 41410
rect 56478 41358 56530 41410
rect 2942 41246 2994 41298
rect 5070 41246 5122 41298
rect 5742 41246 5794 41298
rect 6526 41246 6578 41298
rect 18286 41246 18338 41298
rect 20750 41246 20802 41298
rect 21758 41246 21810 41298
rect 24222 41246 24274 41298
rect 30942 41246 30994 41298
rect 32846 41246 32898 41298
rect 39342 41246 39394 41298
rect 51998 41246 52050 41298
rect 54798 41246 54850 41298
rect 60734 41246 60786 41298
rect 61070 41246 61122 41298
rect 2270 41134 2322 41186
rect 6190 41134 6242 41186
rect 7086 41134 7138 41186
rect 7534 41134 7586 41186
rect 8318 41134 8370 41186
rect 9326 41134 9378 41186
rect 9886 41134 9938 41186
rect 15262 41134 15314 41186
rect 15486 41134 15538 41186
rect 15822 41134 15874 41186
rect 15934 41134 15986 41186
rect 16046 41134 16098 41186
rect 16718 41134 16770 41186
rect 16942 41134 16994 41186
rect 19182 41134 19234 41186
rect 22094 41134 22146 41186
rect 22654 41134 22706 41186
rect 24334 41134 24386 41186
rect 28478 41134 28530 41186
rect 29374 41134 29426 41186
rect 29822 41134 29874 41186
rect 30606 41134 30658 41186
rect 31390 41134 31442 41186
rect 32174 41134 32226 41186
rect 32510 41134 32562 41186
rect 34302 41134 34354 41186
rect 34750 41134 34802 41186
rect 37886 41134 37938 41186
rect 40126 41134 40178 41186
rect 40350 41134 40402 41186
rect 41134 41134 41186 41186
rect 41470 41134 41522 41186
rect 45726 41134 45778 41186
rect 47182 41134 47234 41186
rect 48638 41134 48690 41186
rect 50094 41134 50146 41186
rect 51326 41134 51378 41186
rect 52670 41134 52722 41186
rect 52894 41134 52946 41186
rect 53790 41134 53842 41186
rect 56030 41134 56082 41186
rect 60510 41134 60562 41186
rect 61742 41134 61794 41186
rect 7758 41022 7810 41074
rect 9550 41022 9602 41074
rect 10782 41022 10834 41074
rect 12462 41022 12514 41074
rect 12910 41022 12962 41074
rect 13806 41022 13858 41074
rect 14142 41022 14194 41074
rect 14366 41022 14418 41074
rect 14926 41022 14978 41074
rect 15038 41022 15090 41074
rect 17166 41022 17218 41074
rect 19406 41022 19458 41074
rect 19742 41022 19794 41074
rect 21646 41022 21698 41074
rect 21758 41022 21810 41074
rect 21870 41022 21922 41074
rect 22990 41022 23042 41074
rect 31054 41022 31106 41074
rect 31726 41022 31778 41074
rect 32734 41022 32786 41074
rect 33406 41022 33458 41074
rect 34974 41022 35026 41074
rect 37214 41022 37266 41074
rect 40574 41022 40626 41074
rect 42590 41022 42642 41074
rect 44942 41022 44994 41074
rect 45390 41022 45442 41074
rect 49870 41022 49922 41074
rect 55358 41022 55410 41074
rect 55918 41022 55970 41074
rect 56366 41022 56418 41074
rect 56478 41022 56530 41074
rect 59726 41022 59778 41074
rect 61182 41022 61234 41074
rect 1934 40910 1986 40962
rect 9774 40910 9826 40962
rect 12350 40910 12402 40962
rect 12686 40910 12738 40962
rect 14030 40910 14082 40962
rect 16270 40910 16322 40962
rect 16942 40910 16994 40962
rect 17950 40910 18002 40962
rect 18174 40910 18226 40962
rect 18398 40910 18450 40962
rect 18846 40910 18898 40962
rect 20638 40910 20690 40962
rect 27134 40910 27186 40962
rect 32958 40910 33010 40962
rect 33742 40910 33794 40962
rect 35870 40910 35922 40962
rect 36542 40910 36594 40962
rect 36990 40910 37042 40962
rect 37102 40910 37154 40962
rect 37438 40910 37490 40962
rect 38446 40910 38498 40962
rect 40462 40910 40514 40962
rect 40910 40910 40962 40962
rect 41806 40910 41858 40962
rect 46062 40910 46114 40962
rect 50094 40910 50146 40962
rect 50766 40910 50818 40962
rect 51886 40910 51938 40962
rect 52782 40910 52834 40962
rect 53118 40910 53170 40962
rect 54574 40910 54626 40962
rect 57822 40910 57874 40962
rect 60958 40910 61010 40962
rect 61742 40910 61794 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 3726 40574 3778 40626
rect 5182 40574 5234 40626
rect 7758 40574 7810 40626
rect 10334 40574 10386 40626
rect 19518 40574 19570 40626
rect 24446 40574 24498 40626
rect 24670 40574 24722 40626
rect 25342 40574 25394 40626
rect 25902 40574 25954 40626
rect 28702 40574 28754 40626
rect 29486 40574 29538 40626
rect 42814 40574 42866 40626
rect 43038 40574 43090 40626
rect 44270 40574 44322 40626
rect 45390 40574 45442 40626
rect 55470 40574 55522 40626
rect 2718 40462 2770 40514
rect 7086 40462 7138 40514
rect 7534 40462 7586 40514
rect 15598 40462 15650 40514
rect 17726 40462 17778 40514
rect 21982 40462 22034 40514
rect 24110 40462 24162 40514
rect 24334 40462 24386 40514
rect 25678 40462 25730 40514
rect 26014 40462 26066 40514
rect 27694 40462 27746 40514
rect 30270 40462 30322 40514
rect 33630 40462 33682 40514
rect 36094 40462 36146 40514
rect 36542 40462 36594 40514
rect 37214 40462 37266 40514
rect 39230 40462 39282 40514
rect 40238 40462 40290 40514
rect 42478 40462 42530 40514
rect 42702 40462 42754 40514
rect 49310 40462 49362 40514
rect 49982 40462 50034 40514
rect 52446 40462 52498 40514
rect 54238 40462 54290 40514
rect 54574 40462 54626 40514
rect 55694 40462 55746 40514
rect 55806 40462 55858 40514
rect 57598 40462 57650 40514
rect 60622 40462 60674 40514
rect 2606 40350 2658 40402
rect 6302 40350 6354 40402
rect 6750 40350 6802 40402
rect 7422 40350 7474 40402
rect 8542 40350 8594 40402
rect 8990 40350 9042 40402
rect 11342 40350 11394 40402
rect 12126 40350 12178 40402
rect 12798 40350 12850 40402
rect 14590 40350 14642 40402
rect 15710 40350 15762 40402
rect 16830 40350 16882 40402
rect 20190 40350 20242 40402
rect 21422 40350 21474 40402
rect 22094 40350 22146 40402
rect 22542 40350 22594 40402
rect 26238 40350 26290 40402
rect 26798 40350 26850 40402
rect 28926 40350 28978 40402
rect 29150 40350 29202 40402
rect 29486 40350 29538 40402
rect 30046 40350 30098 40402
rect 30494 40350 30546 40402
rect 31278 40350 31330 40402
rect 34862 40350 34914 40402
rect 35646 40350 35698 40402
rect 40126 40350 40178 40402
rect 40462 40350 40514 40402
rect 40798 40350 40850 40402
rect 41134 40350 41186 40402
rect 41358 40350 41410 40402
rect 46846 40350 46898 40402
rect 47294 40350 47346 40402
rect 47630 40350 47682 40402
rect 49646 40350 49698 40402
rect 53230 40350 53282 40402
rect 55134 40350 55186 40402
rect 57822 40350 57874 40402
rect 58606 40350 58658 40402
rect 58942 40350 58994 40402
rect 60510 40350 60562 40402
rect 61406 40350 61458 40402
rect 62078 40350 62130 40402
rect 2270 40238 2322 40290
rect 3390 40238 3442 40290
rect 9886 40238 9938 40290
rect 11454 40238 11506 40290
rect 14702 40238 14754 40290
rect 16270 40238 16322 40290
rect 23886 40238 23938 40290
rect 27358 40238 27410 40290
rect 27918 40238 27970 40290
rect 29038 40238 29090 40290
rect 31166 40238 31218 40290
rect 32622 40238 32674 40290
rect 35422 40238 35474 40290
rect 41022 40238 41074 40290
rect 41918 40238 41970 40290
rect 42702 40238 42754 40290
rect 46062 40238 46114 40290
rect 50318 40238 50370 40290
rect 61182 40238 61234 40290
rect 11006 40126 11058 40178
rect 14590 40126 14642 40178
rect 15598 40126 15650 40178
rect 16494 40126 16546 40178
rect 28254 40126 28306 40178
rect 29822 40126 29874 40178
rect 31614 40126 31666 40178
rect 48750 40126 48802 40178
rect 49086 40126 49138 40178
rect 54798 40126 54850 40178
rect 57262 40126 57314 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 8318 39790 8370 39842
rect 12350 39790 12402 39842
rect 16830 39790 16882 39842
rect 21422 39790 21474 39842
rect 28478 39790 28530 39842
rect 30942 39790 30994 39842
rect 44942 39790 44994 39842
rect 49310 39790 49362 39842
rect 52110 39790 52162 39842
rect 62078 39790 62130 39842
rect 4174 39678 4226 39730
rect 6078 39678 6130 39730
rect 7758 39678 7810 39730
rect 12462 39678 12514 39730
rect 13694 39678 13746 39730
rect 14814 39678 14866 39730
rect 24558 39678 24610 39730
rect 26126 39678 26178 39730
rect 28142 39678 28194 39730
rect 31166 39678 31218 39730
rect 32958 39678 33010 39730
rect 40014 39678 40066 39730
rect 41582 39678 41634 39730
rect 43934 39678 43986 39730
rect 44270 39678 44322 39730
rect 53230 39678 53282 39730
rect 53566 39678 53618 39730
rect 53790 39678 53842 39730
rect 57934 39678 57986 39730
rect 59502 39678 59554 39730
rect 61070 39678 61122 39730
rect 4398 39566 4450 39618
rect 6414 39566 6466 39618
rect 6862 39566 6914 39618
rect 7870 39566 7922 39618
rect 8878 39566 8930 39618
rect 9662 39566 9714 39618
rect 9998 39566 10050 39618
rect 10334 39566 10386 39618
rect 11006 39566 11058 39618
rect 11454 39566 11506 39618
rect 14030 39566 14082 39618
rect 15262 39566 15314 39618
rect 18398 39566 18450 39618
rect 19294 39566 19346 39618
rect 20414 39566 20466 39618
rect 21310 39566 21362 39618
rect 23102 39566 23154 39618
rect 23550 39566 23602 39618
rect 24110 39566 24162 39618
rect 26350 39566 26402 39618
rect 27470 39566 27522 39618
rect 28254 39566 28306 39618
rect 29598 39566 29650 39618
rect 31054 39566 31106 39618
rect 31502 39566 31554 39618
rect 32846 39566 32898 39618
rect 33518 39566 33570 39618
rect 33854 39566 33906 39618
rect 35086 39566 35138 39618
rect 37214 39566 37266 39618
rect 40798 39566 40850 39618
rect 41918 39566 41970 39618
rect 42926 39566 42978 39618
rect 47518 39566 47570 39618
rect 47966 39566 48018 39618
rect 49422 39566 49474 39618
rect 49982 39566 50034 39618
rect 50430 39566 50482 39618
rect 51998 39566 52050 39618
rect 56142 39566 56194 39618
rect 58270 39566 58322 39618
rect 59054 39566 59106 39618
rect 59278 39566 59330 39618
rect 59614 39566 59666 39618
rect 59838 39566 59890 39618
rect 60510 39566 60562 39618
rect 61518 39566 61570 39618
rect 2382 39454 2434 39506
rect 6302 39454 6354 39506
rect 7310 39454 7362 39506
rect 8654 39454 8706 39506
rect 12798 39454 12850 39506
rect 14142 39454 14194 39506
rect 14814 39454 14866 39506
rect 16046 39454 16098 39506
rect 16606 39454 16658 39506
rect 17614 39454 17666 39506
rect 17950 39454 18002 39506
rect 22318 39454 22370 39506
rect 22654 39454 22706 39506
rect 27358 39454 27410 39506
rect 29934 39454 29986 39506
rect 30382 39454 30434 39506
rect 33966 39454 34018 39506
rect 35982 39454 36034 39506
rect 37886 39454 37938 39506
rect 41134 39454 41186 39506
rect 41470 39454 41522 39506
rect 42702 39454 42754 39506
rect 46286 39454 46338 39506
rect 47294 39454 47346 39506
rect 48862 39454 48914 39506
rect 54686 39454 54738 39506
rect 54798 39454 54850 39506
rect 56366 39454 56418 39506
rect 60622 39454 60674 39506
rect 62190 39454 62242 39506
rect 3726 39342 3778 39394
rect 4734 39342 4786 39394
rect 9774 39342 9826 39394
rect 10782 39342 10834 39394
rect 17166 39342 17218 39394
rect 18510 39342 18562 39394
rect 22878 39342 22930 39394
rect 29262 39342 29314 39394
rect 32510 39342 32562 39394
rect 33070 39342 33122 39394
rect 40462 39342 40514 39394
rect 43598 39342 43650 39394
rect 47406 39342 47458 39394
rect 52670 39342 52722 39394
rect 54910 39342 54962 39394
rect 55022 39342 55074 39394
rect 55134 39342 55186 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 3838 39006 3890 39058
rect 8878 39006 8930 39058
rect 10110 39006 10162 39058
rect 12014 39006 12066 39058
rect 16830 39006 16882 39058
rect 17502 39006 17554 39058
rect 18510 39006 18562 39058
rect 20414 39006 20466 39058
rect 24558 39006 24610 39058
rect 25566 39006 25618 39058
rect 26126 39006 26178 39058
rect 27246 39006 27298 39058
rect 38670 39006 38722 39058
rect 41134 39006 41186 39058
rect 46510 39006 46562 39058
rect 47854 39006 47906 39058
rect 47966 39006 48018 39058
rect 2158 38894 2210 38946
rect 4734 38894 4786 38946
rect 5070 38894 5122 38946
rect 6974 38894 7026 38946
rect 7310 38894 7362 38946
rect 11118 38894 11170 38946
rect 13022 38894 13074 38946
rect 16270 38894 16322 38946
rect 17614 38894 17666 38946
rect 17726 38894 17778 38946
rect 17838 38894 17890 38946
rect 21534 38894 21586 38946
rect 23550 38894 23602 38946
rect 23998 38894 24050 38946
rect 30382 38894 30434 38946
rect 30718 38894 30770 38946
rect 36878 38894 36930 38946
rect 40238 38894 40290 38946
rect 40350 38894 40402 38946
rect 41358 38894 41410 38946
rect 45502 38894 45554 38946
rect 47518 38894 47570 38946
rect 47630 38894 47682 38946
rect 47742 38894 47794 38946
rect 48750 38894 48802 38946
rect 51774 38894 51826 38946
rect 52670 38894 52722 38946
rect 53006 38894 53058 38946
rect 53454 38894 53506 38946
rect 54798 38894 54850 38946
rect 60510 38894 60562 38946
rect 4062 38782 4114 38834
rect 4510 38782 4562 38834
rect 5406 38782 5458 38834
rect 5630 38782 5682 38834
rect 5966 38782 6018 38834
rect 7534 38782 7586 38834
rect 8542 38782 8594 38834
rect 9550 38782 9602 38834
rect 9998 38782 10050 38834
rect 10222 38782 10274 38834
rect 11230 38782 11282 38834
rect 13358 38782 13410 38834
rect 14366 38782 14418 38834
rect 16494 38782 16546 38834
rect 17390 38782 17442 38834
rect 18734 38782 18786 38834
rect 19182 38782 19234 38834
rect 19406 38782 19458 38834
rect 19854 38782 19906 38834
rect 24222 38782 24274 38834
rect 28590 38782 28642 38834
rect 29038 38782 29090 38834
rect 29262 38782 29314 38834
rect 31054 38782 31106 38834
rect 32174 38782 32226 38834
rect 32510 38782 32562 38834
rect 32958 38782 33010 38834
rect 33406 38782 33458 38834
rect 33518 38782 33570 38834
rect 35534 38782 35586 38834
rect 35982 38782 36034 38834
rect 36430 38782 36482 38834
rect 42142 38782 42194 38834
rect 45838 38782 45890 38834
rect 46062 38782 46114 38834
rect 46734 38782 46786 38834
rect 49086 38782 49138 38834
rect 49870 38782 49922 38834
rect 51998 38782 52050 38834
rect 52446 38782 52498 38834
rect 53342 38782 53394 38834
rect 55918 38782 55970 38834
rect 56814 38782 56866 38834
rect 57710 38782 57762 38834
rect 59614 38782 59666 38834
rect 59726 38782 59778 38834
rect 60734 38782 60786 38834
rect 61406 38782 61458 38834
rect 4286 38670 4338 38722
rect 6302 38670 6354 38722
rect 8318 38670 8370 38722
rect 11678 38670 11730 38722
rect 14702 38670 14754 38722
rect 18622 38670 18674 38722
rect 22542 38670 22594 38722
rect 22654 38670 22706 38722
rect 25678 38670 25730 38722
rect 31278 38670 31330 38722
rect 33182 38670 33234 38722
rect 41246 38670 41298 38722
rect 41582 38670 41634 38722
rect 42926 38670 42978 38722
rect 45054 38670 45106 38722
rect 46622 38670 46674 38722
rect 49198 38670 49250 38722
rect 50318 38670 50370 38722
rect 50878 38670 50930 38722
rect 52894 38670 52946 38722
rect 57262 38670 57314 38722
rect 61854 38670 61906 38722
rect 7870 38558 7922 38610
rect 12686 38558 12738 38610
rect 28702 38558 28754 38610
rect 37438 38558 37490 38610
rect 39790 38558 39842 38610
rect 41806 38558 41858 38610
rect 51214 38558 51266 38610
rect 53454 38558 53506 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 13582 38222 13634 38274
rect 17278 38222 17330 38274
rect 25230 38222 25282 38274
rect 34190 38222 34242 38274
rect 42702 38222 42754 38274
rect 55806 38222 55858 38274
rect 58494 38222 58546 38274
rect 2046 38110 2098 38162
rect 2382 38110 2434 38162
rect 3614 38110 3666 38162
rect 4958 38110 5010 38162
rect 11678 38110 11730 38162
rect 12686 38110 12738 38162
rect 20302 38110 20354 38162
rect 22990 38110 23042 38162
rect 28142 38110 28194 38162
rect 32062 38110 32114 38162
rect 34414 38110 34466 38162
rect 43934 38110 43986 38162
rect 44942 38110 44994 38162
rect 46398 38110 46450 38162
rect 3726 37998 3778 38050
rect 4734 37998 4786 38050
rect 8094 37998 8146 38050
rect 8318 37998 8370 38050
rect 8654 37998 8706 38050
rect 8990 37998 9042 38050
rect 9550 37998 9602 38050
rect 10446 37998 10498 38050
rect 11006 37998 11058 38050
rect 13694 37998 13746 38050
rect 15150 37998 15202 38050
rect 15598 37998 15650 38050
rect 19854 37998 19906 38050
rect 20414 37998 20466 38050
rect 21198 37998 21250 38050
rect 21534 37998 21586 38050
rect 22430 37998 22482 38050
rect 23326 37998 23378 38050
rect 24110 37998 24162 38050
rect 25566 37998 25618 38050
rect 25790 37998 25842 38050
rect 28478 37998 28530 38050
rect 29822 37998 29874 38050
rect 30158 37998 30210 38050
rect 31950 37998 32002 38050
rect 34078 37998 34130 38050
rect 34862 37998 34914 38050
rect 35086 37998 35138 38050
rect 36094 37998 36146 38050
rect 37998 37998 38050 38050
rect 41694 37998 41746 38050
rect 42702 37998 42754 38050
rect 43822 37998 43874 38050
rect 45278 37998 45330 38050
rect 46062 37998 46114 38050
rect 46622 37998 46674 38050
rect 47182 37998 47234 38050
rect 48414 37998 48466 38050
rect 48974 37998 49026 38050
rect 50766 37998 50818 38050
rect 52110 37998 52162 38050
rect 52670 37998 52722 38050
rect 53230 37998 53282 38050
rect 53790 37998 53842 38050
rect 54798 37998 54850 38050
rect 55918 37998 55970 38050
rect 57822 37998 57874 38050
rect 58830 37998 58882 38050
rect 59502 37998 59554 38050
rect 60510 37998 60562 38050
rect 61294 37998 61346 38050
rect 61966 37998 62018 38050
rect 2606 37886 2658 37938
rect 2718 37886 2770 37938
rect 3390 37886 3442 37938
rect 6078 37886 6130 37938
rect 9102 37886 9154 37938
rect 14366 37886 14418 37938
rect 18510 37886 18562 37938
rect 19518 37886 19570 37938
rect 21422 37886 21474 37938
rect 21870 37886 21922 37938
rect 22878 37886 22930 37938
rect 24558 37886 24610 37938
rect 29150 37886 29202 37938
rect 29486 37886 29538 37938
rect 32958 37886 33010 37938
rect 37214 37886 37266 37938
rect 38222 37886 38274 37938
rect 38670 37886 38722 37938
rect 40014 37886 40066 37938
rect 43038 37886 43090 37938
rect 43262 37886 43314 37938
rect 44158 37886 44210 37938
rect 45726 37886 45778 37938
rect 45838 37886 45890 37938
rect 46286 37886 46338 37938
rect 46846 37886 46898 37938
rect 47294 37886 47346 37938
rect 47854 37886 47906 37938
rect 48078 37886 48130 37938
rect 48190 37886 48242 37938
rect 49310 37886 49362 37938
rect 50318 37886 50370 37938
rect 53454 37886 53506 37938
rect 53902 37886 53954 37938
rect 57150 37886 57202 37938
rect 59614 37886 59666 37938
rect 60846 37886 60898 37938
rect 2270 37774 2322 37826
rect 2494 37774 2546 37826
rect 7758 37774 7810 37826
rect 9326 37774 9378 37826
rect 12238 37774 12290 37826
rect 20190 37774 20242 37826
rect 20638 37774 20690 37826
rect 27806 37774 27858 37826
rect 35870 37774 35922 37826
rect 36878 37774 36930 37826
rect 37102 37774 37154 37826
rect 37662 37774 37714 37826
rect 43150 37774 43202 37826
rect 48302 37774 48354 37826
rect 60622 37774 60674 37826
rect 60734 37774 60786 37826
rect 61630 37774 61682 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 2046 37438 2098 37490
rect 3054 37438 3106 37490
rect 6414 37438 6466 37490
rect 8318 37438 8370 37490
rect 8654 37438 8706 37490
rect 15710 37438 15762 37490
rect 15822 37438 15874 37490
rect 15934 37438 15986 37490
rect 25342 37438 25394 37490
rect 32510 37438 32562 37490
rect 40910 37438 40962 37490
rect 41134 37438 41186 37490
rect 43486 37438 43538 37490
rect 47966 37438 48018 37490
rect 48862 37438 48914 37490
rect 51214 37438 51266 37490
rect 52670 37438 52722 37490
rect 54014 37438 54066 37490
rect 61854 37438 61906 37490
rect 2494 37326 2546 37378
rect 2718 37326 2770 37378
rect 2830 37326 2882 37378
rect 7422 37326 7474 37378
rect 8878 37326 8930 37378
rect 8990 37326 9042 37378
rect 10222 37326 10274 37378
rect 14478 37326 14530 37378
rect 16046 37326 16098 37378
rect 16158 37326 16210 37378
rect 18622 37326 18674 37378
rect 21646 37326 21698 37378
rect 25678 37326 25730 37378
rect 26574 37326 26626 37378
rect 37438 37326 37490 37378
rect 39678 37326 39730 37378
rect 41358 37326 41410 37378
rect 41918 37326 41970 37378
rect 42142 37326 42194 37378
rect 43374 37326 43426 37378
rect 45838 37326 45890 37378
rect 46398 37326 46450 37378
rect 46734 37326 46786 37378
rect 49422 37326 49474 37378
rect 50318 37326 50370 37378
rect 55806 37326 55858 37378
rect 56590 37326 56642 37378
rect 56702 37326 56754 37378
rect 60062 37326 60114 37378
rect 3614 37214 3666 37266
rect 5294 37214 5346 37266
rect 6638 37214 6690 37266
rect 7198 37214 7250 37266
rect 12014 37214 12066 37266
rect 12574 37214 12626 37266
rect 14254 37214 14306 37266
rect 14702 37214 14754 37266
rect 17502 37214 17554 37266
rect 17950 37214 18002 37266
rect 25902 37214 25954 37266
rect 27022 37214 27074 37266
rect 27694 37214 27746 37266
rect 28590 37214 28642 37266
rect 29374 37214 29426 37266
rect 31166 37214 31218 37266
rect 31502 37214 31554 37266
rect 33406 37214 33458 37266
rect 33630 37214 33682 37266
rect 36430 37214 36482 37266
rect 37998 37214 38050 37266
rect 39342 37214 39394 37266
rect 40350 37214 40402 37266
rect 41022 37214 41074 37266
rect 43150 37214 43202 37266
rect 43598 37214 43650 37266
rect 43710 37214 43762 37266
rect 44270 37214 44322 37266
rect 46622 37214 46674 37266
rect 47518 37214 47570 37266
rect 47742 37214 47794 37266
rect 48190 37214 48242 37266
rect 48750 37214 48802 37266
rect 49310 37214 49362 37266
rect 50206 37214 50258 37266
rect 51102 37214 51154 37266
rect 51550 37214 51602 37266
rect 51886 37214 51938 37266
rect 52222 37214 52274 37266
rect 52558 37214 52610 37266
rect 53566 37214 53618 37266
rect 54238 37214 54290 37266
rect 54910 37214 54962 37266
rect 56030 37214 56082 37266
rect 56926 37214 56978 37266
rect 58494 37214 58546 37266
rect 60398 37214 60450 37266
rect 61070 37214 61122 37266
rect 62078 37214 62130 37266
rect 2718 37102 2770 37154
rect 3502 37102 3554 37154
rect 5742 37102 5794 37154
rect 20750 37102 20802 37154
rect 24670 37102 24722 37154
rect 26238 37102 26290 37154
rect 27918 37102 27970 37154
rect 28926 37102 28978 37154
rect 33854 37102 33906 37154
rect 36206 37102 36258 37154
rect 38782 37102 38834 37154
rect 39790 37102 39842 37154
rect 44382 37102 44434 37154
rect 47182 37102 47234 37154
rect 48078 37102 48130 37154
rect 51774 37102 51826 37154
rect 54126 37102 54178 37154
rect 55358 37102 55410 37154
rect 58382 37102 58434 37154
rect 61518 37102 61570 37154
rect 7982 36990 8034 37042
rect 11342 36990 11394 37042
rect 23662 36990 23714 37042
rect 26686 36990 26738 37042
rect 26910 36990 26962 37042
rect 33182 36990 33234 37042
rect 35982 36990 36034 37042
rect 42030 36990 42082 37042
rect 42478 36990 42530 37042
rect 42702 36990 42754 37042
rect 57710 36990 57762 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 4174 36654 4226 36706
rect 6526 36654 6578 36706
rect 12798 36654 12850 36706
rect 24670 36654 24722 36706
rect 48750 36654 48802 36706
rect 57374 36654 57426 36706
rect 2494 36542 2546 36594
rect 3950 36542 4002 36594
rect 5070 36542 5122 36594
rect 8990 36542 9042 36594
rect 13918 36542 13970 36594
rect 17502 36542 17554 36594
rect 18286 36542 18338 36594
rect 20526 36542 20578 36594
rect 23326 36542 23378 36594
rect 27918 36542 27970 36594
rect 32174 36542 32226 36594
rect 37886 36542 37938 36594
rect 46174 36542 46226 36594
rect 46846 36542 46898 36594
rect 56030 36542 56082 36594
rect 60622 36542 60674 36594
rect 3278 36430 3330 36482
rect 4398 36430 4450 36482
rect 11006 36430 11058 36482
rect 11230 36430 11282 36482
rect 11790 36430 11842 36482
rect 16830 36430 16882 36482
rect 17614 36430 17666 36482
rect 18398 36430 18450 36482
rect 19294 36430 19346 36482
rect 19742 36430 19794 36482
rect 20750 36430 20802 36482
rect 21646 36430 21698 36482
rect 22318 36430 22370 36482
rect 23998 36430 24050 36482
rect 25454 36430 25506 36482
rect 25678 36430 25730 36482
rect 28030 36430 28082 36482
rect 28254 36430 28306 36482
rect 28366 36430 28418 36482
rect 29374 36430 29426 36482
rect 30382 36430 30434 36482
rect 31614 36430 31666 36482
rect 31950 36430 32002 36482
rect 35086 36430 35138 36482
rect 35870 36430 35922 36482
rect 37438 36430 37490 36482
rect 37774 36430 37826 36482
rect 39902 36430 39954 36482
rect 41470 36430 41522 36482
rect 42030 36430 42082 36482
rect 44830 36430 44882 36482
rect 45054 36430 45106 36482
rect 46398 36430 46450 36482
rect 47182 36430 47234 36482
rect 47854 36430 47906 36482
rect 48190 36430 48242 36482
rect 48750 36430 48802 36482
rect 50206 36430 50258 36482
rect 50430 36430 50482 36482
rect 52782 36430 52834 36482
rect 52894 36430 52946 36482
rect 53118 36430 53170 36482
rect 54014 36430 54066 36482
rect 54462 36430 54514 36482
rect 55806 36430 55858 36482
rect 56702 36430 56754 36482
rect 61294 36430 61346 36482
rect 61630 36430 61682 36482
rect 61966 36430 62018 36482
rect 2158 36318 2210 36370
rect 2942 36318 2994 36370
rect 5630 36318 5682 36370
rect 9214 36318 9266 36370
rect 12014 36318 12066 36370
rect 16046 36318 16098 36370
rect 17950 36318 18002 36370
rect 22542 36318 22594 36370
rect 24334 36318 24386 36370
rect 27806 36318 27858 36370
rect 29150 36318 29202 36370
rect 32958 36318 33010 36370
rect 34526 36318 34578 36370
rect 34862 36318 34914 36370
rect 36430 36318 36482 36370
rect 39678 36318 39730 36370
rect 40910 36318 40962 36370
rect 43934 36318 43986 36370
rect 46286 36318 46338 36370
rect 48078 36318 48130 36370
rect 49086 36318 49138 36370
rect 53230 36318 53282 36370
rect 54798 36318 54850 36370
rect 56030 36318 56082 36370
rect 56478 36318 56530 36370
rect 59278 36318 59330 36370
rect 60958 36318 61010 36370
rect 61518 36318 61570 36370
rect 2382 36206 2434 36258
rect 2606 36206 2658 36258
rect 5966 36206 6018 36258
rect 7870 36206 7922 36258
rect 13582 36206 13634 36258
rect 21534 36206 21586 36258
rect 21982 36206 22034 36258
rect 22878 36206 22930 36258
rect 35422 36206 35474 36258
rect 45390 36206 45442 36258
rect 53678 36206 53730 36258
rect 60510 36206 60562 36258
rect 60734 36206 60786 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 2046 35870 2098 35922
rect 8878 35870 8930 35922
rect 11006 35870 11058 35922
rect 11454 35870 11506 35922
rect 13022 35870 13074 35922
rect 13134 35870 13186 35922
rect 17502 35870 17554 35922
rect 18286 35870 18338 35922
rect 18398 35870 18450 35922
rect 22430 35870 22482 35922
rect 29150 35870 29202 35922
rect 30606 35870 30658 35922
rect 32510 35870 32562 35922
rect 35198 35870 35250 35922
rect 35422 35870 35474 35922
rect 40126 35870 40178 35922
rect 40238 35870 40290 35922
rect 42926 35870 42978 35922
rect 56702 35870 56754 35922
rect 58382 35870 58434 35922
rect 62190 35870 62242 35922
rect 2382 35758 2434 35810
rect 3390 35758 3442 35810
rect 7310 35758 7362 35810
rect 7982 35758 8034 35810
rect 10110 35758 10162 35810
rect 12574 35758 12626 35810
rect 12798 35758 12850 35810
rect 12910 35758 12962 35810
rect 14142 35758 14194 35810
rect 21086 35758 21138 35810
rect 22990 35758 23042 35810
rect 26014 35758 26066 35810
rect 33854 35758 33906 35810
rect 34190 35758 34242 35810
rect 35086 35758 35138 35810
rect 39790 35758 39842 35810
rect 40014 35758 40066 35810
rect 40350 35758 40402 35810
rect 41134 35758 41186 35810
rect 43710 35758 43762 35810
rect 44270 35758 44322 35810
rect 45054 35758 45106 35810
rect 46846 35758 46898 35810
rect 47630 35758 47682 35810
rect 48750 35758 48802 35810
rect 48862 35758 48914 35810
rect 53342 35758 53394 35810
rect 57374 35758 57426 35810
rect 59614 35758 59666 35810
rect 1934 35646 1986 35698
rect 2158 35646 2210 35698
rect 3502 35646 3554 35698
rect 4734 35646 4786 35698
rect 5966 35646 6018 35698
rect 7086 35646 7138 35698
rect 7758 35646 7810 35698
rect 8542 35646 8594 35698
rect 9774 35646 9826 35698
rect 10670 35646 10722 35698
rect 11342 35646 11394 35698
rect 11566 35646 11618 35698
rect 12014 35646 12066 35698
rect 14590 35646 14642 35698
rect 15150 35646 15202 35698
rect 15374 35646 15426 35698
rect 17390 35646 17442 35698
rect 17614 35646 17666 35698
rect 18062 35646 18114 35698
rect 18510 35646 18562 35698
rect 18846 35646 18898 35698
rect 19630 35646 19682 35698
rect 23214 35646 23266 35698
rect 24110 35646 24162 35698
rect 25230 35646 25282 35698
rect 33182 35646 33234 35698
rect 33518 35646 33570 35698
rect 34414 35646 34466 35698
rect 36318 35646 36370 35698
rect 36654 35646 36706 35698
rect 38558 35646 38610 35698
rect 38782 35646 38834 35698
rect 40910 35646 40962 35698
rect 42030 35646 42082 35698
rect 42366 35646 42418 35698
rect 42814 35646 42866 35698
rect 43486 35646 43538 35698
rect 44494 35646 44546 35698
rect 45390 35646 45442 35698
rect 47182 35646 47234 35698
rect 47854 35646 47906 35698
rect 48190 35646 48242 35698
rect 49310 35646 49362 35698
rect 50094 35646 50146 35698
rect 51886 35646 51938 35698
rect 51998 35646 52050 35698
rect 52222 35646 52274 35698
rect 53230 35646 53282 35698
rect 54462 35646 54514 35698
rect 57262 35646 57314 35698
rect 58830 35646 58882 35698
rect 4286 35534 4338 35586
rect 10446 35534 10498 35586
rect 19966 35534 20018 35586
rect 24446 35534 24498 35586
rect 28142 35534 28194 35586
rect 31950 35534 32002 35586
rect 36542 35534 36594 35586
rect 41470 35534 41522 35586
rect 47742 35534 47794 35586
rect 53566 35534 53618 35586
rect 54014 35534 54066 35586
rect 55470 35534 55522 35586
rect 61742 35534 61794 35586
rect 14366 35422 14418 35474
rect 23550 35422 23602 35474
rect 48862 35422 48914 35474
rect 55694 35422 55746 35474
rect 56030 35422 56082 35474
rect 58046 35422 58098 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 3054 35086 3106 35138
rect 5854 35086 5906 35138
rect 13582 35086 13634 35138
rect 13918 35086 13970 35138
rect 23326 35086 23378 35138
rect 40574 35086 40626 35138
rect 44830 35086 44882 35138
rect 44942 35086 44994 35138
rect 45166 35086 45218 35138
rect 45278 35086 45330 35138
rect 49086 35086 49138 35138
rect 50094 35086 50146 35138
rect 53006 35086 53058 35138
rect 53566 35086 53618 35138
rect 53790 35086 53842 35138
rect 55470 35086 55522 35138
rect 55582 35086 55634 35138
rect 61070 35086 61122 35138
rect 61742 35086 61794 35138
rect 4062 34974 4114 35026
rect 22542 34974 22594 35026
rect 28478 34974 28530 35026
rect 31390 34974 31442 35026
rect 34414 34974 34466 35026
rect 37102 34974 37154 35026
rect 43710 34974 43762 35026
rect 51774 34974 51826 35026
rect 2606 34862 2658 34914
rect 4174 34862 4226 34914
rect 4510 34862 4562 34914
rect 6190 34862 6242 34914
rect 6862 34862 6914 34914
rect 7534 34862 7586 34914
rect 7870 34862 7922 34914
rect 7982 34862 8034 34914
rect 8094 34862 8146 34914
rect 8654 34862 8706 34914
rect 9102 34862 9154 34914
rect 9326 34862 9378 34914
rect 9662 34862 9714 34914
rect 9998 34862 10050 34914
rect 11118 34862 11170 34914
rect 11790 34862 11842 34914
rect 14590 34862 14642 34914
rect 15262 34862 15314 34914
rect 15598 34862 15650 34914
rect 15822 34862 15874 34914
rect 16046 34862 16098 34914
rect 17390 34862 17442 34914
rect 21534 34862 21586 34914
rect 22206 34862 22258 34914
rect 23102 34862 23154 34914
rect 23662 34862 23714 34914
rect 23998 34862 24050 34914
rect 25118 34862 25170 34914
rect 25678 34862 25730 34914
rect 27134 34862 27186 34914
rect 28142 34862 28194 34914
rect 28366 34862 28418 34914
rect 28590 34862 28642 34914
rect 30158 34862 30210 34914
rect 31838 34862 31890 34914
rect 33070 34862 33122 34914
rect 33966 34862 34018 34914
rect 35086 34862 35138 34914
rect 37550 34862 37602 34914
rect 38110 34862 38162 34914
rect 39566 34862 39618 34914
rect 41022 34862 41074 34914
rect 42254 34862 42306 34914
rect 42814 34862 42866 34914
rect 43598 34862 43650 34914
rect 46286 34862 46338 34914
rect 47742 34862 47794 34914
rect 48190 34862 48242 34914
rect 49198 34862 49250 34914
rect 50430 34862 50482 34914
rect 51214 34862 51266 34914
rect 51662 34862 51714 34914
rect 54238 34862 54290 34914
rect 55806 34862 55858 34914
rect 56926 34862 56978 34914
rect 58046 34862 58098 34914
rect 58270 34862 58322 34914
rect 59838 34862 59890 34914
rect 60734 34862 60786 34914
rect 2382 34750 2434 34802
rect 6750 34750 6802 34802
rect 12798 34750 12850 34802
rect 14478 34750 14530 34802
rect 15374 34750 15426 34802
rect 18286 34750 18338 34802
rect 20750 34750 20802 34802
rect 21422 34750 21474 34802
rect 24894 34750 24946 34802
rect 27582 34750 27634 34802
rect 29150 34750 29202 34802
rect 30270 34750 30322 34802
rect 35534 34750 35586 34802
rect 35870 34750 35922 34802
rect 40574 34750 40626 34802
rect 42926 34750 42978 34802
rect 50990 34750 51042 34802
rect 53230 34750 53282 34802
rect 53342 34750 53394 34802
rect 54574 34750 54626 34802
rect 54686 34750 54738 34802
rect 55918 34750 55970 34802
rect 56590 34750 56642 34802
rect 57150 34750 57202 34802
rect 59614 34750 59666 34802
rect 60510 34750 60562 34802
rect 61966 34750 62018 34802
rect 1934 34638 1986 34690
rect 3390 34638 3442 34690
rect 4734 34638 4786 34690
rect 8318 34638 8370 34690
rect 8766 34638 8818 34690
rect 10110 34638 10162 34690
rect 12686 34638 12738 34690
rect 16382 34638 16434 34690
rect 16718 34638 16770 34690
rect 16830 34638 16882 34690
rect 16942 34638 16994 34690
rect 20078 34638 20130 34690
rect 20414 34638 20466 34690
rect 29262 34638 29314 34690
rect 29374 34638 29426 34690
rect 35086 34638 35138 34690
rect 37774 34638 37826 34690
rect 41918 34638 41970 34690
rect 45838 34638 45890 34690
rect 54350 34638 54402 34690
rect 54462 34638 54514 34690
rect 56254 34638 56306 34690
rect 61406 34638 61458 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 2494 34302 2546 34354
rect 11790 34302 11842 34354
rect 12910 34302 12962 34354
rect 15486 34302 15538 34354
rect 17278 34302 17330 34354
rect 22654 34302 22706 34354
rect 24670 34302 24722 34354
rect 27358 34302 27410 34354
rect 32398 34302 32450 34354
rect 36206 34302 36258 34354
rect 40350 34302 40402 34354
rect 41470 34302 41522 34354
rect 41694 34302 41746 34354
rect 42702 34302 42754 34354
rect 43598 34302 43650 34354
rect 46846 34302 46898 34354
rect 47742 34302 47794 34354
rect 55246 34302 55298 34354
rect 59166 34302 59218 34354
rect 3390 34190 3442 34242
rect 10782 34190 10834 34242
rect 12126 34190 12178 34242
rect 13470 34190 13522 34242
rect 14030 34190 14082 34242
rect 15038 34190 15090 34242
rect 15374 34190 15426 34242
rect 17502 34190 17554 34242
rect 18174 34190 18226 34242
rect 18398 34190 18450 34242
rect 18510 34190 18562 34242
rect 19854 34190 19906 34242
rect 28254 34190 28306 34242
rect 29822 34190 29874 34242
rect 30382 34190 30434 34242
rect 32174 34190 32226 34242
rect 32286 34190 32338 34242
rect 33406 34190 33458 34242
rect 35982 34190 36034 34242
rect 36094 34190 36146 34242
rect 36654 34190 36706 34242
rect 38894 34190 38946 34242
rect 41022 34190 41074 34242
rect 42590 34190 42642 34242
rect 43150 34190 43202 34242
rect 45390 34190 45442 34242
rect 48750 34190 48802 34242
rect 49086 34190 49138 34242
rect 52110 34190 52162 34242
rect 55918 34190 55970 34242
rect 57038 34190 57090 34242
rect 60734 34190 60786 34242
rect 61742 34190 61794 34242
rect 2158 34078 2210 34130
rect 2382 34078 2434 34130
rect 2718 34078 2770 34130
rect 3166 34078 3218 34130
rect 4734 34078 4786 34130
rect 6078 34078 6130 34130
rect 6862 34078 6914 34130
rect 7646 34078 7698 34130
rect 15822 34078 15874 34130
rect 16270 34078 16322 34130
rect 17614 34078 17666 34130
rect 18734 34078 18786 34130
rect 22990 34078 23042 34130
rect 23438 34078 23490 34130
rect 26126 34078 26178 34130
rect 27694 34078 27746 34130
rect 29598 34078 29650 34130
rect 31054 34078 31106 34130
rect 31726 34078 31778 34130
rect 32510 34078 32562 34130
rect 35646 34078 35698 34130
rect 36318 34078 36370 34130
rect 36878 34078 36930 34130
rect 37774 34078 37826 34130
rect 39006 34078 39058 34130
rect 39678 34078 39730 34130
rect 39902 34078 39954 34130
rect 40798 34078 40850 34130
rect 41134 34078 41186 34130
rect 41918 34078 41970 34130
rect 42142 34078 42194 34130
rect 42814 34078 42866 34130
rect 44158 34078 44210 34130
rect 46510 34078 46562 34130
rect 47182 34078 47234 34130
rect 49870 34078 49922 34130
rect 49982 34078 50034 34130
rect 51886 34078 51938 34130
rect 52334 34078 52386 34130
rect 53342 34078 53394 34130
rect 53790 34078 53842 34130
rect 54014 34078 54066 34130
rect 54462 34078 54514 34130
rect 54686 34078 54738 34130
rect 54910 34078 54962 34130
rect 55022 34078 55074 34130
rect 55582 34078 55634 34130
rect 62078 34078 62130 34130
rect 4062 33966 4114 34018
rect 7534 33966 7586 34018
rect 8990 33966 9042 34018
rect 16830 33966 16882 34018
rect 18398 33966 18450 34018
rect 23214 33966 23266 34018
rect 24110 33966 24162 34018
rect 24334 33966 24386 34018
rect 25678 33966 25730 34018
rect 26462 33966 26514 34018
rect 28142 33966 28194 34018
rect 28814 33966 28866 34018
rect 30830 33966 30882 34018
rect 31390 33966 31442 34018
rect 38222 33966 38274 34018
rect 38334 33966 38386 34018
rect 42254 33966 42306 34018
rect 46286 33966 46338 34018
rect 48078 33966 48130 34018
rect 53566 33966 53618 34018
rect 53902 33966 53954 34018
rect 7086 33854 7138 33906
rect 9662 33854 9714 33906
rect 13246 33854 13298 33906
rect 21422 33854 21474 33906
rect 22878 33854 22930 33906
rect 23662 33854 23714 33906
rect 26686 33854 26738 33906
rect 27022 33854 27074 33906
rect 28030 33854 28082 33906
rect 29262 33854 29314 33906
rect 35310 33854 35362 33906
rect 39342 33854 39394 33906
rect 48190 33854 48242 33906
rect 55582 33854 55634 33906
rect 58830 33854 58882 33906
rect 59614 33854 59666 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 1934 33518 1986 33570
rect 17726 33518 17778 33570
rect 25454 33518 25506 33570
rect 30382 33518 30434 33570
rect 37102 33518 37154 33570
rect 37326 33518 37378 33570
rect 37886 33518 37938 33570
rect 40574 33518 40626 33570
rect 46062 33518 46114 33570
rect 50766 33518 50818 33570
rect 51326 33518 51378 33570
rect 53118 33518 53170 33570
rect 54462 33518 54514 33570
rect 7086 33406 7138 33458
rect 10558 33406 10610 33458
rect 12798 33406 12850 33458
rect 14142 33406 14194 33458
rect 19070 33406 19122 33458
rect 21646 33406 21698 33458
rect 21982 33406 22034 33458
rect 28254 33406 28306 33458
rect 30046 33406 30098 33458
rect 32734 33406 32786 33458
rect 36206 33406 36258 33458
rect 47406 33406 47458 33458
rect 53454 33406 53506 33458
rect 55470 33406 55522 33458
rect 4062 33294 4114 33346
rect 5630 33294 5682 33346
rect 6190 33294 6242 33346
rect 7198 33294 7250 33346
rect 10222 33294 10274 33346
rect 11006 33294 11058 33346
rect 12014 33294 12066 33346
rect 12350 33294 12402 33346
rect 14030 33294 14082 33346
rect 14590 33294 14642 33346
rect 16046 33294 16098 33346
rect 16830 33294 16882 33346
rect 18622 33294 18674 33346
rect 19294 33294 19346 33346
rect 20526 33294 20578 33346
rect 20750 33294 20802 33346
rect 22542 33294 22594 33346
rect 25230 33294 25282 33346
rect 29262 33294 29314 33346
rect 29934 33294 29986 33346
rect 31726 33294 31778 33346
rect 33070 33294 33122 33346
rect 34414 33294 34466 33346
rect 35086 33294 35138 33346
rect 35422 33294 35474 33346
rect 38222 33294 38274 33346
rect 39678 33294 39730 33346
rect 40126 33294 40178 33346
rect 41358 33294 41410 33346
rect 44158 33294 44210 33346
rect 45054 33294 45106 33346
rect 45726 33294 45778 33346
rect 51550 33294 51602 33346
rect 52782 33294 52834 33346
rect 53342 33294 53394 33346
rect 53902 33294 53954 33346
rect 54126 33294 54178 33346
rect 55022 33294 55074 33346
rect 56478 33294 56530 33346
rect 56814 33294 56866 33346
rect 58158 33294 58210 33346
rect 60734 33294 60786 33346
rect 61742 33294 61794 33346
rect 6862 33182 6914 33234
rect 9550 33182 9602 33234
rect 10782 33182 10834 33234
rect 11342 33182 11394 33234
rect 12686 33182 12738 33234
rect 17390 33182 17442 33234
rect 18510 33182 18562 33234
rect 19070 33182 19122 33234
rect 21870 33182 21922 33234
rect 23214 33182 23266 33234
rect 25790 33182 25842 33234
rect 26014 33182 26066 33234
rect 27134 33182 27186 33234
rect 33294 33182 33346 33234
rect 33742 33182 33794 33234
rect 34302 33182 34354 33234
rect 35870 33182 35922 33234
rect 37662 33182 37714 33234
rect 42254 33182 42306 33234
rect 45166 33182 45218 33234
rect 46846 33182 46898 33234
rect 48750 33182 48802 33234
rect 53566 33182 53618 33234
rect 59390 33182 59442 33234
rect 60510 33182 60562 33234
rect 61966 33182 62018 33234
rect 5182 33070 5234 33122
rect 7758 33070 7810 33122
rect 10222 33070 10274 33122
rect 11454 33070 11506 33122
rect 13806 33070 13858 33122
rect 14254 33070 14306 33122
rect 20190 33070 20242 33122
rect 22094 33070 22146 33122
rect 25006 33070 25058 33122
rect 25566 33070 25618 33122
rect 33854 33070 33906 33122
rect 36094 33070 36146 33122
rect 36990 33070 37042 33122
rect 46510 33070 46562 33122
rect 47854 33070 47906 33122
rect 61406 33070 61458 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 8990 32734 9042 32786
rect 9886 32734 9938 32786
rect 11230 32734 11282 32786
rect 22766 32734 22818 32786
rect 23438 32734 23490 32786
rect 28254 32734 28306 32786
rect 28814 32734 28866 32786
rect 30494 32734 30546 32786
rect 31502 32734 31554 32786
rect 33518 32734 33570 32786
rect 34526 32734 34578 32786
rect 38334 32734 38386 32786
rect 38446 32734 38498 32786
rect 38782 32734 38834 32786
rect 39790 32734 39842 32786
rect 40238 32734 40290 32786
rect 40462 32734 40514 32786
rect 43598 32734 43650 32786
rect 48974 32734 49026 32786
rect 49198 32734 49250 32786
rect 54462 32734 54514 32786
rect 56030 32734 56082 32786
rect 57486 32734 57538 32786
rect 58382 32734 58434 32786
rect 3054 32622 3106 32674
rect 4846 32622 4898 32674
rect 15598 32622 15650 32674
rect 16270 32622 16322 32674
rect 16606 32622 16658 32674
rect 17950 32622 18002 32674
rect 22206 32622 22258 32674
rect 22878 32622 22930 32674
rect 24558 32622 24610 32674
rect 27918 32622 27970 32674
rect 36206 32622 36258 32674
rect 38558 32622 38610 32674
rect 42366 32622 42418 32674
rect 44158 32622 44210 32674
rect 44494 32622 44546 32674
rect 46062 32622 46114 32674
rect 48862 32622 48914 32674
rect 51998 32622 52050 32674
rect 57934 32622 57986 32674
rect 61630 32622 61682 32674
rect 2046 32510 2098 32562
rect 2382 32510 2434 32562
rect 3614 32510 3666 32562
rect 4062 32510 4114 32562
rect 5854 32510 5906 32562
rect 6190 32510 6242 32562
rect 7534 32510 7586 32562
rect 9550 32510 9602 32562
rect 9886 32510 9938 32562
rect 10222 32510 10274 32562
rect 13358 32510 13410 32562
rect 14814 32510 14866 32562
rect 15486 32510 15538 32562
rect 16046 32510 16098 32562
rect 16494 32510 16546 32562
rect 17614 32510 17666 32562
rect 19070 32510 19122 32562
rect 19294 32510 19346 32562
rect 21534 32510 21586 32562
rect 22318 32510 22370 32562
rect 24446 32510 24498 32562
rect 26238 32510 26290 32562
rect 26462 32510 26514 32562
rect 27022 32510 27074 32562
rect 28926 32510 28978 32562
rect 29374 32510 29426 32562
rect 31838 32510 31890 32562
rect 32062 32510 32114 32562
rect 33070 32510 33122 32562
rect 33294 32510 33346 32562
rect 33854 32510 33906 32562
rect 37774 32510 37826 32562
rect 37998 32510 38050 32562
rect 39454 32510 39506 32562
rect 40126 32510 40178 32562
rect 41694 32510 41746 32562
rect 42254 32510 42306 32562
rect 42702 32510 42754 32562
rect 44718 32510 44770 32562
rect 45390 32510 45442 32562
rect 50542 32510 50594 32562
rect 51214 32510 51266 32562
rect 54686 32510 54738 32562
rect 57038 32510 57090 32562
rect 57710 32510 57762 32562
rect 58494 32510 58546 32562
rect 60174 32510 60226 32562
rect 60510 32510 60562 32562
rect 61070 32510 61122 32562
rect 2270 32398 2322 32450
rect 4510 32398 4562 32450
rect 8542 32398 8594 32450
rect 12574 32398 12626 32450
rect 13134 32398 13186 32450
rect 14030 32398 14082 32450
rect 16158 32398 16210 32450
rect 26686 32398 26738 32450
rect 32510 32398 32562 32450
rect 37102 32398 37154 32450
rect 39230 32398 39282 32450
rect 48190 32398 48242 32450
rect 49534 32398 49586 32450
rect 50430 32398 50482 32450
rect 54126 32398 54178 32450
rect 55470 32398 55522 32450
rect 56926 32398 56978 32450
rect 14478 32286 14530 32338
rect 17502 32286 17554 32338
rect 21198 32286 21250 32338
rect 23774 32286 23826 32338
rect 33630 32286 33682 32338
rect 37438 32286 37490 32338
rect 43934 32286 43986 32338
rect 49534 32286 49586 32338
rect 49982 32286 50034 32338
rect 50206 32286 50258 32338
rect 55694 32286 55746 32338
rect 57374 32286 57426 32338
rect 58382 32286 58434 32338
rect 61294 32286 61346 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 2718 31950 2770 32002
rect 3502 31950 3554 32002
rect 6190 31950 6242 32002
rect 10222 31950 10274 32002
rect 17502 31950 17554 32002
rect 22318 31950 22370 32002
rect 33294 31950 33346 32002
rect 34190 31950 34242 32002
rect 51326 31950 51378 32002
rect 52110 31950 52162 32002
rect 57150 31950 57202 32002
rect 61070 31950 61122 32002
rect 1934 31838 1986 31890
rect 3726 31838 3778 31890
rect 4734 31838 4786 31890
rect 8542 31838 8594 31890
rect 9214 31838 9266 31890
rect 9886 31838 9938 31890
rect 19518 31838 19570 31890
rect 28030 31838 28082 31890
rect 28366 31838 28418 31890
rect 34974 31838 35026 31890
rect 36430 31838 36482 31890
rect 43598 31838 43650 31890
rect 45726 31838 45778 31890
rect 47182 31838 47234 31890
rect 51998 31838 52050 31890
rect 57486 31838 57538 31890
rect 2158 31726 2210 31778
rect 2382 31726 2434 31778
rect 2718 31726 2770 31778
rect 4846 31726 4898 31778
rect 5630 31726 5682 31778
rect 5966 31726 6018 31778
rect 6190 31726 6242 31778
rect 7086 31726 7138 31778
rect 7982 31726 8034 31778
rect 8318 31726 8370 31778
rect 8990 31726 9042 31778
rect 9438 31726 9490 31778
rect 11566 31726 11618 31778
rect 13470 31726 13522 31778
rect 14366 31726 14418 31778
rect 14478 31726 14530 31778
rect 16494 31726 16546 31778
rect 16830 31726 16882 31778
rect 17838 31726 17890 31778
rect 18062 31726 18114 31778
rect 18510 31726 18562 31778
rect 20190 31726 20242 31778
rect 21534 31726 21586 31778
rect 22542 31726 22594 31778
rect 22766 31726 22818 31778
rect 22878 31726 22930 31778
rect 23998 31726 24050 31778
rect 24334 31726 24386 31778
rect 25230 31726 25282 31778
rect 28478 31726 28530 31778
rect 33406 31726 33458 31778
rect 34302 31726 34354 31778
rect 34750 31726 34802 31778
rect 35534 31726 35586 31778
rect 35758 31726 35810 31778
rect 35982 31726 36034 31778
rect 37998 31726 38050 31778
rect 38222 31726 38274 31778
rect 38558 31726 38610 31778
rect 39678 31726 39730 31778
rect 40686 31726 40738 31778
rect 45278 31726 45330 31778
rect 46622 31726 46674 31778
rect 47518 31726 47570 31778
rect 53678 31726 53730 31778
rect 54574 31726 54626 31778
rect 60510 31726 60562 31778
rect 61406 31726 61458 31778
rect 61630 31726 61682 31778
rect 3278 31614 3330 31666
rect 6862 31614 6914 31666
rect 7422 31614 7474 31666
rect 7758 31614 7810 31666
rect 8094 31614 8146 31666
rect 11118 31614 11170 31666
rect 11790 31614 11842 31666
rect 12686 31614 12738 31666
rect 18734 31614 18786 31666
rect 21310 31614 21362 31666
rect 23102 31614 23154 31666
rect 23550 31614 23602 31666
rect 23662 31614 23714 31666
rect 24446 31614 24498 31666
rect 24558 31614 24610 31666
rect 25902 31614 25954 31666
rect 29710 31614 29762 31666
rect 31166 31614 31218 31666
rect 32734 31614 32786 31666
rect 32958 31614 33010 31666
rect 34526 31614 34578 31666
rect 36318 31614 36370 31666
rect 37326 31614 37378 31666
rect 37662 31614 37714 31666
rect 38894 31614 38946 31666
rect 41134 31614 41186 31666
rect 42254 31614 42306 31666
rect 44158 31614 44210 31666
rect 49310 31614 49362 31666
rect 53006 31614 53058 31666
rect 53342 31614 53394 31666
rect 55358 31614 55410 31666
rect 58830 31614 58882 31666
rect 61854 31614 61906 31666
rect 2942 31502 2994 31554
rect 6414 31502 6466 31554
rect 6974 31502 7026 31554
rect 9102 31502 9154 31554
rect 10110 31502 10162 31554
rect 11006 31502 11058 31554
rect 12126 31502 12178 31554
rect 23326 31502 23378 31554
rect 24670 31502 24722 31554
rect 29150 31502 29202 31554
rect 30270 31502 30322 31554
rect 32286 31502 32338 31554
rect 33518 31502 33570 31554
rect 35870 31502 35922 31554
rect 46062 31502 46114 31554
rect 48190 31502 48242 31554
rect 52670 31502 52722 31554
rect 54462 31502 54514 31554
rect 59950 31502 60002 31554
rect 61518 31502 61570 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 2270 31166 2322 31218
rect 2494 31166 2546 31218
rect 6974 31166 7026 31218
rect 7646 31166 7698 31218
rect 8542 31166 8594 31218
rect 8766 31166 8818 31218
rect 10558 31166 10610 31218
rect 11678 31166 11730 31218
rect 12574 31166 12626 31218
rect 12798 31166 12850 31218
rect 15150 31166 15202 31218
rect 2046 31054 2098 31106
rect 2158 31054 2210 31106
rect 5630 31054 5682 31106
rect 13358 31054 13410 31106
rect 14814 31054 14866 31106
rect 15374 31110 15426 31162
rect 16270 31166 16322 31218
rect 16382 31166 16434 31218
rect 17502 31166 17554 31218
rect 18846 31166 18898 31218
rect 20190 31166 20242 31218
rect 20862 31166 20914 31218
rect 24558 31166 24610 31218
rect 27694 31166 27746 31218
rect 30382 31166 30434 31218
rect 30718 31166 30770 31218
rect 31166 31166 31218 31218
rect 33070 31166 33122 31218
rect 33406 31166 33458 31218
rect 33854 31166 33906 31218
rect 37550 31166 37602 31218
rect 39678 31166 39730 31218
rect 41470 31166 41522 31218
rect 43710 31166 43762 31218
rect 44830 31166 44882 31218
rect 46510 31166 46562 31218
rect 47070 31166 47122 31218
rect 47630 31166 47682 31218
rect 50542 31166 50594 31218
rect 51102 31166 51154 31218
rect 57598 31166 57650 31218
rect 15486 31054 15538 31106
rect 15710 31054 15762 31106
rect 17838 31054 17890 31106
rect 22542 31054 22594 31106
rect 23102 31054 23154 31106
rect 24110 31054 24162 31106
rect 29934 31054 29986 31106
rect 32174 31054 32226 31106
rect 38782 31054 38834 31106
rect 45614 31054 45666 31106
rect 45950 31054 46002 31106
rect 47742 31054 47794 31106
rect 49310 31054 49362 31106
rect 51774 31054 51826 31106
rect 52446 31054 52498 31106
rect 53566 31054 53618 31106
rect 53902 31054 53954 31106
rect 54238 31054 54290 31106
rect 56030 31054 56082 31106
rect 56590 31054 56642 31106
rect 58158 31054 58210 31106
rect 58718 31054 58770 31106
rect 3166 30942 3218 30994
rect 3726 30942 3778 30994
rect 5966 30942 6018 30994
rect 7870 30942 7922 30994
rect 8094 30942 8146 30994
rect 8318 30942 8370 30994
rect 8878 30942 8930 30994
rect 12462 30942 12514 30994
rect 12910 30942 12962 30994
rect 13694 30942 13746 30994
rect 16494 30942 16546 30994
rect 16942 30942 16994 30994
rect 20750 30942 20802 30994
rect 21086 30942 21138 30994
rect 21310 30942 21362 30994
rect 22094 30942 22146 30994
rect 23214 30942 23266 30994
rect 23550 30942 23602 30994
rect 23886 30942 23938 30994
rect 24334 30942 24386 30994
rect 24670 30942 24722 30994
rect 25790 30942 25842 30994
rect 27358 30942 27410 30994
rect 28926 30942 28978 30994
rect 29598 30942 29650 30994
rect 31502 30942 31554 30994
rect 32286 30942 32338 30994
rect 34190 30930 34242 30982
rect 41806 30942 41858 30994
rect 42254 30942 42306 30994
rect 46174 30942 46226 30994
rect 47406 30942 47458 30994
rect 48190 30942 48242 30994
rect 51438 30942 51490 30994
rect 52110 30942 52162 30994
rect 54574 30942 54626 30994
rect 55806 30942 55858 30994
rect 56814 30942 56866 30994
rect 57262 30942 57314 30994
rect 57934 30942 57986 30994
rect 59614 30942 59666 30994
rect 3838 30830 3890 30882
rect 6862 30830 6914 30882
rect 7758 30830 7810 30882
rect 15934 30830 15986 30882
rect 22430 30830 22482 30882
rect 23662 30830 23714 30882
rect 26126 30830 26178 30882
rect 27022 30830 27074 30882
rect 27806 30830 27858 30882
rect 28702 30830 28754 30882
rect 34974 30830 35026 30882
rect 37102 30830 37154 30882
rect 40126 30830 40178 30882
rect 40910 30830 40962 30882
rect 47742 30830 47794 30882
rect 53006 30830 53058 30882
rect 53230 30830 53282 30882
rect 55022 30830 55074 30882
rect 57038 30830 57090 30882
rect 59278 30830 59330 30882
rect 61966 30830 62018 30882
rect 14590 30718 14642 30770
rect 25678 30718 25730 30770
rect 29486 30718 29538 30770
rect 55470 30718 55522 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 4958 30382 5010 30434
rect 15150 30382 15202 30434
rect 19518 30382 19570 30434
rect 24670 30382 24722 30434
rect 32062 30382 32114 30434
rect 43262 30382 43314 30434
rect 43934 30382 43986 30434
rect 50878 30382 50930 30434
rect 56702 30382 56754 30434
rect 4622 30270 4674 30322
rect 10670 30270 10722 30322
rect 16718 30270 16770 30322
rect 25230 30270 25282 30322
rect 30942 30270 30994 30322
rect 34302 30270 34354 30322
rect 39342 30270 39394 30322
rect 4734 30158 4786 30210
rect 5742 30158 5794 30210
rect 6078 30158 6130 30210
rect 7310 30158 7362 30210
rect 7758 30158 7810 30210
rect 11230 30158 11282 30210
rect 11566 30158 11618 30210
rect 12798 30158 12850 30210
rect 13806 30158 13858 30210
rect 14254 30158 14306 30210
rect 15038 30158 15090 30210
rect 16606 30158 16658 30210
rect 19854 30158 19906 30210
rect 20302 30158 20354 30210
rect 21422 30158 21474 30210
rect 22654 30158 22706 30210
rect 24558 30158 24610 30210
rect 26014 30158 26066 30210
rect 28478 30158 28530 30210
rect 29710 30158 29762 30210
rect 31166 30158 31218 30210
rect 34190 30158 34242 30210
rect 34414 30158 34466 30210
rect 34750 30158 34802 30210
rect 34974 30158 35026 30210
rect 35646 30158 35698 30210
rect 36094 30158 36146 30210
rect 37214 30158 37266 30210
rect 37662 30158 37714 30210
rect 38558 30158 38610 30210
rect 41470 30158 41522 30210
rect 43038 30158 43090 30210
rect 44158 30158 44210 30210
rect 48638 30158 48690 30210
rect 49422 30158 49474 30210
rect 51214 30158 51266 30210
rect 51886 30158 51938 30210
rect 54462 30158 54514 30210
rect 55358 30158 55410 30210
rect 56030 30158 56082 30210
rect 56478 30158 56530 30210
rect 56926 30158 56978 30210
rect 57374 30158 57426 30210
rect 61518 30158 61570 30210
rect 2270 30046 2322 30098
rect 6302 30046 6354 30098
rect 6638 30046 6690 30098
rect 7422 30046 7474 30098
rect 8542 30046 8594 30098
rect 11342 30046 11394 30098
rect 12126 30046 12178 30098
rect 12350 30046 12402 30098
rect 13022 30046 13074 30098
rect 15598 30046 15650 30098
rect 18958 30046 19010 30098
rect 19294 30046 19346 30098
rect 20750 30046 20802 30098
rect 23886 30046 23938 30098
rect 29934 30046 29986 30098
rect 41918 30046 41970 30098
rect 47630 30046 47682 30098
rect 49758 30046 49810 30098
rect 51998 30046 52050 30098
rect 53342 30046 53394 30098
rect 55582 30046 55634 30098
rect 61854 30046 61906 30098
rect 62190 30046 62242 30098
rect 3502 29934 3554 29986
rect 20526 29934 20578 29986
rect 20862 29934 20914 29986
rect 25678 29934 25730 29986
rect 26126 29934 26178 29986
rect 26350 29934 26402 29986
rect 27358 29934 27410 29986
rect 33182 29934 33234 29986
rect 33406 29934 33458 29986
rect 33630 29934 33682 29986
rect 35086 29934 35138 29986
rect 35310 29934 35362 29986
rect 35758 29934 35810 29986
rect 35982 29934 36034 29986
rect 37998 29934 38050 29986
rect 38894 29934 38946 29986
rect 39790 29934 39842 29986
rect 40126 29934 40178 29986
rect 40462 29934 40514 29986
rect 40798 29934 40850 29986
rect 42478 29934 42530 29986
rect 43598 29934 43650 29986
rect 45054 29934 45106 29986
rect 46062 29934 46114 29986
rect 47182 29934 47234 29986
rect 50542 29934 50594 29986
rect 55022 29934 55074 29986
rect 55806 29934 55858 29986
rect 58718 29934 58770 29986
rect 59838 29934 59890 29986
rect 60510 29934 60562 29986
rect 60622 29934 60674 29986
rect 60734 29934 60786 29986
rect 60958 29934 61010 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 7982 29598 8034 29650
rect 9886 29598 9938 29650
rect 12350 29598 12402 29650
rect 14142 29598 14194 29650
rect 15822 29598 15874 29650
rect 16382 29598 16434 29650
rect 25566 29598 25618 29650
rect 25790 29598 25842 29650
rect 31950 29598 32002 29650
rect 32398 29598 32450 29650
rect 33406 29598 33458 29650
rect 36654 29598 36706 29650
rect 38446 29598 38498 29650
rect 41470 29598 41522 29650
rect 42366 29598 42418 29650
rect 43822 29598 43874 29650
rect 46958 29598 47010 29650
rect 49310 29598 49362 29650
rect 3838 29486 3890 29538
rect 5518 29486 5570 29538
rect 7870 29486 7922 29538
rect 10782 29486 10834 29538
rect 15038 29486 15090 29538
rect 15710 29486 15762 29538
rect 16494 29486 16546 29538
rect 17950 29486 18002 29538
rect 25454 29486 25506 29538
rect 28814 29486 28866 29538
rect 31278 29486 31330 29538
rect 33294 29486 33346 29538
rect 33854 29486 33906 29538
rect 34526 29486 34578 29538
rect 36542 29486 36594 29538
rect 38110 29486 38162 29538
rect 39006 29486 39058 29538
rect 48078 29486 48130 29538
rect 50206 29486 50258 29538
rect 52334 29486 52386 29538
rect 55918 29486 55970 29538
rect 56702 29486 56754 29538
rect 58382 29486 58434 29538
rect 61294 29486 61346 29538
rect 4510 29374 4562 29426
rect 7758 29374 7810 29426
rect 8430 29374 8482 29426
rect 8990 29374 9042 29426
rect 9550 29374 9602 29426
rect 15262 29374 15314 29426
rect 16046 29374 16098 29426
rect 16270 29374 16322 29426
rect 16942 29374 16994 29426
rect 17390 29374 17442 29426
rect 17726 29374 17778 29426
rect 18174 29374 18226 29426
rect 18734 29374 18786 29426
rect 19854 29374 19906 29426
rect 20526 29374 20578 29426
rect 20750 29374 20802 29426
rect 22206 29374 22258 29426
rect 23102 29374 23154 29426
rect 23998 29374 24050 29426
rect 24222 29374 24274 29426
rect 26238 29374 26290 29426
rect 26798 29374 26850 29426
rect 28702 29374 28754 29426
rect 29038 29374 29090 29426
rect 30494 29374 30546 29426
rect 31166 29374 31218 29426
rect 32510 29374 32562 29426
rect 33182 29374 33234 29426
rect 34750 29374 34802 29426
rect 35534 29374 35586 29426
rect 35982 29374 36034 29426
rect 36206 29374 36258 29426
rect 36878 29374 36930 29426
rect 37214 29374 37266 29426
rect 39678 29374 39730 29426
rect 40126 29374 40178 29426
rect 40350 29374 40402 29426
rect 41918 29374 41970 29426
rect 42702 29374 42754 29426
rect 42926 29374 42978 29426
rect 44158 29374 44210 29426
rect 46286 29374 46338 29426
rect 47294 29374 47346 29426
rect 47854 29374 47906 29426
rect 53230 29374 53282 29426
rect 54574 29374 54626 29426
rect 55134 29374 55186 29426
rect 55470 29374 55522 29426
rect 55806 29374 55858 29426
rect 56590 29374 56642 29426
rect 57598 29374 57650 29426
rect 58046 29374 58098 29426
rect 58830 29374 58882 29426
rect 60286 29374 60338 29426
rect 61406 29374 61458 29426
rect 1710 29262 1762 29314
rect 6974 29262 7026 29314
rect 13358 29262 13410 29314
rect 13694 29262 13746 29314
rect 17950 29262 18002 29314
rect 23438 29262 23490 29314
rect 30158 29262 30210 29314
rect 35198 29262 35250 29314
rect 35310 29262 35362 29314
rect 40238 29262 40290 29314
rect 41022 29262 41074 29314
rect 43262 29262 43314 29314
rect 44718 29262 44770 29314
rect 45054 29262 45106 29314
rect 46510 29262 46562 29314
rect 48750 29262 48802 29314
rect 51998 29262 52050 29314
rect 53678 29262 53730 29314
rect 54910 29262 54962 29314
rect 14478 29150 14530 29202
rect 21758 29150 21810 29202
rect 22766 29150 22818 29202
rect 38782 29150 38834 29202
rect 42030 29150 42082 29202
rect 45278 29150 45330 29202
rect 45614 29150 45666 29202
rect 45950 29150 46002 29202
rect 48974 29150 49026 29202
rect 55918 29150 55970 29202
rect 56702 29150 56754 29202
rect 57262 29150 57314 29202
rect 61966 29150 62018 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 2382 28814 2434 28866
rect 15598 28814 15650 28866
rect 20302 28814 20354 28866
rect 25006 28814 25058 28866
rect 31054 28814 31106 28866
rect 36430 28814 36482 28866
rect 37326 28814 37378 28866
rect 40686 28814 40738 28866
rect 47070 28814 47122 28866
rect 49870 28814 49922 28866
rect 51326 28814 51378 28866
rect 52782 28814 52834 28866
rect 55358 28814 55410 28866
rect 58158 28814 58210 28866
rect 1710 28702 1762 28754
rect 6974 28702 7026 28754
rect 9102 28702 9154 28754
rect 10558 28702 10610 28754
rect 13806 28702 13858 28754
rect 14702 28702 14754 28754
rect 18958 28702 19010 28754
rect 19742 28702 19794 28754
rect 24558 28702 24610 28754
rect 29150 28702 29202 28754
rect 30494 28702 30546 28754
rect 33070 28702 33122 28754
rect 35198 28702 35250 28754
rect 37214 28702 37266 28754
rect 37774 28702 37826 28754
rect 40126 28702 40178 28754
rect 45726 28702 45778 28754
rect 56254 28702 56306 28754
rect 57150 28702 57202 28754
rect 60734 28702 60786 28754
rect 1822 28590 1874 28642
rect 5966 28590 6018 28642
rect 6190 28590 6242 28642
rect 9774 28590 9826 28642
rect 12798 28590 12850 28642
rect 14142 28590 14194 28642
rect 14366 28590 14418 28642
rect 16382 28590 16434 28642
rect 16942 28590 16994 28642
rect 17278 28590 17330 28642
rect 19070 28590 19122 28642
rect 19518 28590 19570 28642
rect 19966 28590 20018 28642
rect 20862 28590 20914 28642
rect 21758 28590 21810 28642
rect 28478 28590 28530 28642
rect 29710 28590 29762 28642
rect 30382 28590 30434 28642
rect 31166 28590 31218 28642
rect 32958 28590 33010 28642
rect 34974 28590 35026 28642
rect 35534 28590 35586 28642
rect 35758 28590 35810 28642
rect 35982 28590 36034 28642
rect 36990 28590 37042 28642
rect 38222 28590 38274 28642
rect 39230 28590 39282 28642
rect 39790 28590 39842 28642
rect 39902 28590 39954 28642
rect 40350 28590 40402 28642
rect 41470 28590 41522 28642
rect 42702 28590 42754 28642
rect 43934 28590 43986 28642
rect 45166 28590 45218 28642
rect 45390 28590 45442 28642
rect 46734 28590 46786 28642
rect 47070 28590 47122 28642
rect 50542 28590 50594 28642
rect 50990 28590 51042 28642
rect 51774 28590 51826 28642
rect 53118 28590 53170 28642
rect 55022 28590 55074 28642
rect 55582 28590 55634 28642
rect 56590 28590 56642 28642
rect 57374 28590 57426 28642
rect 60510 28590 60562 28642
rect 61182 28590 61234 28642
rect 61630 28590 61682 28642
rect 62190 28590 62242 28642
rect 4398 28478 4450 28530
rect 5630 28478 5682 28530
rect 5742 28478 5794 28530
rect 9438 28478 9490 28530
rect 11342 28478 11394 28530
rect 14814 28478 14866 28530
rect 15822 28478 15874 28530
rect 22430 28478 22482 28530
rect 26238 28478 26290 28530
rect 27806 28478 27858 28530
rect 28366 28478 28418 28530
rect 31726 28478 31778 28530
rect 38334 28478 38386 28530
rect 41358 28478 41410 28530
rect 46062 28478 46114 28530
rect 46510 28478 46562 28530
rect 47966 28478 48018 28530
rect 50206 28478 50258 28530
rect 52110 28478 52162 28530
rect 53342 28478 53394 28530
rect 53902 28478 53954 28530
rect 54350 28478 54402 28530
rect 54686 28478 54738 28530
rect 55806 28478 55858 28530
rect 57710 28478 57762 28530
rect 59278 28478 59330 28530
rect 60846 28478 60898 28530
rect 14590 28366 14642 28418
rect 18846 28366 18898 28418
rect 28030 28366 28082 28418
rect 34638 28366 34690 28418
rect 39118 28366 39170 28418
rect 44830 28366 44882 28418
rect 45838 28366 45890 28418
rect 47294 28366 47346 28418
rect 55022 28366 55074 28418
rect 60734 28366 60786 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 2270 28030 2322 28082
rect 3166 28030 3218 28082
rect 4286 28030 4338 28082
rect 6302 28030 6354 28082
rect 7646 28030 7698 28082
rect 10558 28030 10610 28082
rect 21422 28030 21474 28082
rect 21646 28030 21698 28082
rect 22654 28030 22706 28082
rect 24558 28030 24610 28082
rect 25230 28030 25282 28082
rect 27582 28030 27634 28082
rect 31166 28030 31218 28082
rect 31390 28030 31442 28082
rect 32510 28030 32562 28082
rect 33070 28030 33122 28082
rect 33182 28030 33234 28082
rect 33854 28030 33906 28082
rect 34078 28030 34130 28082
rect 36654 28030 36706 28082
rect 37774 28030 37826 28082
rect 38446 28030 38498 28082
rect 38558 28030 38610 28082
rect 38670 28030 38722 28082
rect 43150 28030 43202 28082
rect 48862 28030 48914 28082
rect 54126 28030 54178 28082
rect 56814 28030 56866 28082
rect 56926 28030 56978 28082
rect 61518 28030 61570 28082
rect 3502 27918 3554 27970
rect 4510 27918 4562 27970
rect 4622 27918 4674 27970
rect 5406 27918 5458 27970
rect 11678 27918 11730 27970
rect 12462 27918 12514 27970
rect 13358 27918 13410 27970
rect 14702 27918 14754 27970
rect 16270 27918 16322 27970
rect 23438 27918 23490 27970
rect 24670 27918 24722 27970
rect 26014 27918 26066 27970
rect 26350 27918 26402 27970
rect 28590 27918 28642 27970
rect 32398 27918 32450 27970
rect 34750 27918 34802 27970
rect 34862 27918 34914 27970
rect 40014 27918 40066 27970
rect 41022 27918 41074 27970
rect 44046 27918 44098 27970
rect 47518 27918 47570 27970
rect 50206 27918 50258 27970
rect 52110 27918 52162 27970
rect 52670 27918 52722 27970
rect 55694 27918 55746 27970
rect 57038 27918 57090 27970
rect 1934 27806 1986 27858
rect 2606 27806 2658 27858
rect 3726 27806 3778 27858
rect 4958 27806 5010 27858
rect 5630 27806 5682 27858
rect 12238 27806 12290 27858
rect 13806 27806 13858 27858
rect 14926 27806 14978 27858
rect 15934 27806 15986 27858
rect 17502 27806 17554 27858
rect 18622 27806 18674 27858
rect 19630 27806 19682 27858
rect 20974 27806 21026 27858
rect 21870 27806 21922 27858
rect 22206 27806 22258 27858
rect 22542 27806 22594 27858
rect 22766 27806 22818 27858
rect 23214 27806 23266 27858
rect 23662 27806 23714 27858
rect 24222 27806 24274 27858
rect 24334 27806 24386 27858
rect 25342 27806 25394 27858
rect 25678 27806 25730 27858
rect 26574 27806 26626 27858
rect 26798 27806 26850 27858
rect 27694 27806 27746 27858
rect 30382 27806 30434 27858
rect 31614 27806 31666 27858
rect 31950 27806 32002 27858
rect 33294 27806 33346 27858
rect 33630 27806 33682 27858
rect 34190 27806 34242 27858
rect 35534 27806 35586 27858
rect 35758 27806 35810 27858
rect 35982 27806 36034 27858
rect 36430 27806 36482 27858
rect 37326 27806 37378 27858
rect 37550 27806 37602 27858
rect 37998 27806 38050 27858
rect 40126 27806 40178 27858
rect 41134 27806 41186 27858
rect 42030 27806 42082 27858
rect 42814 27806 42866 27858
rect 44158 27806 44210 27858
rect 45614 27806 45666 27858
rect 46734 27806 46786 27858
rect 47294 27806 47346 27858
rect 51550 27806 51602 27858
rect 51998 27806 52050 27858
rect 52446 27806 52498 27858
rect 53006 27806 53058 27858
rect 53566 27806 53618 27858
rect 54798 27806 54850 27858
rect 55806 27806 55858 27858
rect 57262 27806 57314 27858
rect 57598 27806 57650 27858
rect 58158 27806 58210 27858
rect 58718 27806 58770 27858
rect 59726 27806 59778 27858
rect 4622 27694 4674 27746
rect 9102 27694 9154 27746
rect 14254 27694 14306 27746
rect 16046 27694 16098 27746
rect 16718 27694 16770 27746
rect 18286 27694 18338 27746
rect 20638 27694 20690 27746
rect 21758 27694 21810 27746
rect 31278 27694 31330 27746
rect 37886 27694 37938 27746
rect 41582 27694 41634 27746
rect 41694 27694 41746 27746
rect 43934 27694 43986 27746
rect 48078 27694 48130 27746
rect 51326 27694 51378 27746
rect 52558 27694 52610 27746
rect 52894 27694 52946 27746
rect 55246 27694 55298 27746
rect 55358 27694 55410 27746
rect 13022 27582 13074 27634
rect 16830 27582 16882 27634
rect 25454 27582 25506 27634
rect 26686 27582 26738 27634
rect 36766 27582 36818 27634
rect 39118 27582 39170 27634
rect 39454 27582 39506 27634
rect 46398 27582 46450 27634
rect 51998 27582 52050 27634
rect 58046 27582 58098 27634
rect 59390 27582 59442 27634
rect 60174 27582 60226 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 11342 27246 11394 27298
rect 11678 27246 11730 27298
rect 27694 27246 27746 27298
rect 44942 27246 44994 27298
rect 45390 27246 45442 27298
rect 45614 27246 45666 27298
rect 49758 27246 49810 27298
rect 50094 27246 50146 27298
rect 52110 27246 52162 27298
rect 53118 27246 53170 27298
rect 58270 27246 58322 27298
rect 59390 27246 59442 27298
rect 62078 27246 62130 27298
rect 2606 27134 2658 27186
rect 4398 27134 4450 27186
rect 6190 27134 6242 27186
rect 7758 27134 7810 27186
rect 9326 27134 9378 27186
rect 9886 27134 9938 27186
rect 10222 27134 10274 27186
rect 18062 27134 18114 27186
rect 19070 27134 19122 27186
rect 25118 27134 25170 27186
rect 26014 27134 26066 27186
rect 31166 27134 31218 27186
rect 33406 27134 33458 27186
rect 36318 27134 36370 27186
rect 37102 27134 37154 27186
rect 37774 27134 37826 27186
rect 41694 27134 41746 27186
rect 43150 27134 43202 27186
rect 50542 27134 50594 27186
rect 53902 27134 53954 27186
rect 56814 27134 56866 27186
rect 57822 27134 57874 27186
rect 60622 27134 60674 27186
rect 60846 27134 60898 27186
rect 62190 27134 62242 27186
rect 1934 27022 1986 27074
rect 3054 27022 3106 27074
rect 3390 27022 3442 27074
rect 3726 27022 3778 27074
rect 4622 27022 4674 27074
rect 5630 27022 5682 27074
rect 6974 27022 7026 27074
rect 7646 27022 7698 27074
rect 7870 27022 7922 27074
rect 10894 27022 10946 27074
rect 16158 27022 16210 27074
rect 16942 27022 16994 27074
rect 17614 27022 17666 27074
rect 20526 27022 20578 27074
rect 22430 27022 22482 27074
rect 22990 27022 23042 27074
rect 23662 27022 23714 27074
rect 24110 27022 24162 27074
rect 25006 27022 25058 27074
rect 25342 27022 25394 27074
rect 25902 27022 25954 27074
rect 26686 27022 26738 27074
rect 29934 27022 29986 27074
rect 31390 27022 31442 27074
rect 32174 27022 32226 27074
rect 32510 27022 32562 27074
rect 32958 27022 33010 27074
rect 34862 27022 34914 27074
rect 35758 27022 35810 27074
rect 37662 27022 37714 27074
rect 38670 27022 38722 27074
rect 39118 27022 39170 27074
rect 40686 27022 40738 27074
rect 41470 27022 41522 27074
rect 46174 27022 46226 27074
rect 47070 27022 47122 27074
rect 50430 27022 50482 27074
rect 50766 27022 50818 27074
rect 50990 27022 51042 27074
rect 51438 27022 51490 27074
rect 51662 27022 51714 27074
rect 51886 27022 51938 27074
rect 52894 27022 52946 27074
rect 53454 27022 53506 27074
rect 53790 27022 53842 27074
rect 54574 27022 54626 27074
rect 54686 27022 54738 27074
rect 55246 27022 55298 27074
rect 55470 27022 55522 27074
rect 55582 27022 55634 27074
rect 55806 27022 55858 27074
rect 56702 27022 56754 27074
rect 57486 27022 57538 27074
rect 58046 27022 58098 27074
rect 58830 27022 58882 27074
rect 61406 27022 61458 27074
rect 2158 26910 2210 26962
rect 4734 26910 4786 26962
rect 6750 26910 6802 26962
rect 7310 26910 7362 26962
rect 8206 26910 8258 26962
rect 11902 26910 11954 26962
rect 12462 26910 12514 26962
rect 14030 26910 14082 26962
rect 15486 26910 15538 26962
rect 18734 26910 18786 26962
rect 19294 26910 19346 26962
rect 19630 26910 19682 26962
rect 20750 26910 20802 26962
rect 21646 26910 21698 26962
rect 21982 26910 22034 26962
rect 23326 26910 23378 26962
rect 24334 26910 24386 26962
rect 24670 26910 24722 26962
rect 25678 26910 25730 26962
rect 27918 26910 27970 26962
rect 28478 26910 28530 26962
rect 29150 26910 29202 26962
rect 29262 26910 29314 26962
rect 30494 26910 30546 26962
rect 31502 26910 31554 26962
rect 33966 26910 34018 26962
rect 34526 26910 34578 26962
rect 35198 26910 35250 26962
rect 37550 26910 37602 26962
rect 40238 26910 40290 26962
rect 41022 26910 41074 26962
rect 43486 26910 43538 26962
rect 43598 26910 43650 26962
rect 6862 26798 6914 26850
rect 8542 26798 8594 26850
rect 8878 26798 8930 26850
rect 10558 26798 10610 26850
rect 27358 26798 27410 26850
rect 43710 26854 43762 26906
rect 44830 26910 44882 26962
rect 45054 26910 45106 26962
rect 48750 26910 48802 26962
rect 49870 26910 49922 26962
rect 51550 26910 51602 26962
rect 52670 26910 52722 26962
rect 56590 26910 56642 26962
rect 59838 26910 59890 26962
rect 29486 26798 29538 26850
rect 35534 26798 35586 26850
rect 43934 26798 43986 26850
rect 52782 26798 52834 26850
rect 54350 26798 54402 26850
rect 54798 26798 54850 26850
rect 61182 26798 61234 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 2046 26462 2098 26514
rect 11790 26462 11842 26514
rect 12238 26462 12290 26514
rect 13134 26462 13186 26514
rect 14590 26462 14642 26514
rect 14926 26462 14978 26514
rect 15038 26462 15090 26514
rect 16830 26462 16882 26514
rect 19630 26462 19682 26514
rect 26238 26462 26290 26514
rect 26350 26462 26402 26514
rect 26798 26462 26850 26514
rect 31726 26462 31778 26514
rect 33182 26462 33234 26514
rect 39902 26462 39954 26514
rect 40126 26462 40178 26514
rect 42926 26462 42978 26514
rect 48750 26462 48802 26514
rect 49758 26462 49810 26514
rect 57710 26462 57762 26514
rect 61630 26462 61682 26514
rect 61742 26462 61794 26514
rect 61966 26462 62018 26514
rect 1710 26350 1762 26402
rect 2942 26350 2994 26402
rect 5182 26350 5234 26402
rect 5630 26350 5682 26402
rect 9998 26350 10050 26402
rect 17950 26350 18002 26402
rect 21310 26350 21362 26402
rect 22318 26350 22370 26402
rect 23326 26350 23378 26402
rect 25790 26350 25842 26402
rect 26126 26350 26178 26402
rect 28030 26350 28082 26402
rect 33070 26350 33122 26402
rect 36318 26350 36370 26402
rect 41134 26350 41186 26402
rect 44718 26350 44770 26402
rect 46174 26350 46226 26402
rect 46622 26350 46674 26402
rect 50094 26350 50146 26402
rect 51662 26350 51714 26402
rect 55806 26350 55858 26402
rect 58606 26350 58658 26402
rect 62190 26350 62242 26402
rect 6750 26238 6802 26290
rect 6862 26238 6914 26290
rect 7310 26238 7362 26290
rect 7758 26238 7810 26290
rect 7982 26238 8034 26290
rect 8206 26238 8258 26290
rect 8542 26238 8594 26290
rect 8766 26238 8818 26290
rect 12574 26238 12626 26290
rect 13134 26238 13186 26290
rect 13694 26238 13746 26290
rect 13918 26238 13970 26290
rect 14814 26238 14866 26290
rect 15822 26238 15874 26290
rect 16270 26238 16322 26290
rect 22206 26238 22258 26290
rect 22542 26238 22594 26290
rect 25902 26238 25954 26290
rect 27918 26238 27970 26290
rect 29038 26238 29090 26290
rect 30494 26238 30546 26290
rect 31166 26238 31218 26290
rect 32174 26238 32226 26290
rect 34526 26238 34578 26290
rect 38110 26238 38162 26290
rect 39454 26238 39506 26290
rect 39678 26238 39730 26290
rect 41022 26238 41074 26290
rect 42254 26238 42306 26290
rect 42478 26238 42530 26290
rect 47294 26238 47346 26290
rect 47518 26238 47570 26290
rect 47742 26238 47794 26290
rect 48974 26238 49026 26290
rect 49646 26238 49698 26290
rect 49870 26238 49922 26290
rect 50990 26238 51042 26290
rect 54462 26238 54514 26290
rect 54798 26238 54850 26290
rect 56030 26238 56082 26290
rect 57038 26238 57090 26290
rect 59054 26238 59106 26290
rect 59726 26238 59778 26290
rect 60174 26238 60226 26290
rect 5854 26126 5906 26178
rect 7870 26126 7922 26178
rect 8430 26126 8482 26178
rect 12798 26126 12850 26178
rect 15374 26126 15426 26178
rect 31390 26126 31442 26178
rect 32398 26126 32450 26178
rect 33630 26126 33682 26178
rect 34190 26126 34242 26178
rect 34750 26126 34802 26178
rect 38558 26126 38610 26178
rect 40014 26126 40066 26178
rect 41694 26126 41746 26178
rect 47630 26126 47682 26178
rect 53790 26126 53842 26178
rect 55358 26126 55410 26178
rect 56702 26126 56754 26178
rect 4734 26014 4786 26066
rect 6190 26014 6242 26066
rect 7422 26014 7474 26066
rect 13358 26014 13410 26066
rect 16494 26014 16546 26066
rect 20078 26014 20130 26066
rect 24558 26014 24610 26066
rect 29150 26014 29202 26066
rect 35086 26014 35138 26066
rect 37438 26014 37490 26066
rect 45502 26014 45554 26066
rect 45838 26014 45890 26066
rect 47070 26014 47122 26066
rect 60398 26014 60450 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 16494 25678 16546 25730
rect 20302 25678 20354 25730
rect 22766 25678 22818 25730
rect 24222 25678 24274 25730
rect 26462 25678 26514 25730
rect 27582 25678 27634 25730
rect 31390 25678 31442 25730
rect 34414 25678 34466 25730
rect 34750 25678 34802 25730
rect 44830 25678 44882 25730
rect 45390 25678 45442 25730
rect 45614 25678 45666 25730
rect 46062 25678 46114 25730
rect 54574 25678 54626 25730
rect 58606 25678 58658 25730
rect 9662 25566 9714 25618
rect 10334 25566 10386 25618
rect 10670 25566 10722 25618
rect 17950 25566 18002 25618
rect 25678 25566 25730 25618
rect 28702 25566 28754 25618
rect 34862 25566 34914 25618
rect 39118 25566 39170 25618
rect 45166 25566 45218 25618
rect 46622 25566 46674 25618
rect 48750 25566 48802 25618
rect 54238 25566 54290 25618
rect 55134 25566 55186 25618
rect 58718 25566 58770 25618
rect 60958 25566 61010 25618
rect 4958 25454 5010 25506
rect 5742 25454 5794 25506
rect 6414 25454 6466 25506
rect 6750 25454 6802 25506
rect 12014 25454 12066 25506
rect 12686 25454 12738 25506
rect 13470 25454 13522 25506
rect 17054 25454 17106 25506
rect 17614 25454 17666 25506
rect 18510 25454 18562 25506
rect 18846 25454 18898 25506
rect 19630 25454 19682 25506
rect 21870 25454 21922 25506
rect 22430 25454 22482 25506
rect 23550 25454 23602 25506
rect 24782 25454 24834 25506
rect 25230 25454 25282 25506
rect 26014 25454 26066 25506
rect 26238 25454 26290 25506
rect 27022 25454 27074 25506
rect 32398 25454 32450 25506
rect 33070 25454 33122 25506
rect 34190 25454 34242 25506
rect 35422 25454 35474 25506
rect 36990 25454 37042 25506
rect 37662 25454 37714 25506
rect 38558 25454 38610 25506
rect 39566 25454 39618 25506
rect 41358 25454 41410 25506
rect 41694 25454 41746 25506
rect 42590 25454 42642 25506
rect 42926 25454 42978 25506
rect 44270 25454 44322 25506
rect 45054 25454 45106 25506
rect 49422 25454 49474 25506
rect 50878 25454 50930 25506
rect 52782 25454 52834 25506
rect 54014 25454 54066 25506
rect 54910 25454 54962 25506
rect 55806 25454 55858 25506
rect 56030 25454 56082 25506
rect 57150 25454 57202 25506
rect 58606 25454 58658 25506
rect 2382 25342 2434 25394
rect 4286 25342 4338 25394
rect 4398 25342 4450 25394
rect 5966 25342 6018 25394
rect 7534 25342 7586 25394
rect 10782 25342 10834 25394
rect 11230 25342 11282 25394
rect 11342 25342 11394 25394
rect 11678 25342 11730 25394
rect 12350 25342 12402 25394
rect 12910 25342 12962 25394
rect 14702 25342 14754 25394
rect 18286 25342 18338 25394
rect 19518 25342 19570 25394
rect 21534 25342 21586 25394
rect 22206 25342 22258 25394
rect 23886 25342 23938 25394
rect 24334 25342 24386 25394
rect 28142 25342 28194 25394
rect 33518 25342 33570 25394
rect 35086 25342 35138 25394
rect 36094 25342 36146 25394
rect 37326 25342 37378 25394
rect 38222 25342 38274 25394
rect 43150 25342 43202 25394
rect 43486 25342 43538 25394
rect 46174 25342 46226 25394
rect 50318 25342 50370 25394
rect 50542 25342 50594 25394
rect 50654 25342 50706 25394
rect 51102 25342 51154 25394
rect 52894 25342 52946 25394
rect 57262 25342 57314 25394
rect 60622 25342 60674 25394
rect 61294 25342 61346 25394
rect 61518 25342 61570 25394
rect 3726 25230 3778 25282
rect 4062 25230 4114 25282
rect 4734 25230 4786 25282
rect 5630 25230 5682 25282
rect 5854 25230 5906 25282
rect 11006 25230 11058 25282
rect 12462 25230 12514 25282
rect 13806 25230 13858 25282
rect 17166 25230 17218 25282
rect 17390 25230 17442 25282
rect 18510 25230 18562 25282
rect 20638 25230 20690 25282
rect 30046 25230 30098 25282
rect 35758 25230 35810 25282
rect 49758 25230 49810 25282
rect 49870 25230 49922 25282
rect 50094 25230 50146 25282
rect 51438 25230 51490 25282
rect 51774 25230 51826 25282
rect 53006 25230 53058 25282
rect 53230 25230 53282 25282
rect 53678 25230 53730 25282
rect 55470 25230 55522 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 6414 24894 6466 24946
rect 7534 24894 7586 24946
rect 8990 24894 9042 24946
rect 15038 24894 15090 24946
rect 16158 24894 16210 24946
rect 16606 24894 16658 24946
rect 24670 24894 24722 24946
rect 30382 24894 30434 24946
rect 30494 24894 30546 24946
rect 30606 24894 30658 24946
rect 37550 24894 37602 24946
rect 38334 24894 38386 24946
rect 41022 24894 41074 24946
rect 43150 24894 43202 24946
rect 49310 24894 49362 24946
rect 56814 24894 56866 24946
rect 57038 24894 57090 24946
rect 58830 24894 58882 24946
rect 5630 24782 5682 24834
rect 6974 24782 7026 24834
rect 8430 24782 8482 24834
rect 13134 24782 13186 24834
rect 14030 24782 14082 24834
rect 17838 24782 17890 24834
rect 18062 24782 18114 24834
rect 19630 24782 19682 24834
rect 21310 24782 21362 24834
rect 22766 24782 22818 24834
rect 25902 24782 25954 24834
rect 29150 24782 29202 24834
rect 31950 24782 32002 24834
rect 32062 24782 32114 24834
rect 33406 24782 33458 24834
rect 36318 24782 36370 24834
rect 38110 24782 38162 24834
rect 38894 24782 38946 24834
rect 40238 24782 40290 24834
rect 41918 24782 41970 24834
rect 47070 24782 47122 24834
rect 47294 24782 47346 24834
rect 48078 24782 48130 24834
rect 51326 24782 51378 24834
rect 51886 24782 51938 24834
rect 55246 24782 55298 24834
rect 57150 24782 57202 24834
rect 57822 24782 57874 24834
rect 58270 24782 58322 24834
rect 60062 24782 60114 24834
rect 3838 24670 3890 24722
rect 5070 24670 5122 24722
rect 5854 24670 5906 24722
rect 6638 24670 6690 24722
rect 7198 24670 7250 24722
rect 7870 24670 7922 24722
rect 8206 24670 8258 24722
rect 9550 24670 9602 24722
rect 13022 24670 13074 24722
rect 13358 24670 13410 24722
rect 13470 24670 13522 24722
rect 13918 24670 13970 24722
rect 15822 24670 15874 24722
rect 16830 24670 16882 24722
rect 17502 24670 17554 24722
rect 18398 24670 18450 24722
rect 18846 24670 18898 24722
rect 19182 24670 19234 24722
rect 19966 24670 20018 24722
rect 21422 24670 21474 24722
rect 22206 24670 22258 24722
rect 23662 24670 23714 24722
rect 24446 24670 24498 24722
rect 25230 24670 25282 24722
rect 25790 24670 25842 24722
rect 26798 24670 26850 24722
rect 27918 24670 27970 24722
rect 29822 24670 29874 24722
rect 30942 24670 30994 24722
rect 31390 24670 31442 24722
rect 31726 24670 31778 24722
rect 32174 24670 32226 24722
rect 37998 24670 38050 24722
rect 38670 24670 38722 24722
rect 39342 24670 39394 24722
rect 44494 24670 44546 24722
rect 45054 24670 45106 24722
rect 45502 24670 45554 24722
rect 46398 24670 46450 24722
rect 47966 24670 48018 24722
rect 48302 24670 48354 24722
rect 49534 24670 49586 24722
rect 49758 24670 49810 24722
rect 50990 24670 51042 24722
rect 51998 24670 52050 24722
rect 53006 24670 53058 24722
rect 53342 24670 53394 24722
rect 54686 24670 54738 24722
rect 55134 24670 55186 24722
rect 55470 24670 55522 24722
rect 57262 24670 57314 24722
rect 58494 24670 58546 24722
rect 59278 24670 59330 24722
rect 10334 24558 10386 24610
rect 12462 24558 12514 24610
rect 15598 24558 15650 24610
rect 17614 24558 17666 24610
rect 19070 24558 19122 24610
rect 25678 24558 25730 24610
rect 30942 24558 30994 24610
rect 31166 24558 31218 24610
rect 44718 24558 44770 24610
rect 48862 24558 48914 24610
rect 49646 24558 49698 24610
rect 52446 24558 52498 24610
rect 62190 24558 62242 24610
rect 1934 24446 1986 24498
rect 4734 24446 4786 24498
rect 6750 24446 6802 24498
rect 7646 24446 7698 24498
rect 14702 24446 14754 24498
rect 16494 24446 16546 24498
rect 18734 24446 18786 24498
rect 20414 24446 20466 24498
rect 20750 24446 20802 24498
rect 23102 24446 23154 24498
rect 23438 24446 23490 24498
rect 27134 24446 27186 24498
rect 35310 24446 35362 24498
rect 40126 24446 40178 24498
rect 46734 24446 46786 24498
rect 50206 24446 50258 24498
rect 50542 24446 50594 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 3502 24110 3554 24162
rect 6526 24110 6578 24162
rect 8094 24110 8146 24162
rect 11790 24110 11842 24162
rect 12238 24110 12290 24162
rect 12462 24110 12514 24162
rect 13694 24110 13746 24162
rect 15374 24110 15426 24162
rect 18062 24110 18114 24162
rect 26014 24110 26066 24162
rect 26350 24110 26402 24162
rect 27582 24110 27634 24162
rect 33182 24110 33234 24162
rect 35198 24110 35250 24162
rect 39230 24110 39282 24162
rect 44382 24110 44434 24162
rect 53566 24110 53618 24162
rect 60062 24110 60114 24162
rect 5070 23998 5122 24050
rect 5854 23998 5906 24050
rect 6974 23998 7026 24050
rect 10894 23998 10946 24050
rect 24334 23998 24386 24050
rect 29262 23998 29314 24050
rect 40126 23998 40178 24050
rect 44942 23998 44994 24050
rect 47854 23998 47906 24050
rect 54910 23998 54962 24050
rect 57150 23998 57202 24050
rect 4062 23886 4114 23938
rect 4286 23886 4338 23938
rect 6750 23886 6802 23938
rect 7086 23886 7138 23938
rect 7310 23886 7362 23938
rect 11902 23886 11954 23938
rect 13582 23886 13634 23938
rect 14254 23886 14306 23938
rect 15038 23886 15090 23938
rect 18398 23886 18450 23938
rect 19182 23886 19234 23938
rect 19630 23886 19682 23938
rect 19966 23886 20018 23938
rect 20078 23886 20130 23938
rect 20190 23886 20242 23938
rect 24110 23886 24162 23938
rect 24446 23886 24498 23938
rect 24670 23886 24722 23938
rect 25678 23886 25730 23938
rect 26126 23886 26178 23938
rect 27022 23886 27074 23938
rect 28366 23886 28418 23938
rect 29822 23886 29874 23938
rect 31614 23886 31666 23938
rect 32062 23886 32114 23938
rect 32174 23886 32226 23938
rect 33518 23886 33570 23938
rect 34190 23886 34242 23938
rect 39006 23886 39058 23938
rect 39342 23886 39394 23938
rect 39790 23886 39842 23938
rect 41582 23886 41634 23938
rect 45950 23886 46002 23938
rect 46734 23886 46786 23938
rect 47518 23886 47570 23938
rect 48638 23886 48690 23938
rect 49422 23886 49474 23938
rect 50654 23886 50706 23938
rect 51102 23886 51154 23938
rect 51438 23886 51490 23938
rect 51662 23886 51714 23938
rect 52894 23886 52946 23938
rect 54798 23886 54850 23938
rect 57038 23886 57090 23938
rect 60958 23886 61010 23938
rect 2382 23774 2434 23826
rect 6302 23774 6354 23826
rect 7758 23774 7810 23826
rect 7982 23774 8034 23826
rect 9774 23774 9826 23826
rect 11118 23774 11170 23826
rect 11454 23774 11506 23826
rect 11678 23774 11730 23826
rect 14030 23774 14082 23826
rect 17278 23774 17330 23826
rect 18958 23774 19010 23826
rect 21870 23774 21922 23826
rect 24894 23774 24946 23826
rect 25454 23774 25506 23826
rect 25902 23774 25954 23826
rect 27918 23774 27970 23826
rect 28478 23774 28530 23826
rect 29486 23774 29538 23826
rect 31838 23774 31890 23826
rect 34302 23774 34354 23826
rect 35422 23774 35474 23826
rect 35758 23774 35810 23826
rect 37326 23774 37378 23826
rect 42590 23774 42642 23826
rect 45278 23774 45330 23826
rect 46846 23774 46898 23826
rect 47630 23774 47682 23826
rect 49310 23774 49362 23826
rect 49982 23774 50034 23826
rect 50878 23774 50930 23826
rect 53454 23774 53506 23826
rect 56590 23774 56642 23826
rect 56702 23774 56754 23826
rect 58158 23774 58210 23826
rect 60622 23774 60674 23826
rect 61182 23774 61234 23826
rect 61630 23774 61682 23826
rect 4622 23662 4674 23714
rect 6414 23662 6466 23714
rect 8766 23662 8818 23714
rect 9214 23662 9266 23714
rect 9438 23662 9490 23714
rect 9662 23662 9714 23714
rect 10334 23662 10386 23714
rect 11230 23662 11282 23714
rect 14142 23662 14194 23714
rect 14814 23662 14866 23714
rect 19742 23662 19794 23714
rect 23102 23662 23154 23714
rect 28702 23662 28754 23714
rect 29150 23662 29202 23714
rect 29374 23662 29426 23714
rect 30382 23662 30434 23714
rect 30606 23662 30658 23714
rect 30718 23662 30770 23714
rect 30830 23662 30882 23714
rect 31390 23662 31442 23714
rect 32398 23662 32450 23714
rect 34862 23662 34914 23714
rect 36990 23662 37042 23714
rect 41694 23662 41746 23714
rect 41918 23662 41970 23714
rect 44830 23662 44882 23714
rect 45054 23662 45106 23714
rect 45950 23662 46002 23714
rect 51326 23662 51378 23714
rect 56366 23662 56418 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 2046 23326 2098 23378
rect 6862 23326 6914 23378
rect 9774 23326 9826 23378
rect 17614 23326 17666 23378
rect 18174 23326 18226 23378
rect 19406 23326 19458 23378
rect 25230 23326 25282 23378
rect 29934 23326 29986 23378
rect 34302 23326 34354 23378
rect 35422 23326 35474 23378
rect 36766 23326 36818 23378
rect 37438 23326 37490 23378
rect 40126 23326 40178 23378
rect 40238 23326 40290 23378
rect 46286 23326 46338 23378
rect 47518 23326 47570 23378
rect 56590 23326 56642 23378
rect 1710 23214 1762 23266
rect 2606 23214 2658 23266
rect 11566 23214 11618 23266
rect 14814 23214 14866 23266
rect 15374 23214 15426 23266
rect 16046 23214 16098 23266
rect 16830 23214 16882 23266
rect 17838 23214 17890 23266
rect 20526 23214 20578 23266
rect 23438 23214 23490 23266
rect 23662 23214 23714 23266
rect 31726 23214 31778 23266
rect 33182 23214 33234 23266
rect 35870 23214 35922 23266
rect 36990 23214 37042 23266
rect 37550 23214 37602 23266
rect 39118 23214 39170 23266
rect 40014 23214 40066 23266
rect 44606 23214 44658 23266
rect 46622 23214 46674 23266
rect 47182 23214 47234 23266
rect 47406 23214 47458 23266
rect 49646 23214 49698 23266
rect 53566 23214 53618 23266
rect 60958 23214 61010 23266
rect 2830 23102 2882 23154
rect 3502 23102 3554 23154
rect 5966 23102 6018 23154
rect 6190 23102 6242 23154
rect 7086 23102 7138 23154
rect 7534 23102 7586 23154
rect 8430 23102 8482 23154
rect 10110 23102 10162 23154
rect 14366 23102 14418 23154
rect 15150 23102 15202 23154
rect 16158 23102 16210 23154
rect 16606 23102 16658 23154
rect 18286 23102 18338 23154
rect 18510 23102 18562 23154
rect 18958 23102 19010 23154
rect 19630 23102 19682 23154
rect 21086 23102 21138 23154
rect 22430 23102 22482 23154
rect 22990 23102 23042 23154
rect 23214 23102 23266 23154
rect 24558 23102 24610 23154
rect 25790 23102 25842 23154
rect 27582 23102 27634 23154
rect 27806 23102 27858 23154
rect 28478 23102 28530 23154
rect 29598 23102 29650 23154
rect 36094 23102 36146 23154
rect 36654 23102 36706 23154
rect 38334 23102 38386 23154
rect 39006 23102 39058 23154
rect 39566 23102 39618 23154
rect 40350 23102 40402 23154
rect 41806 23102 41858 23154
rect 42366 23102 42418 23154
rect 43038 23102 43090 23154
rect 44270 23102 44322 23154
rect 44942 23102 44994 23154
rect 45726 23102 45778 23154
rect 46846 23102 46898 23154
rect 47854 23102 47906 23154
rect 48750 23102 48802 23154
rect 49870 23102 49922 23154
rect 51550 23102 51602 23154
rect 52222 23102 52274 23154
rect 52894 23102 52946 23154
rect 54574 23102 54626 23154
rect 56926 23102 56978 23154
rect 58606 23102 58658 23154
rect 59054 23102 59106 23154
rect 59950 23102 60002 23154
rect 3166 22990 3218 23042
rect 3838 22990 3890 23042
rect 8094 22990 8146 23042
rect 8990 22990 9042 23042
rect 10558 22990 10610 23042
rect 14702 22990 14754 23042
rect 21646 22990 21698 23042
rect 24446 22990 24498 23042
rect 45950 22990 46002 23042
rect 48190 22990 48242 23042
rect 54798 22990 54850 23042
rect 57150 22990 57202 23042
rect 57822 22990 57874 23042
rect 13470 22878 13522 22930
rect 16046 22878 16098 22930
rect 17502 22878 17554 22930
rect 19070 22878 19122 22930
rect 29262 22878 29314 22930
rect 33070 22878 33122 22930
rect 37998 22878 38050 22930
rect 41022 22878 41074 22930
rect 52782 22878 52834 22930
rect 62078 22878 62130 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 22318 22542 22370 22594
rect 24782 22542 24834 22594
rect 25678 22542 25730 22594
rect 32622 22542 32674 22594
rect 39006 22542 39058 22594
rect 49982 22542 50034 22594
rect 51102 22542 51154 22594
rect 60622 22542 60674 22594
rect 60958 22542 61010 22594
rect 4622 22430 4674 22482
rect 9102 22430 9154 22482
rect 9550 22430 9602 22482
rect 10670 22430 10722 22482
rect 12462 22430 12514 22482
rect 13582 22430 13634 22482
rect 14030 22430 14082 22482
rect 14926 22430 14978 22482
rect 18398 22430 18450 22482
rect 20526 22430 20578 22482
rect 21422 22430 21474 22482
rect 29374 22430 29426 22482
rect 39790 22430 39842 22482
rect 45278 22430 45330 22482
rect 45838 22430 45890 22482
rect 47966 22430 48018 22482
rect 54238 22430 54290 22482
rect 5630 22318 5682 22370
rect 6974 22318 7026 22370
rect 8654 22318 8706 22370
rect 9774 22318 9826 22370
rect 10222 22318 10274 22370
rect 11006 22318 11058 22370
rect 11790 22318 11842 22370
rect 13022 22318 13074 22370
rect 13918 22318 13970 22370
rect 14142 22318 14194 22370
rect 14478 22318 14530 22370
rect 15038 22318 15090 22370
rect 15374 22318 15426 22370
rect 15710 22318 15762 22370
rect 17614 22318 17666 22370
rect 21870 22318 21922 22370
rect 22430 22318 22482 22370
rect 25230 22318 25282 22370
rect 26462 22318 26514 22370
rect 27358 22318 27410 22370
rect 30046 22318 30098 22370
rect 30494 22318 30546 22370
rect 31502 22318 31554 22370
rect 32062 22318 32114 22370
rect 32398 22318 32450 22370
rect 33518 22318 33570 22370
rect 33854 22318 33906 22370
rect 35198 22318 35250 22370
rect 35870 22318 35922 22370
rect 36318 22318 36370 22370
rect 39454 22318 39506 22370
rect 40686 22318 40738 22370
rect 41694 22318 41746 22370
rect 44830 22318 44882 22370
rect 45166 22318 45218 22370
rect 45390 22318 45442 22370
rect 47630 22318 47682 22370
rect 47854 22318 47906 22370
rect 49310 22318 49362 22370
rect 49758 22318 49810 22370
rect 50542 22318 50594 22370
rect 52670 22318 52722 22370
rect 53454 22318 53506 22370
rect 53790 22318 53842 22370
rect 54350 22318 54402 22370
rect 57486 22318 57538 22370
rect 58158 22318 58210 22370
rect 3502 22206 3554 22258
rect 6414 22206 6466 22258
rect 7534 22206 7586 22258
rect 9550 22206 9602 22258
rect 10894 22206 10946 22258
rect 12350 22206 12402 22258
rect 14814 22206 14866 22258
rect 17278 22206 17330 22258
rect 22318 22206 22370 22258
rect 28030 22206 28082 22258
rect 31838 22206 31890 22258
rect 32174 22206 32226 22258
rect 33070 22206 33122 22258
rect 33294 22206 33346 22258
rect 34526 22206 34578 22258
rect 37550 22206 37602 22258
rect 40910 22206 40962 22258
rect 42702 22206 42754 22258
rect 48862 22206 48914 22258
rect 51550 22206 51602 22258
rect 53118 22206 53170 22258
rect 54014 22206 54066 22258
rect 55134 22206 55186 22258
rect 57262 22206 57314 22258
rect 59390 22206 59442 22258
rect 61294 22206 61346 22258
rect 61518 22206 61570 22258
rect 1710 22094 1762 22146
rect 5070 22094 5122 22146
rect 12014 22094 12066 22146
rect 12574 22094 12626 22146
rect 15822 22094 15874 22146
rect 16942 22094 16994 22146
rect 23438 22094 23490 22146
rect 33854 22094 33906 22146
rect 34190 22094 34242 22146
rect 34862 22094 34914 22146
rect 35982 22094 36034 22146
rect 36430 22094 36482 22146
rect 41582 22094 41634 22146
rect 44158 22094 44210 22146
rect 52110 22094 52162 22146
rect 53230 22094 53282 22146
rect 53342 22094 53394 22146
rect 57038 22094 57090 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 2382 21758 2434 21810
rect 4622 21758 4674 21810
rect 4846 21758 4898 21810
rect 7646 21758 7698 21810
rect 11342 21758 11394 21810
rect 14926 21758 14978 21810
rect 17726 21758 17778 21810
rect 19518 21758 19570 21810
rect 19630 21758 19682 21810
rect 20302 21758 20354 21810
rect 22654 21758 22706 21810
rect 23886 21758 23938 21810
rect 29710 21758 29762 21810
rect 31054 21758 31106 21810
rect 33294 21758 33346 21810
rect 33966 21758 34018 21810
rect 40014 21758 40066 21810
rect 41582 21758 41634 21810
rect 41918 21758 41970 21810
rect 42142 21758 42194 21810
rect 43262 21758 43314 21810
rect 44494 21758 44546 21810
rect 45390 21758 45442 21810
rect 45838 21758 45890 21810
rect 46622 21758 46674 21810
rect 55358 21758 55410 21810
rect 55694 21758 55746 21810
rect 61518 21758 61570 21810
rect 3502 21646 3554 21698
rect 4398 21646 4450 21698
rect 5182 21646 5234 21698
rect 8318 21646 8370 21698
rect 8766 21646 8818 21698
rect 11790 21646 11842 21698
rect 15598 21646 15650 21698
rect 17614 21646 17666 21698
rect 18398 21646 18450 21698
rect 19406 21646 19458 21698
rect 19966 21646 20018 21698
rect 20974 21646 21026 21698
rect 21310 21646 21362 21698
rect 21646 21646 21698 21698
rect 23550 21646 23602 21698
rect 23662 21646 23714 21698
rect 26462 21646 26514 21698
rect 28030 21646 28082 21698
rect 30270 21646 30322 21698
rect 31614 21646 31666 21698
rect 32174 21646 32226 21698
rect 33630 21646 33682 21698
rect 39678 21646 39730 21698
rect 42366 21646 42418 21698
rect 43822 21646 43874 21698
rect 44158 21646 44210 21698
rect 47742 21646 47794 21698
rect 48750 21646 48802 21698
rect 48974 21646 49026 21698
rect 49086 21646 49138 21698
rect 49310 21646 49362 21698
rect 51326 21646 51378 21698
rect 58382 21646 58434 21698
rect 59614 21646 59666 21698
rect 5406 21534 5458 21586
rect 6190 21534 6242 21586
rect 6638 21534 6690 21586
rect 11118 21534 11170 21586
rect 12014 21534 12066 21586
rect 13582 21534 13634 21586
rect 13806 21534 13858 21586
rect 14478 21534 14530 21586
rect 14702 21534 14754 21586
rect 15486 21534 15538 21586
rect 17390 21534 17442 21586
rect 18846 21534 18898 21586
rect 19182 21534 19234 21586
rect 20638 21534 20690 21586
rect 22318 21534 22370 21586
rect 22878 21534 22930 21586
rect 23326 21534 23378 21586
rect 24558 21534 24610 21586
rect 25342 21534 25394 21586
rect 33070 21534 33122 21586
rect 33294 21534 33346 21586
rect 34526 21534 34578 21586
rect 34974 21534 35026 21586
rect 35758 21534 35810 21586
rect 38670 21534 38722 21586
rect 39118 21534 39170 21586
rect 40238 21534 40290 21586
rect 41022 21534 41074 21586
rect 42030 21534 42082 21586
rect 43598 21534 43650 21586
rect 44830 21534 44882 21586
rect 45054 21534 45106 21586
rect 45726 21534 45778 21586
rect 46958 21534 47010 21586
rect 47630 21534 47682 21586
rect 49870 21534 49922 21586
rect 53006 21534 53058 21586
rect 54686 21534 54738 21586
rect 55022 21534 55074 21586
rect 55246 21534 55298 21586
rect 55918 21534 55970 21586
rect 57262 21534 57314 21586
rect 58270 21534 58322 21586
rect 59054 21534 59106 21586
rect 59278 21534 59330 21586
rect 4734 21422 4786 21474
rect 6078 21422 6130 21474
rect 9886 21422 9938 21474
rect 10782 21422 10834 21474
rect 12574 21422 12626 21474
rect 14142 21422 14194 21474
rect 14590 21422 14642 21474
rect 21982 21422 22034 21474
rect 22766 21422 22818 21474
rect 24222 21422 24274 21474
rect 29262 21422 29314 21474
rect 30046 21422 30098 21474
rect 34302 21422 34354 21474
rect 37886 21422 37938 21474
rect 38222 21422 38274 21474
rect 42926 21422 42978 21474
rect 48862 21422 48914 21474
rect 49982 21422 50034 21474
rect 53454 21422 53506 21474
rect 54014 21422 54066 21474
rect 57598 21422 57650 21474
rect 58382 21422 58434 21474
rect 59502 21422 59554 21474
rect 7982 21310 8034 21362
rect 10222 21310 10274 21362
rect 10558 21310 10610 21362
rect 12798 21310 12850 21362
rect 13134 21310 13186 21362
rect 16270 21310 16322 21362
rect 16606 21310 16658 21362
rect 31390 21310 31442 21362
rect 41246 21310 41298 21362
rect 52558 21310 52610 21362
rect 54126 21310 54178 21362
rect 54462 21310 54514 21362
rect 59054 21310 59106 21362
rect 60174 21310 60226 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 3278 20974 3330 21026
rect 4174 20974 4226 21026
rect 4510 20974 4562 21026
rect 5630 20974 5682 21026
rect 12014 20974 12066 21026
rect 17390 20974 17442 21026
rect 27134 20974 27186 21026
rect 27470 20974 27522 21026
rect 29374 20974 29426 21026
rect 48302 20974 48354 21026
rect 58606 20974 58658 21026
rect 60510 20974 60562 21026
rect 61630 20974 61682 21026
rect 61966 20974 62018 21026
rect 5742 20862 5794 20914
rect 7758 20862 7810 20914
rect 9214 20862 9266 20914
rect 12462 20862 12514 20914
rect 14030 20862 14082 20914
rect 15598 20862 15650 20914
rect 17838 20862 17890 20914
rect 21310 20862 21362 20914
rect 22542 20862 22594 20914
rect 24670 20862 24722 20914
rect 29934 20862 29986 20914
rect 31726 20862 31778 20914
rect 31950 20862 32002 20914
rect 33070 20862 33122 20914
rect 35198 20862 35250 20914
rect 36318 20862 36370 20914
rect 38446 20862 38498 20914
rect 39454 20862 39506 20914
rect 49534 20862 49586 20914
rect 53118 20862 53170 20914
rect 54238 20862 54290 20914
rect 62190 20862 62242 20914
rect 1822 20750 1874 20802
rect 2718 20750 2770 20802
rect 3054 20750 3106 20802
rect 3950 20750 4002 20802
rect 4846 20750 4898 20802
rect 6974 20750 7026 20802
rect 7870 20750 7922 20802
rect 8094 20750 8146 20802
rect 8990 20750 9042 20802
rect 9550 20750 9602 20802
rect 13694 20750 13746 20802
rect 14590 20750 14642 20802
rect 17278 20750 17330 20802
rect 17950 20750 18002 20802
rect 20078 20750 20130 20802
rect 20414 20750 20466 20802
rect 20638 20750 20690 20802
rect 21422 20750 21474 20802
rect 21870 20750 21922 20802
rect 24894 20750 24946 20802
rect 25678 20750 25730 20802
rect 27918 20750 27970 20802
rect 29262 20750 29314 20802
rect 31054 20750 31106 20802
rect 31614 20750 31666 20802
rect 32398 20750 32450 20802
rect 36206 20750 36258 20802
rect 37102 20750 37154 20802
rect 38110 20750 38162 20802
rect 39006 20750 39058 20802
rect 40126 20750 40178 20802
rect 40574 20750 40626 20802
rect 40910 20750 40962 20802
rect 43038 20750 43090 20802
rect 45166 20750 45218 20802
rect 46286 20750 46338 20802
rect 47630 20750 47682 20802
rect 52670 20750 52722 20802
rect 53902 20750 53954 20802
rect 54014 20750 54066 20802
rect 54462 20750 54514 20802
rect 55694 20750 55746 20802
rect 56142 20750 56194 20802
rect 56366 20750 56418 20802
rect 56590 20750 56642 20802
rect 58382 20750 58434 20802
rect 58830 20750 58882 20802
rect 59054 20750 59106 20802
rect 59166 20750 59218 20802
rect 59838 20750 59890 20802
rect 60734 20750 60786 20802
rect 6302 20638 6354 20690
rect 6638 20638 6690 20690
rect 8318 20638 8370 20690
rect 9438 20638 9490 20690
rect 14478 20638 14530 20690
rect 15150 20638 15202 20690
rect 15374 20638 15426 20690
rect 15486 20638 15538 20690
rect 15710 20638 15762 20690
rect 16606 20638 16658 20690
rect 25118 20638 25170 20690
rect 25230 20638 25282 20690
rect 26126 20638 26178 20690
rect 26574 20638 26626 20690
rect 28254 20638 28306 20690
rect 29822 20638 29874 20690
rect 30158 20638 30210 20690
rect 30382 20638 30434 20690
rect 30718 20638 30770 20690
rect 31278 20638 31330 20690
rect 35870 20638 35922 20690
rect 40798 20638 40850 20690
rect 41358 20638 41410 20690
rect 42254 20638 42306 20690
rect 42814 20638 42866 20690
rect 47518 20638 47570 20690
rect 50990 20638 51042 20690
rect 56254 20638 56306 20690
rect 59502 20638 59554 20690
rect 1934 20526 1986 20578
rect 2158 20526 2210 20578
rect 2606 20526 2658 20578
rect 3614 20526 3666 20578
rect 4958 20526 5010 20578
rect 5182 20526 5234 20578
rect 7310 20526 7362 20578
rect 8542 20526 8594 20578
rect 10670 20526 10722 20578
rect 12574 20526 12626 20578
rect 20526 20526 20578 20578
rect 25902 20526 25954 20578
rect 30942 20526 30994 20578
rect 35534 20526 35586 20578
rect 35758 20526 35810 20578
rect 37214 20526 37266 20578
rect 40350 20526 40402 20578
rect 41694 20526 41746 20578
rect 43374 20526 43426 20578
rect 43822 20526 43874 20578
rect 44158 20526 44210 20578
rect 48750 20526 48802 20578
rect 49086 20526 49138 20578
rect 51998 20526 52050 20578
rect 60958 20526 61010 20578
rect 61070 20526 61122 20578
rect 61182 20526 61234 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 43038 20190 43090 20242
rect 44158 20190 44210 20242
rect 50542 20190 50594 20242
rect 57598 20190 57650 20242
rect 2494 20078 2546 20130
rect 5182 20078 5234 20130
rect 5294 20078 5346 20130
rect 5518 20078 5570 20130
rect 6078 20078 6130 20130
rect 7534 20078 7586 20130
rect 7758 20078 7810 20130
rect 8430 20078 8482 20130
rect 8766 20078 8818 20130
rect 8990 20078 9042 20130
rect 11230 20078 11282 20130
rect 11790 20078 11842 20130
rect 22094 20078 22146 20130
rect 25902 20078 25954 20130
rect 29710 20078 29762 20130
rect 30494 20078 30546 20130
rect 30718 20078 30770 20130
rect 31054 20078 31106 20130
rect 31726 20078 31778 20130
rect 34862 20078 34914 20130
rect 39902 20078 39954 20130
rect 41806 20078 41858 20130
rect 45950 20078 46002 20130
rect 47854 20078 47906 20130
rect 47966 20078 48018 20130
rect 48862 20078 48914 20130
rect 51662 20078 51714 20130
rect 52222 20078 52274 20130
rect 53902 20078 53954 20130
rect 54350 20078 54402 20130
rect 54574 20078 54626 20130
rect 57710 20078 57762 20130
rect 58942 20078 58994 20130
rect 61518 20078 61570 20130
rect 1710 19966 1762 20018
rect 5742 19966 5794 20018
rect 6302 19966 6354 20018
rect 7198 19966 7250 20018
rect 8542 19966 8594 20018
rect 9550 19966 9602 20018
rect 9774 19966 9826 20018
rect 10670 19966 10722 20018
rect 12014 19966 12066 20018
rect 12686 19966 12738 20018
rect 13470 19966 13522 20018
rect 14702 19966 14754 20018
rect 15374 19966 15426 20018
rect 16494 19966 16546 20018
rect 17390 19966 17442 20018
rect 20302 19966 20354 20018
rect 20526 19966 20578 20018
rect 21422 19966 21474 20018
rect 24782 19966 24834 20018
rect 25454 19966 25506 20018
rect 26350 19966 26402 20018
rect 28254 19966 28306 20018
rect 29822 19966 29874 20018
rect 30382 19966 30434 20018
rect 30942 19966 30994 20018
rect 31950 19966 32002 20018
rect 32510 19966 32562 20018
rect 33630 19966 33682 20018
rect 34190 19966 34242 20018
rect 36094 19966 36146 20018
rect 37326 19966 37378 20018
rect 37662 19966 37714 20018
rect 39118 19966 39170 20018
rect 39454 19966 39506 20018
rect 45502 19966 45554 20018
rect 47070 19966 47122 20018
rect 48750 19966 48802 20018
rect 48974 19966 49026 20018
rect 49310 19966 49362 20018
rect 53678 19966 53730 20018
rect 55022 19966 55074 20018
rect 55918 19966 55970 20018
rect 57038 19966 57090 20018
rect 58158 19966 58210 20018
rect 61406 19966 61458 20018
rect 61630 19966 61682 20018
rect 61966 19966 62018 20018
rect 4622 19854 4674 19906
rect 10110 19854 10162 19906
rect 12238 19854 12290 19906
rect 12350 19854 12402 19906
rect 18062 19854 18114 19906
rect 20078 19854 20130 19906
rect 24222 19854 24274 19906
rect 25566 19854 25618 19906
rect 26238 19854 26290 19906
rect 27246 19854 27298 19906
rect 27694 19854 27746 19906
rect 33518 19854 33570 19906
rect 46398 19854 46450 19906
rect 46846 19854 46898 19906
rect 54462 19854 54514 19906
rect 55470 19854 55522 19906
rect 56590 19854 56642 19906
rect 61070 19854 61122 19906
rect 16606 19742 16658 19794
rect 27358 19742 27410 19794
rect 28702 19742 28754 19794
rect 29038 19742 29090 19794
rect 34078 19742 34130 19794
rect 47406 19742 47458 19794
rect 47854 19742 47906 19794
rect 52110 19742 52162 19794
rect 52782 19742 52834 19794
rect 53118 19742 53170 19794
rect 57486 19742 57538 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 21422 19406 21474 19458
rect 21758 19406 21810 19458
rect 26686 19406 26738 19458
rect 42030 19406 42082 19458
rect 45054 19406 45106 19458
rect 52782 19406 52834 19458
rect 56814 19406 56866 19458
rect 59838 19406 59890 19458
rect 60510 19406 60562 19458
rect 5966 19294 6018 19346
rect 14142 19294 14194 19346
rect 16942 19294 16994 19346
rect 19518 19294 19570 19346
rect 23214 19294 23266 19346
rect 29374 19294 29426 19346
rect 30158 19294 30210 19346
rect 36206 19294 36258 19346
rect 42254 19294 42306 19346
rect 47182 19294 47234 19346
rect 50542 19294 50594 19346
rect 51662 19294 51714 19346
rect 53230 19294 53282 19346
rect 4734 19182 4786 19234
rect 6414 19182 6466 19234
rect 6638 19182 6690 19234
rect 6974 19182 7026 19234
rect 7310 19182 7362 19234
rect 7758 19182 7810 19234
rect 9662 19182 9714 19234
rect 9886 19182 9938 19234
rect 10334 19182 10386 19234
rect 11790 19182 11842 19234
rect 12350 19182 12402 19234
rect 13918 19182 13970 19234
rect 14590 19182 14642 19234
rect 15710 19182 15762 19234
rect 16830 19182 16882 19234
rect 19630 19182 19682 19234
rect 20414 19182 20466 19234
rect 24222 19182 24274 19234
rect 25566 19182 25618 19234
rect 26686 19182 26738 19234
rect 27022 19182 27074 19234
rect 27134 19182 27186 19234
rect 29598 19182 29650 19234
rect 33070 19182 33122 19234
rect 34190 19182 34242 19234
rect 34974 19182 35026 19234
rect 35758 19182 35810 19234
rect 36094 19182 36146 19234
rect 42366 19182 42418 19234
rect 43038 19182 43090 19234
rect 44270 19182 44322 19234
rect 44830 19182 44882 19234
rect 45950 19182 46002 19234
rect 46398 19182 46450 19234
rect 47742 19182 47794 19234
rect 51214 19182 51266 19234
rect 52222 19182 52274 19234
rect 52558 19182 52610 19234
rect 53566 19182 53618 19234
rect 54350 19182 54402 19234
rect 55694 19182 55746 19234
rect 56254 19182 56306 19234
rect 56478 19182 56530 19234
rect 58158 19182 58210 19234
rect 58494 19182 58546 19234
rect 59502 19182 59554 19234
rect 60734 19182 60786 19234
rect 2942 19070 2994 19122
rect 5630 19070 5682 19122
rect 11118 19070 11170 19122
rect 11454 19070 11506 19122
rect 12574 19070 12626 19122
rect 14254 19070 14306 19122
rect 14926 19070 14978 19122
rect 15374 19070 15426 19122
rect 15486 19070 15538 19122
rect 16494 19070 16546 19122
rect 21982 19070 22034 19122
rect 22318 19070 22370 19122
rect 23774 19070 23826 19122
rect 24558 19070 24610 19122
rect 24670 19070 24722 19122
rect 31166 19070 31218 19122
rect 33294 19070 33346 19122
rect 33854 19070 33906 19122
rect 34750 19070 34802 19122
rect 38558 19070 38610 19122
rect 40238 19070 40290 19122
rect 42702 19070 42754 19122
rect 43710 19070 43762 19122
rect 44046 19070 44098 19122
rect 45390 19070 45442 19122
rect 45502 19070 45554 19122
rect 45614 19070 45666 19122
rect 46846 19070 46898 19122
rect 48414 19070 48466 19122
rect 50878 19070 50930 19122
rect 58606 19070 58658 19122
rect 59726 19070 59778 19122
rect 61406 19070 61458 19122
rect 61854 19070 61906 19122
rect 2046 18958 2098 19010
rect 6750 18958 6802 19010
rect 11902 18958 11954 19010
rect 15934 18958 15986 19010
rect 23662 18958 23714 19010
rect 24782 18958 24834 19010
rect 24894 18958 24946 19010
rect 32510 18958 32562 19010
rect 37102 18958 37154 19010
rect 42814 18958 42866 19010
rect 43934 18958 43986 19010
rect 47070 18958 47122 19010
rect 51550 18958 51602 19010
rect 51774 18958 51826 19010
rect 59838 18958 59890 19010
rect 61518 18958 61570 19010
rect 62190 18958 62242 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 8430 18622 8482 18674
rect 10334 18622 10386 18674
rect 13358 18622 13410 18674
rect 13582 18622 13634 18674
rect 24110 18622 24162 18674
rect 24334 18622 24386 18674
rect 33182 18622 33234 18674
rect 36878 18622 36930 18674
rect 41022 18622 41074 18674
rect 50206 18622 50258 18674
rect 53790 18622 53842 18674
rect 57710 18622 57762 18674
rect 60846 18622 60898 18674
rect 4846 18510 4898 18562
rect 8654 18510 8706 18562
rect 10558 18510 10610 18562
rect 11342 18510 11394 18562
rect 13918 18510 13970 18562
rect 16046 18510 16098 18562
rect 16606 18510 16658 18562
rect 22430 18510 22482 18562
rect 25790 18510 25842 18562
rect 33742 18510 33794 18562
rect 35758 18510 35810 18562
rect 42030 18510 42082 18562
rect 44942 18510 44994 18562
rect 46062 18510 46114 18562
rect 49422 18510 49474 18562
rect 49534 18510 49586 18562
rect 50990 18510 51042 18562
rect 51326 18510 51378 18562
rect 53678 18510 53730 18562
rect 54014 18510 54066 18562
rect 57038 18510 57090 18562
rect 59950 18510 60002 18562
rect 61854 18510 61906 18562
rect 2718 18398 2770 18450
rect 3054 18398 3106 18450
rect 3614 18398 3666 18450
rect 6526 18398 6578 18450
rect 7534 18398 7586 18450
rect 7870 18398 7922 18450
rect 8206 18398 8258 18450
rect 9998 18398 10050 18450
rect 13470 18398 13522 18450
rect 13806 18398 13858 18450
rect 15374 18398 15426 18450
rect 16718 18398 16770 18450
rect 18062 18398 18114 18450
rect 18958 18398 19010 18450
rect 19854 18398 19906 18450
rect 20190 18398 20242 18450
rect 20526 18398 20578 18450
rect 22206 18398 22258 18450
rect 22766 18398 22818 18450
rect 24222 18398 24274 18450
rect 24670 18398 24722 18450
rect 28254 18398 28306 18450
rect 28366 18398 28418 18450
rect 30494 18398 30546 18450
rect 30718 18398 30770 18450
rect 32398 18398 32450 18450
rect 33070 18398 33122 18450
rect 33630 18398 33682 18450
rect 35086 18398 35138 18450
rect 36206 18398 36258 18450
rect 37438 18398 37490 18450
rect 42142 18398 42194 18450
rect 42702 18398 42754 18450
rect 42814 18398 42866 18450
rect 43150 18398 43202 18450
rect 44046 18398 44098 18450
rect 45166 18398 45218 18450
rect 46286 18398 46338 18450
rect 47630 18398 47682 18450
rect 48750 18398 48802 18450
rect 49758 18398 49810 18450
rect 49982 18398 50034 18450
rect 50654 18398 50706 18450
rect 51998 18398 52050 18450
rect 52334 18398 52386 18450
rect 53118 18398 53170 18450
rect 53342 18398 53394 18450
rect 54126 18398 54178 18450
rect 54910 18398 54962 18450
rect 56030 18398 56082 18450
rect 57374 18398 57426 18450
rect 57934 18398 57986 18450
rect 61182 18398 61234 18450
rect 62078 18398 62130 18450
rect 2270 18286 2322 18338
rect 3950 18286 4002 18338
rect 8318 18286 8370 18338
rect 9774 18286 9826 18338
rect 10446 18286 10498 18338
rect 15038 18286 15090 18338
rect 16942 18286 16994 18338
rect 17614 18286 17666 18338
rect 23326 18286 23378 18338
rect 23886 18286 23938 18338
rect 27022 18286 27074 18338
rect 28702 18286 28754 18338
rect 31950 18286 32002 18338
rect 35422 18286 35474 18338
rect 38222 18286 38274 18338
rect 40350 18286 40402 18338
rect 43038 18286 43090 18338
rect 43598 18286 43650 18338
rect 46398 18286 46450 18338
rect 48862 18286 48914 18338
rect 50094 18286 50146 18338
rect 13134 18174 13186 18226
rect 18510 18174 18562 18226
rect 35086 18174 35138 18226
rect 41358 18174 41410 18226
rect 44382 18174 44434 18226
rect 52222 18174 52274 18226
rect 54350 18174 54402 18226
rect 55806 18174 55858 18226
rect 58494 18174 58546 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 12014 17838 12066 17890
rect 14702 17838 14754 17890
rect 15262 17838 15314 17890
rect 15822 17838 15874 17890
rect 18734 17838 18786 17890
rect 25678 17838 25730 17890
rect 33966 17838 34018 17890
rect 39566 17838 39618 17890
rect 40014 17838 40066 17890
rect 41470 17838 41522 17890
rect 44830 17838 44882 17890
rect 45278 17838 45330 17890
rect 51774 17838 51826 17890
rect 55806 17838 55858 17890
rect 60622 17838 60674 17890
rect 2046 17726 2098 17778
rect 5966 17726 6018 17778
rect 6862 17726 6914 17778
rect 11342 17726 11394 17778
rect 14366 17726 14418 17778
rect 19630 17726 19682 17778
rect 20078 17726 20130 17778
rect 24894 17726 24946 17778
rect 29598 17726 29650 17778
rect 30382 17726 30434 17778
rect 30718 17726 30770 17778
rect 35758 17726 35810 17778
rect 37886 17726 37938 17778
rect 44942 17726 44994 17778
rect 48302 17726 48354 17778
rect 50318 17726 50370 17778
rect 52558 17726 52610 17778
rect 56814 17726 56866 17778
rect 7310 17614 7362 17666
rect 7982 17614 8034 17666
rect 9662 17614 9714 17666
rect 9886 17614 9938 17666
rect 10110 17614 10162 17666
rect 12686 17614 12738 17666
rect 18174 17614 18226 17666
rect 19070 17614 19122 17666
rect 19294 17614 19346 17666
rect 20190 17614 20242 17666
rect 21982 17614 22034 17666
rect 26350 17614 26402 17666
rect 26686 17614 26738 17666
rect 27134 17614 27186 17666
rect 28478 17614 28530 17666
rect 29150 17614 29202 17666
rect 30270 17614 30322 17666
rect 30830 17614 30882 17666
rect 34974 17614 35026 17666
rect 36990 17614 37042 17666
rect 37550 17614 37602 17666
rect 38222 17614 38274 17666
rect 40238 17614 40290 17666
rect 41134 17614 41186 17666
rect 41358 17614 41410 17666
rect 42814 17614 42866 17666
rect 43822 17614 43874 17666
rect 47854 17614 47906 17666
rect 48190 17614 48242 17666
rect 49086 17614 49138 17666
rect 49422 17614 49474 17666
rect 50654 17614 50706 17666
rect 51662 17614 51714 17666
rect 51886 17614 51938 17666
rect 53790 17614 53842 17666
rect 54238 17614 54290 17666
rect 54686 17614 54738 17666
rect 55022 17614 55074 17666
rect 56366 17614 56418 17666
rect 57038 17614 57090 17666
rect 60510 17614 60562 17666
rect 60734 17614 60786 17666
rect 61630 17614 61682 17666
rect 61854 17614 61906 17666
rect 62190 17614 62242 17666
rect 3838 17502 3890 17554
rect 12798 17502 12850 17554
rect 13582 17502 13634 17554
rect 14142 17502 14194 17554
rect 15262 17502 15314 17554
rect 15374 17502 15426 17554
rect 17054 17502 17106 17554
rect 21310 17502 21362 17554
rect 21646 17502 21698 17554
rect 22766 17502 22818 17554
rect 32398 17502 32450 17554
rect 36094 17502 36146 17554
rect 38446 17502 38498 17554
rect 39454 17502 39506 17554
rect 39678 17502 39730 17554
rect 40798 17502 40850 17554
rect 40910 17502 40962 17554
rect 42254 17502 42306 17554
rect 42590 17502 42642 17554
rect 43710 17502 43762 17554
rect 47182 17502 47234 17554
rect 48414 17502 48466 17554
rect 49534 17502 49586 17554
rect 52110 17502 52162 17554
rect 53230 17502 53282 17554
rect 53678 17502 53730 17554
rect 54462 17502 54514 17554
rect 55358 17502 55410 17554
rect 59390 17502 59442 17554
rect 60958 17502 61010 17554
rect 61294 17502 61346 17554
rect 2494 17390 2546 17442
rect 2830 17390 2882 17442
rect 4958 17390 5010 17442
rect 5854 17390 5906 17442
rect 6302 17390 6354 17442
rect 11678 17390 11730 17442
rect 35086 17390 35138 17442
rect 35310 17390 35362 17442
rect 35646 17390 35698 17442
rect 35870 17390 35922 17442
rect 38894 17390 38946 17442
rect 41470 17390 41522 17442
rect 43150 17390 43202 17442
rect 43598 17390 43650 17442
rect 44046 17390 44098 17442
rect 48862 17390 48914 17442
rect 48974 17390 49026 17442
rect 49982 17390 50034 17442
rect 54350 17390 54402 17442
rect 57934 17390 57986 17442
rect 62078 17390 62130 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 2606 17054 2658 17106
rect 2942 17054 2994 17106
rect 3950 17054 4002 17106
rect 4398 17054 4450 17106
rect 5630 17054 5682 17106
rect 5854 17054 5906 17106
rect 8878 17054 8930 17106
rect 11006 17054 11058 17106
rect 13918 17054 13970 17106
rect 15486 17054 15538 17106
rect 16606 17054 16658 17106
rect 17614 17054 17666 17106
rect 18734 17054 18786 17106
rect 18958 17054 19010 17106
rect 24334 17054 24386 17106
rect 24558 17054 24610 17106
rect 26014 17054 26066 17106
rect 30382 17054 30434 17106
rect 33854 17054 33906 17106
rect 34078 17054 34130 17106
rect 36766 17054 36818 17106
rect 40350 17054 40402 17106
rect 46174 17054 46226 17106
rect 47070 17054 47122 17106
rect 49310 17054 49362 17106
rect 53790 17054 53842 17106
rect 54574 17054 54626 17106
rect 56030 17054 56082 17106
rect 56590 17054 56642 17106
rect 60510 17054 60562 17106
rect 60846 17054 60898 17106
rect 61182 17054 61234 17106
rect 61518 17054 61570 17106
rect 62190 17054 62242 17106
rect 4846 16942 4898 16994
rect 5070 16942 5122 16994
rect 6414 16942 6466 16994
rect 6974 16942 7026 16994
rect 7982 16942 8034 16994
rect 8318 16942 8370 16994
rect 14478 16942 14530 16994
rect 14926 16942 14978 16994
rect 16270 16942 16322 16994
rect 16718 16942 16770 16994
rect 17950 16942 18002 16994
rect 19070 16942 19122 16994
rect 20414 16942 20466 16994
rect 23886 16942 23938 16994
rect 24670 16942 24722 16994
rect 25454 16942 25506 16994
rect 25790 16942 25842 16994
rect 26686 16942 26738 16994
rect 27022 16942 27074 16994
rect 28142 16942 28194 16994
rect 31614 16942 31666 16994
rect 32062 16942 32114 16994
rect 32174 16942 32226 16994
rect 33518 16942 33570 16994
rect 34750 16942 34802 16994
rect 37214 16942 37266 16994
rect 38894 16942 38946 16994
rect 39006 16942 39058 16994
rect 41358 16942 41410 16994
rect 41918 16942 41970 16994
rect 43262 16942 43314 16994
rect 46510 16942 46562 16994
rect 47406 16942 47458 16994
rect 54798 16942 54850 16994
rect 55470 16942 55522 16994
rect 55806 16942 55858 16994
rect 55918 16942 55970 16994
rect 57598 16942 57650 16994
rect 57710 16942 57762 16994
rect 59390 16942 59442 16994
rect 61854 16942 61906 16994
rect 5182 16830 5234 16882
rect 5518 16830 5570 16882
rect 6190 16830 6242 16882
rect 6862 16830 6914 16882
rect 7422 16830 7474 16882
rect 10110 16830 10162 16882
rect 12910 16830 12962 16882
rect 14254 16830 14306 16882
rect 15486 16830 15538 16882
rect 15934 16830 15986 16882
rect 18174 16830 18226 16882
rect 18398 16830 18450 16882
rect 19518 16830 19570 16882
rect 20526 16830 20578 16882
rect 21982 16830 22034 16882
rect 23550 16830 23602 16882
rect 24110 16830 24162 16882
rect 25566 16830 25618 16882
rect 27246 16830 27298 16882
rect 27582 16830 27634 16882
rect 29038 16830 29090 16882
rect 29934 16830 29986 16882
rect 30942 16830 30994 16882
rect 31278 16830 31330 16882
rect 33294 16830 33346 16882
rect 34526 16830 34578 16882
rect 34974 16830 35026 16882
rect 35310 16830 35362 16882
rect 35534 16830 35586 16882
rect 35870 16830 35922 16882
rect 36094 16830 36146 16882
rect 37550 16830 37602 16882
rect 37886 16830 37938 16882
rect 39230 16830 39282 16882
rect 39678 16830 39730 16882
rect 39902 16830 39954 16882
rect 41134 16830 41186 16882
rect 41470 16830 41522 16882
rect 41806 16830 41858 16882
rect 42142 16830 42194 16882
rect 42590 16830 42642 16882
rect 44270 16830 44322 16882
rect 45726 16830 45778 16882
rect 47630 16830 47682 16882
rect 47966 16830 48018 16882
rect 48750 16830 48802 16882
rect 49758 16830 49810 16882
rect 50206 16830 50258 16882
rect 53678 16830 53730 16882
rect 54350 16830 54402 16882
rect 55582 16830 55634 16882
rect 57150 16830 57202 16882
rect 57374 16830 57426 16882
rect 2158 16718 2210 16770
rect 3502 16718 3554 16770
rect 7198 16718 7250 16770
rect 8542 16718 8594 16770
rect 18286 16718 18338 16770
rect 19070 16718 19122 16770
rect 21870 16718 21922 16770
rect 23998 16718 24050 16770
rect 25678 16718 25730 16770
rect 33966 16718 34018 16770
rect 34862 16718 34914 16770
rect 35758 16718 35810 16770
rect 39790 16718 39842 16770
rect 46734 16718 46786 16770
rect 50878 16718 50930 16770
rect 53006 16718 53058 16770
rect 54462 16718 54514 16770
rect 2158 16606 2210 16658
rect 3278 16606 3330 16658
rect 15822 16606 15874 16658
rect 20302 16606 20354 16658
rect 28254 16606 28306 16658
rect 29710 16606 29762 16658
rect 32062 16606 32114 16658
rect 38110 16606 38162 16658
rect 38446 16606 38498 16658
rect 38894 16606 38946 16658
rect 42926 16606 42978 16658
rect 47294 16606 47346 16658
rect 48974 16606 49026 16658
rect 58158 16606 58210 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 10222 16270 10274 16322
rect 12126 16270 12178 16322
rect 12350 16270 12402 16322
rect 12910 16270 12962 16322
rect 13918 16270 13970 16322
rect 15374 16270 15426 16322
rect 30270 16270 30322 16322
rect 45054 16270 45106 16322
rect 49086 16270 49138 16322
rect 50206 16270 50258 16322
rect 55470 16270 55522 16322
rect 2270 16158 2322 16210
rect 3166 16158 3218 16210
rect 3614 16158 3666 16210
rect 6638 16158 6690 16210
rect 10670 16158 10722 16210
rect 13582 16158 13634 16210
rect 20638 16158 20690 16210
rect 26686 16158 26738 16210
rect 30718 16158 30770 16210
rect 36430 16158 36482 16210
rect 39342 16158 39394 16210
rect 41470 16158 41522 16210
rect 41918 16158 41970 16210
rect 47406 16158 47458 16210
rect 49534 16158 49586 16210
rect 49870 16158 49922 16210
rect 50766 16158 50818 16210
rect 51438 16158 51490 16210
rect 51886 16158 51938 16210
rect 54574 16158 54626 16210
rect 58046 16158 58098 16210
rect 58382 16158 58434 16210
rect 59278 16158 59330 16210
rect 60622 16158 60674 16210
rect 61518 16158 61570 16210
rect 61966 16158 62018 16210
rect 3950 16046 4002 16098
rect 4622 16046 4674 16098
rect 4734 16046 4786 16098
rect 5182 16046 5234 16098
rect 6078 16046 6130 16098
rect 7422 16046 7474 16098
rect 8990 16046 9042 16098
rect 9886 16046 9938 16098
rect 11118 16046 11170 16098
rect 12686 16046 12738 16098
rect 13470 16046 13522 16098
rect 14030 16046 14082 16098
rect 14478 16046 14530 16098
rect 14702 16046 14754 16098
rect 15710 16046 15762 16098
rect 15934 16046 15986 16098
rect 18958 16046 19010 16098
rect 20302 16046 20354 16098
rect 21310 16046 21362 16098
rect 23102 16046 23154 16098
rect 26126 16046 26178 16098
rect 28366 16046 28418 16098
rect 28478 16046 28530 16098
rect 29150 16046 29202 16098
rect 29486 16046 29538 16098
rect 29598 16046 29650 16098
rect 29934 16046 29986 16098
rect 31502 16046 31554 16098
rect 31726 16046 31778 16098
rect 32062 16046 32114 16098
rect 32622 16046 32674 16098
rect 32958 16046 33010 16098
rect 33518 16046 33570 16098
rect 37550 16046 37602 16098
rect 38558 16046 38610 16098
rect 42366 16046 42418 16098
rect 43038 16046 43090 16098
rect 43150 16046 43202 16098
rect 44270 16046 44322 16098
rect 44830 16046 44882 16098
rect 45614 16046 45666 16098
rect 46622 16046 46674 16098
rect 47070 16046 47122 16098
rect 48190 16046 48242 16098
rect 49310 16046 49362 16098
rect 50430 16046 50482 16098
rect 54686 16046 54738 16098
rect 55358 16046 55410 16098
rect 56590 16046 56642 16098
rect 57598 16046 57650 16098
rect 58830 16046 58882 16098
rect 59502 16046 59554 16098
rect 4174 15934 4226 15986
rect 6190 15934 6242 15986
rect 9662 15934 9714 15986
rect 12574 15934 12626 15986
rect 16382 15934 16434 15986
rect 17390 15934 17442 15986
rect 21758 15934 21810 15986
rect 23438 15934 23490 15986
rect 27358 15934 27410 15986
rect 27694 15934 27746 15986
rect 28030 15934 28082 15986
rect 29262 15934 29314 15986
rect 30158 15934 30210 15986
rect 30942 15934 30994 15986
rect 33070 15934 33122 15986
rect 34302 15934 34354 15986
rect 37102 15934 37154 15986
rect 37774 15934 37826 15986
rect 38110 15934 38162 15986
rect 42142 15934 42194 15986
rect 42814 15934 42866 15986
rect 45390 15934 45442 15986
rect 47854 15934 47906 15986
rect 48414 15934 48466 15986
rect 49646 15934 49698 15986
rect 50878 15934 50930 15986
rect 53118 15934 53170 15986
rect 2718 15822 2770 15874
rect 4958 15822 5010 15874
rect 14814 15822 14866 15874
rect 16270 15822 16322 15874
rect 24110 15822 24162 15874
rect 25230 15822 25282 15874
rect 26574 15822 26626 15874
rect 26798 15822 26850 15874
rect 28142 15822 28194 15874
rect 33294 15822 33346 15874
rect 36990 15822 37042 15874
rect 38222 15822 38274 15874
rect 44830 15822 44882 15874
rect 46062 15822 46114 15874
rect 48078 15822 48130 15874
rect 50654 15822 50706 15874
rect 52782 15822 52834 15874
rect 61070 15822 61122 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 2046 15486 2098 15538
rect 2494 15486 2546 15538
rect 3838 15486 3890 15538
rect 4286 15486 4338 15538
rect 5630 15486 5682 15538
rect 13022 15486 13074 15538
rect 13918 15486 13970 15538
rect 16494 15486 16546 15538
rect 22542 15486 22594 15538
rect 24670 15486 24722 15538
rect 25230 15486 25282 15538
rect 25566 15486 25618 15538
rect 30718 15486 30770 15538
rect 32062 15486 32114 15538
rect 34414 15486 34466 15538
rect 37662 15486 37714 15538
rect 38782 15486 38834 15538
rect 41806 15486 41858 15538
rect 49310 15486 49362 15538
rect 50430 15486 50482 15538
rect 55918 15486 55970 15538
rect 59950 15486 60002 15538
rect 60398 15486 60450 15538
rect 60846 15486 60898 15538
rect 61406 15486 61458 15538
rect 61742 15486 61794 15538
rect 62190 15486 62242 15538
rect 4510 15374 4562 15426
rect 5294 15374 5346 15426
rect 5518 15374 5570 15426
rect 7086 15374 7138 15426
rect 9662 15374 9714 15426
rect 12014 15374 12066 15426
rect 13806 15374 13858 15426
rect 14814 15374 14866 15426
rect 17390 15374 17442 15426
rect 20190 15374 20242 15426
rect 21534 15374 21586 15426
rect 28702 15374 28754 15426
rect 33182 15374 33234 15426
rect 33518 15374 33570 15426
rect 35534 15374 35586 15426
rect 41470 15374 41522 15426
rect 41694 15374 41746 15426
rect 42926 15374 42978 15426
rect 46622 15374 46674 15426
rect 47854 15374 47906 15426
rect 50094 15374 50146 15426
rect 50990 15374 51042 15426
rect 51214 15374 51266 15426
rect 51550 15374 51602 15426
rect 53566 15374 53618 15426
rect 54910 15374 54962 15426
rect 55358 15374 55410 15426
rect 4846 15262 4898 15314
rect 5742 15262 5794 15314
rect 6078 15262 6130 15314
rect 6302 15262 6354 15314
rect 7310 15262 7362 15314
rect 8430 15262 8482 15314
rect 8878 15262 8930 15314
rect 9550 15262 9602 15314
rect 10782 15262 10834 15314
rect 11006 15262 11058 15314
rect 11454 15262 11506 15314
rect 11790 15262 11842 15314
rect 12574 15262 12626 15314
rect 12910 15262 12962 15314
rect 13246 15262 13298 15314
rect 21422 15262 21474 15314
rect 23438 15262 23490 15314
rect 24334 15262 24386 15314
rect 27470 15262 27522 15314
rect 28926 15262 28978 15314
rect 33630 15262 33682 15314
rect 34078 15262 34130 15314
rect 34526 15262 34578 15314
rect 34862 15262 34914 15314
rect 39790 15262 39842 15314
rect 40014 15262 40066 15314
rect 40462 15262 40514 15314
rect 42030 15262 42082 15314
rect 43598 15262 43650 15314
rect 44046 15262 44098 15314
rect 44270 15262 44322 15314
rect 48862 15262 48914 15314
rect 48974 15262 49026 15314
rect 49310 15262 49362 15314
rect 49870 15262 49922 15314
rect 50430 15262 50482 15314
rect 51886 15262 51938 15314
rect 56590 15262 56642 15314
rect 2830 15150 2882 15202
rect 3390 15150 3442 15202
rect 7086 15150 7138 15202
rect 10110 15150 10162 15202
rect 11902 15150 11954 15202
rect 13134 15150 13186 15202
rect 17838 15150 17890 15202
rect 18734 15150 18786 15202
rect 23214 15150 23266 15202
rect 23774 15150 23826 15202
rect 24110 15150 24162 15202
rect 27694 15150 27746 15202
rect 39902 15150 39954 15202
rect 41694 15150 41746 15202
rect 49646 15150 49698 15202
rect 52334 15150 52386 15202
rect 55582 15150 55634 15202
rect 57374 15150 57426 15202
rect 59502 15150 59554 15202
rect 14030 15038 14082 15090
rect 22206 15038 22258 15090
rect 26910 15038 26962 15090
rect 33070 15038 33122 15090
rect 34302 15038 34354 15090
rect 37326 15038 37378 15090
rect 45278 15038 45330 15090
rect 50654 15038 50706 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 13582 14702 13634 14754
rect 22430 14702 22482 14754
rect 22654 14702 22706 14754
rect 31166 14702 31218 14754
rect 33406 14702 33458 14754
rect 34526 14702 34578 14754
rect 35534 14702 35586 14754
rect 44942 14702 44994 14754
rect 47182 14702 47234 14754
rect 53118 14702 53170 14754
rect 53454 14702 53506 14754
rect 53902 14702 53954 14754
rect 2494 14590 2546 14642
rect 3838 14590 3890 14642
rect 4286 14590 4338 14642
rect 4958 14590 5010 14642
rect 6302 14590 6354 14642
rect 10894 14590 10946 14642
rect 13694 14590 13746 14642
rect 18622 14590 18674 14642
rect 21870 14590 21922 14642
rect 29262 14590 29314 14642
rect 33294 14590 33346 14642
rect 35982 14590 36034 14642
rect 37102 14590 37154 14642
rect 41246 14590 41298 14642
rect 43374 14590 43426 14642
rect 44270 14590 44322 14642
rect 48190 14590 48242 14642
rect 48414 14590 48466 14642
rect 55806 14590 55858 14642
rect 57598 14590 57650 14642
rect 58718 14590 58770 14642
rect 61070 14590 61122 14642
rect 61630 14590 61682 14642
rect 62190 14590 62242 14642
rect 3278 14478 3330 14530
rect 5966 14478 6018 14530
rect 6190 14478 6242 14530
rect 6862 14478 6914 14530
rect 7086 14478 7138 14530
rect 9438 14478 9490 14530
rect 11230 14478 11282 14530
rect 11790 14478 11842 14530
rect 12238 14478 12290 14530
rect 14926 14478 14978 14530
rect 16270 14478 16322 14530
rect 17950 14478 18002 14530
rect 21310 14478 21362 14530
rect 21646 14478 21698 14530
rect 22094 14478 22146 14530
rect 25230 14478 25282 14530
rect 26126 14478 26178 14530
rect 26574 14478 26626 14530
rect 28142 14478 28194 14530
rect 28366 14478 28418 14530
rect 28590 14478 28642 14530
rect 29598 14478 29650 14530
rect 29934 14478 29986 14530
rect 31838 14478 31890 14530
rect 32286 14478 32338 14530
rect 33070 14478 33122 14530
rect 34414 14478 34466 14530
rect 35534 14478 35586 14530
rect 37550 14478 37602 14530
rect 38446 14478 38498 14530
rect 39230 14478 39282 14530
rect 40910 14478 40962 14530
rect 41918 14478 41970 14530
rect 42590 14478 42642 14530
rect 47518 14478 47570 14530
rect 48526 14478 48578 14530
rect 55022 14478 55074 14530
rect 55246 14478 55298 14530
rect 55918 14478 55970 14530
rect 57486 14478 57538 14530
rect 60622 14478 60674 14530
rect 4622 14366 4674 14418
rect 9886 14366 9938 14418
rect 12574 14366 12626 14418
rect 12686 14366 12738 14418
rect 13806 14366 13858 14418
rect 15598 14366 15650 14418
rect 19518 14366 19570 14418
rect 24446 14366 24498 14418
rect 30158 14366 30210 14418
rect 30382 14366 30434 14418
rect 31726 14366 31778 14418
rect 34750 14366 34802 14418
rect 34974 14366 35026 14418
rect 35870 14366 35922 14418
rect 36094 14366 36146 14418
rect 40126 14366 40178 14418
rect 41246 14366 41298 14418
rect 41358 14366 41410 14418
rect 42366 14366 42418 14418
rect 43710 14366 43762 14418
rect 46174 14366 46226 14418
rect 47070 14366 47122 14418
rect 47630 14366 47682 14418
rect 49758 14366 49810 14418
rect 52894 14366 52946 14418
rect 57710 14366 57762 14418
rect 1934 14254 1986 14306
rect 2942 14254 2994 14306
rect 4846 14254 4898 14306
rect 5070 14254 5122 14306
rect 6302 14254 6354 14306
rect 9214 14254 9266 14306
rect 14254 14254 14306 14306
rect 14590 14254 14642 14306
rect 15262 14254 15314 14306
rect 17838 14254 17890 14306
rect 20638 14254 20690 14306
rect 21422 14254 21474 14306
rect 25342 14254 25394 14306
rect 28478 14254 28530 14306
rect 29150 14254 29202 14306
rect 29598 14254 29650 14306
rect 30830 14254 30882 14306
rect 34190 14254 34242 14306
rect 37998 14254 38050 14306
rect 41134 14254 41186 14306
rect 51662 14254 51714 14306
rect 51998 14254 52050 14306
rect 57934 14254 57986 14306
rect 58606 14254 58658 14306
rect 59278 14254 59330 14306
rect 59726 14254 59778 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 2158 13918 2210 13970
rect 2718 13918 2770 13970
rect 3054 13918 3106 13970
rect 3614 13918 3666 13970
rect 7198 13918 7250 13970
rect 8878 13918 8930 13970
rect 17950 13918 18002 13970
rect 18958 13918 19010 13970
rect 21758 13918 21810 13970
rect 23998 13918 24050 13970
rect 24334 13918 24386 13970
rect 24558 13918 24610 13970
rect 25454 13918 25506 13970
rect 32286 13918 32338 13970
rect 35646 13918 35698 13970
rect 37214 13918 37266 13970
rect 38446 13918 38498 13970
rect 41134 13918 41186 13970
rect 41358 13918 41410 13970
rect 46734 13918 46786 13970
rect 47854 13918 47906 13970
rect 48862 13918 48914 13970
rect 49758 13918 49810 13970
rect 50654 13918 50706 13970
rect 58046 13918 58098 13970
rect 58494 13918 58546 13970
rect 59390 13918 59442 13970
rect 60286 13918 60338 13970
rect 61182 13918 61234 13970
rect 61742 13918 61794 13970
rect 62190 13918 62242 13970
rect 5630 13806 5682 13858
rect 7310 13806 7362 13858
rect 8542 13806 8594 13858
rect 16270 13806 16322 13858
rect 18622 13806 18674 13858
rect 19742 13806 19794 13858
rect 22318 13806 22370 13858
rect 23102 13806 23154 13858
rect 24670 13806 24722 13858
rect 26462 13806 26514 13858
rect 27582 13806 27634 13858
rect 33406 13806 33458 13858
rect 33966 13806 34018 13858
rect 35422 13806 35474 13858
rect 39342 13806 39394 13858
rect 39566 13806 39618 13858
rect 42142 13806 42194 13858
rect 49086 13806 49138 13858
rect 50206 13806 50258 13858
rect 52334 13806 52386 13858
rect 60734 13806 60786 13858
rect 4846 13694 4898 13746
rect 5854 13694 5906 13746
rect 6302 13694 6354 13746
rect 7086 13694 7138 13746
rect 7534 13694 7586 13746
rect 7870 13694 7922 13746
rect 8766 13694 8818 13746
rect 8990 13694 9042 13746
rect 9662 13694 9714 13746
rect 9998 13694 10050 13746
rect 11006 13694 11058 13746
rect 11566 13694 11618 13746
rect 12350 13694 12402 13746
rect 15038 13694 15090 13746
rect 17390 13694 17442 13746
rect 17614 13694 17666 13746
rect 22094 13694 22146 13746
rect 22878 13694 22930 13746
rect 25678 13694 25730 13746
rect 26238 13694 26290 13746
rect 26910 13694 26962 13746
rect 29934 13694 29986 13746
rect 30494 13694 30546 13746
rect 30830 13694 30882 13746
rect 31838 13694 31890 13746
rect 33294 13694 33346 13746
rect 34526 13694 34578 13746
rect 34862 13694 34914 13746
rect 35198 13694 35250 13746
rect 35982 13694 36034 13746
rect 36878 13694 36930 13746
rect 37550 13694 37602 13746
rect 38110 13694 38162 13746
rect 39902 13694 39954 13746
rect 41022 13694 41074 13746
rect 42254 13694 42306 13746
rect 43262 13694 43314 13746
rect 43710 13694 43762 13746
rect 48750 13694 48802 13746
rect 49198 13694 49250 13746
rect 49534 13694 49586 13746
rect 49982 13694 50034 13746
rect 50990 13694 51042 13746
rect 51214 13694 51266 13746
rect 51438 13694 51490 13746
rect 51774 13694 51826 13746
rect 52558 13694 52610 13746
rect 53342 13694 53394 13746
rect 54574 13694 54626 13746
rect 55358 13694 55410 13746
rect 56590 13694 56642 13746
rect 56814 13694 56866 13746
rect 57150 13694 57202 13746
rect 59838 13694 59890 13746
rect 3950 13582 4002 13634
rect 4174 13582 4226 13634
rect 4622 13582 4674 13634
rect 14478 13582 14530 13634
rect 21534 13582 21586 13634
rect 23662 13582 23714 13634
rect 29710 13582 29762 13634
rect 30382 13582 30434 13634
rect 37886 13582 37938 13634
rect 53902 13582 53954 13634
rect 57598 13582 57650 13634
rect 58942 13582 58994 13634
rect 6638 13470 6690 13522
rect 7982 13470 8034 13522
rect 8206 13470 8258 13522
rect 10782 13470 10834 13522
rect 35646 13470 35698 13522
rect 36318 13470 36370 13522
rect 36654 13470 36706 13522
rect 40238 13470 40290 13522
rect 44494 13470 44546 13522
rect 45390 13470 45442 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 1598 13134 1650 13186
rect 2942 13134 2994 13186
rect 4958 13134 5010 13186
rect 7534 13134 7586 13186
rect 15598 13134 15650 13186
rect 16830 13134 16882 13186
rect 23214 13134 23266 13186
rect 35534 13134 35586 13186
rect 38894 13134 38946 13186
rect 41918 13134 41970 13186
rect 45390 13134 45442 13186
rect 45838 13134 45890 13186
rect 54686 13134 54738 13186
rect 2046 13022 2098 13074
rect 2942 13022 2994 13074
rect 7646 13022 7698 13074
rect 9214 13022 9266 13074
rect 9886 13022 9938 13074
rect 12014 13022 12066 13074
rect 17950 13022 18002 13074
rect 18958 13022 19010 13074
rect 19854 13022 19906 13074
rect 21310 13022 21362 13074
rect 29262 13022 29314 13074
rect 30158 13022 30210 13074
rect 34526 13022 34578 13074
rect 35310 13022 35362 13074
rect 38670 13022 38722 13074
rect 39230 13022 39282 13074
rect 40686 13022 40738 13074
rect 43374 13022 43426 13074
rect 45390 13022 45442 13074
rect 46846 13022 46898 13074
rect 49982 13022 50034 13074
rect 51438 13022 51490 13074
rect 53342 13022 53394 13074
rect 56926 13022 56978 13074
rect 57374 13022 57426 13074
rect 57822 13022 57874 13074
rect 58830 13022 58882 13074
rect 59166 13022 59218 13074
rect 59614 13022 59666 13074
rect 61854 13022 61906 13074
rect 62302 13022 62354 13074
rect 5966 12910 6018 12962
rect 6190 12910 6242 12962
rect 8654 12910 8706 12962
rect 8990 12910 9042 12962
rect 12686 12910 12738 12962
rect 16606 12910 16658 12962
rect 17054 12910 17106 12962
rect 20638 12910 20690 12962
rect 21422 12910 21474 12962
rect 21646 12910 21698 12962
rect 22654 12910 22706 12962
rect 22878 12910 22930 12962
rect 23438 12910 23490 12962
rect 23998 12910 24050 12962
rect 24334 12910 24386 12962
rect 25006 12910 25058 12962
rect 25902 12910 25954 12962
rect 29710 12910 29762 12962
rect 31054 12910 31106 12962
rect 31278 12910 31330 12962
rect 34414 12910 34466 12962
rect 35198 12910 35250 12962
rect 35534 12910 35586 12962
rect 37438 12910 37490 12962
rect 41022 12910 41074 12962
rect 41470 12910 41522 12962
rect 42702 12910 42754 12962
rect 43822 12910 43874 12962
rect 46734 12910 46786 12962
rect 47294 12910 47346 12962
rect 47742 12910 47794 12962
rect 50990 12910 51042 12962
rect 51662 12910 51714 12962
rect 54126 12910 54178 12962
rect 55022 12910 55074 12962
rect 56590 12910 56642 12962
rect 3838 12798 3890 12850
rect 5630 12798 5682 12850
rect 6526 12798 6578 12850
rect 7982 12798 8034 12850
rect 14030 12798 14082 12850
rect 17390 12798 17442 12850
rect 18174 12798 18226 12850
rect 18510 12798 18562 12850
rect 18734 12798 18786 12850
rect 19070 12798 19122 12850
rect 19518 12798 19570 12850
rect 20414 12798 20466 12850
rect 21870 12798 21922 12850
rect 23774 12798 23826 12850
rect 24670 12798 24722 12850
rect 27806 12798 27858 12850
rect 30606 12798 30658 12850
rect 34078 12798 34130 12850
rect 37662 12798 37714 12850
rect 37998 12798 38050 12850
rect 44270 12798 44322 12850
rect 44942 12798 44994 12850
rect 46062 12798 46114 12850
rect 47630 12798 47682 12850
rect 48302 12798 48354 12850
rect 48526 12798 48578 12850
rect 49198 12798 49250 12850
rect 50542 12798 50594 12850
rect 50654 12798 50706 12850
rect 54014 12798 54066 12850
rect 55246 12798 55298 12850
rect 55806 12798 55858 12850
rect 56254 12798 56306 12850
rect 56366 12798 56418 12850
rect 58270 12798 58322 12850
rect 2494 12686 2546 12738
rect 5742 12686 5794 12738
rect 9662 12686 9714 12738
rect 16942 12686 16994 12738
rect 22094 12686 22146 12738
rect 23102 12686 23154 12738
rect 24222 12686 24274 12738
rect 25790 12686 25842 12738
rect 26350 12686 26402 12738
rect 29150 12686 29202 12738
rect 29374 12686 29426 12738
rect 37102 12686 37154 12738
rect 49534 12686 49586 12738
rect 50318 12686 50370 12738
rect 50430 12686 50482 12738
rect 51998 12686 52050 12738
rect 53006 12686 53058 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 3278 12350 3330 12402
rect 4510 12350 4562 12402
rect 11230 12350 11282 12402
rect 16382 12350 16434 12402
rect 17614 12350 17666 12402
rect 18398 12350 18450 12402
rect 23774 12350 23826 12402
rect 25342 12350 25394 12402
rect 27134 12350 27186 12402
rect 28254 12350 28306 12402
rect 29934 12350 29986 12402
rect 35870 12350 35922 12402
rect 38334 12350 38386 12402
rect 40014 12350 40066 12402
rect 41470 12350 41522 12402
rect 44158 12350 44210 12402
rect 45054 12350 45106 12402
rect 49198 12350 49250 12402
rect 55134 12350 55186 12402
rect 55470 12350 55522 12402
rect 56590 12350 56642 12402
rect 57934 12350 57986 12402
rect 58830 12350 58882 12402
rect 59614 12350 59666 12402
rect 2046 12238 2098 12290
rect 4062 12238 4114 12290
rect 10334 12238 10386 12290
rect 13134 12238 13186 12290
rect 13582 12238 13634 12290
rect 15262 12238 15314 12290
rect 15934 12238 15986 12290
rect 16830 12238 16882 12290
rect 18622 12238 18674 12290
rect 18734 12238 18786 12290
rect 19630 12238 19682 12290
rect 20190 12238 20242 12290
rect 22094 12238 22146 12290
rect 22318 12238 22370 12290
rect 22990 12238 23042 12290
rect 23214 12238 23266 12290
rect 24334 12238 24386 12290
rect 26126 12238 26178 12290
rect 29262 12238 29314 12290
rect 33182 12238 33234 12290
rect 33294 12238 33346 12290
rect 33966 12238 34018 12290
rect 39118 12238 39170 12290
rect 41246 12238 41298 12290
rect 41694 12238 41746 12290
rect 43374 12238 43426 12290
rect 44718 12238 44770 12290
rect 47182 12238 47234 12290
rect 49758 12238 49810 12290
rect 51214 12238 51266 12290
rect 52670 12238 52722 12290
rect 53342 12238 53394 12290
rect 56926 12238 56978 12290
rect 1710 12126 1762 12178
rect 6078 12126 6130 12178
rect 8206 12126 8258 12178
rect 8542 12126 8594 12178
rect 9550 12126 9602 12178
rect 10222 12126 10274 12178
rect 12462 12126 12514 12178
rect 13022 12126 13074 12178
rect 13246 12126 13298 12178
rect 13806 12126 13858 12178
rect 14254 12126 14306 12178
rect 14590 12126 14642 12178
rect 15038 12126 15090 12178
rect 15598 12126 15650 12178
rect 16270 12126 16322 12178
rect 16494 12126 16546 12178
rect 17390 12126 17442 12178
rect 17838 12126 17890 12178
rect 17950 12126 18002 12178
rect 19070 12126 19122 12178
rect 19742 12126 19794 12178
rect 20078 12126 20130 12178
rect 20750 12126 20802 12178
rect 21086 12126 21138 12178
rect 22766 12126 22818 12178
rect 23438 12126 23490 12178
rect 23662 12126 23714 12178
rect 24110 12126 24162 12178
rect 24782 12126 24834 12178
rect 25342 12126 25394 12178
rect 25678 12126 25730 12178
rect 25902 12126 25954 12178
rect 28926 12126 28978 12178
rect 30606 12126 30658 12178
rect 31950 12126 32002 12178
rect 32958 12126 33010 12178
rect 36094 12126 36146 12178
rect 37326 12126 37378 12178
rect 37886 12126 37938 12178
rect 38894 12126 38946 12178
rect 39678 12126 39730 12178
rect 41918 12126 41970 12178
rect 42702 12126 42754 12178
rect 44270 12126 44322 12178
rect 45054 12126 45106 12178
rect 45614 12126 45666 12178
rect 46174 12126 46226 12178
rect 46958 12126 47010 12178
rect 47966 12126 48018 12178
rect 48190 12126 48242 12178
rect 48750 12126 48802 12178
rect 48974 12126 49026 12178
rect 49310 12126 49362 12178
rect 50542 12126 50594 12178
rect 52222 12126 52274 12178
rect 55694 12126 55746 12178
rect 58270 12126 58322 12178
rect 2830 12014 2882 12066
rect 3726 12014 3778 12066
rect 4958 12014 5010 12066
rect 5966 12014 6018 12066
rect 7870 12014 7922 12066
rect 10110 12014 10162 12066
rect 11790 12014 11842 12066
rect 14030 12014 14082 12066
rect 19182 12014 19234 12066
rect 20862 12014 20914 12066
rect 22542 12014 22594 12066
rect 24558 12014 24610 12066
rect 41806 12014 41858 12066
rect 42590 12014 42642 12066
rect 47070 12014 47122 12066
rect 57374 12014 57426 12066
rect 59166 12014 59218 12066
rect 4174 11902 4226 11954
rect 11566 11902 11618 11954
rect 12686 11902 12738 11954
rect 14478 11902 14530 11954
rect 19630 11902 19682 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 6862 11566 6914 11618
rect 12126 11566 12178 11618
rect 12798 11566 12850 11618
rect 12910 11566 12962 11618
rect 16830 11566 16882 11618
rect 28030 11566 28082 11618
rect 28366 11566 28418 11618
rect 30606 11566 30658 11618
rect 34302 11566 34354 11618
rect 37550 11566 37602 11618
rect 38110 11566 38162 11618
rect 50542 11566 50594 11618
rect 55582 11566 55634 11618
rect 56254 11566 56306 11618
rect 56702 11566 56754 11618
rect 2494 11454 2546 11506
rect 9886 11454 9938 11506
rect 11790 11454 11842 11506
rect 16270 11454 16322 11506
rect 17838 11454 17890 11506
rect 25118 11454 25170 11506
rect 29598 11454 29650 11506
rect 31838 11454 31890 11506
rect 33406 11454 33458 11506
rect 35870 11454 35922 11506
rect 36990 11454 37042 11506
rect 37214 11454 37266 11506
rect 42814 11454 42866 11506
rect 44942 11454 44994 11506
rect 46174 11454 46226 11506
rect 46846 11454 46898 11506
rect 49086 11454 49138 11506
rect 49422 11454 49474 11506
rect 56254 11454 56306 11506
rect 56702 11454 56754 11506
rect 57150 11454 57202 11506
rect 57598 11454 57650 11506
rect 58046 11454 58098 11506
rect 5742 11342 5794 11394
rect 6526 11342 6578 11394
rect 7422 11342 7474 11394
rect 7758 11342 7810 11394
rect 10782 11342 10834 11394
rect 12350 11342 12402 11394
rect 13358 11342 13410 11394
rect 16718 11342 16770 11394
rect 17054 11342 17106 11394
rect 17614 11342 17666 11394
rect 17950 11342 18002 11394
rect 19070 11342 19122 11394
rect 19518 11342 19570 11394
rect 20302 11342 20354 11394
rect 21870 11342 21922 11394
rect 22318 11342 22370 11394
rect 25678 11342 25730 11394
rect 26574 11342 26626 11394
rect 26798 11342 26850 11394
rect 27358 11342 27410 11394
rect 29150 11342 29202 11394
rect 31390 11342 31442 11394
rect 32286 11342 32338 11394
rect 33294 11342 33346 11394
rect 33518 11342 33570 11394
rect 35086 11342 35138 11394
rect 40350 11342 40402 11394
rect 41246 11342 41298 11394
rect 41806 11342 41858 11394
rect 42030 11342 42082 11394
rect 42366 11342 42418 11394
rect 43038 11342 43090 11394
rect 43262 11342 43314 11394
rect 44158 11342 44210 11394
rect 45390 11342 45442 11394
rect 46398 11342 46450 11394
rect 47630 11342 47682 11394
rect 47966 11342 48018 11394
rect 48974 11342 49026 11394
rect 49870 11342 49922 11394
rect 50878 11342 50930 11394
rect 51102 11342 51154 11394
rect 51774 11342 51826 11394
rect 3614 11230 3666 11282
rect 4958 11230 5010 11282
rect 5854 11230 5906 11282
rect 10446 11230 10498 11282
rect 12686 11230 12738 11282
rect 15150 11230 15202 11282
rect 16494 11230 16546 11282
rect 18622 11230 18674 11282
rect 18958 11230 19010 11282
rect 20750 11230 20802 11282
rect 22990 11230 23042 11282
rect 25902 11230 25954 11282
rect 27246 11230 27298 11282
rect 30382 11230 30434 11282
rect 34862 11230 34914 11282
rect 39454 11230 39506 11282
rect 40686 11230 40738 11282
rect 41470 11230 41522 11282
rect 42702 11230 42754 11282
rect 44830 11230 44882 11282
rect 45166 11230 45218 11282
rect 45726 11230 45778 11282
rect 45950 11230 46002 11282
rect 47182 11230 47234 11282
rect 47406 11230 47458 11282
rect 49086 11230 49138 11282
rect 53118 11230 53170 11282
rect 54238 11230 54290 11282
rect 20638 11118 20690 11170
rect 21310 11118 21362 11170
rect 26350 11118 26402 11170
rect 26686 11118 26738 11170
rect 32734 11118 32786 11170
rect 33070 11118 33122 11170
rect 33966 11118 34018 11170
rect 36430 11118 36482 11170
rect 40574 11118 40626 11170
rect 41918 11118 41970 11170
rect 44046 11118 44098 11170
rect 47518 11118 47570 11170
rect 48302 11118 48354 11170
rect 51438 11118 51490 11170
rect 52670 11118 52722 11170
rect 52782 11118 52834 11170
rect 52894 11118 52946 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4846 10782 4898 10834
rect 5182 10782 5234 10834
rect 5630 10782 5682 10834
rect 6078 10782 6130 10834
rect 6302 10782 6354 10834
rect 7758 10782 7810 10834
rect 8878 10782 8930 10834
rect 12462 10782 12514 10834
rect 13246 10782 13298 10834
rect 13470 10782 13522 10834
rect 21198 10782 21250 10834
rect 21534 10782 21586 10834
rect 21870 10782 21922 10834
rect 22094 10782 22146 10834
rect 24558 10782 24610 10834
rect 25230 10782 25282 10834
rect 25454 10782 25506 10834
rect 26350 10782 26402 10834
rect 33518 10782 33570 10834
rect 36094 10782 36146 10834
rect 36766 10782 36818 10834
rect 39790 10782 39842 10834
rect 42478 10782 42530 10834
rect 45166 10782 45218 10834
rect 46510 10782 46562 10834
rect 48078 10782 48130 10834
rect 56702 10782 56754 10834
rect 57150 10782 57202 10834
rect 5966 10670 6018 10722
rect 7422 10670 7474 10722
rect 8318 10670 8370 10722
rect 8542 10670 8594 10722
rect 11006 10670 11058 10722
rect 16382 10670 16434 10722
rect 17614 10670 17666 10722
rect 18062 10670 18114 10722
rect 22318 10670 22370 10722
rect 23214 10670 23266 10722
rect 24334 10670 24386 10722
rect 26462 10670 26514 10722
rect 27358 10670 27410 10722
rect 33182 10670 33234 10722
rect 34638 10670 34690 10722
rect 37998 10670 38050 10722
rect 41022 10670 41074 10722
rect 41694 10670 41746 10722
rect 43598 10670 43650 10722
rect 46734 10670 46786 10722
rect 47854 10670 47906 10722
rect 48190 10670 48242 10722
rect 49310 10670 49362 10722
rect 53118 10670 53170 10722
rect 6638 10558 6690 10610
rect 6862 10558 6914 10610
rect 7982 10558 8034 10610
rect 8990 10558 9042 10610
rect 9774 10558 9826 10610
rect 10222 10558 10274 10610
rect 10894 10558 10946 10610
rect 11678 10558 11730 10610
rect 11902 10558 11954 10610
rect 12462 10558 12514 10610
rect 12798 10558 12850 10610
rect 13022 10558 13074 10610
rect 15262 10558 15314 10610
rect 15486 10558 15538 10610
rect 16494 10558 16546 10610
rect 18286 10558 18338 10610
rect 18958 10558 19010 10610
rect 19518 10558 19570 10610
rect 20862 10558 20914 10610
rect 23550 10558 23602 10610
rect 23774 10558 23826 10610
rect 25678 10558 25730 10610
rect 26014 10558 26066 10610
rect 27022 10558 27074 10610
rect 28590 10558 28642 10610
rect 29934 10558 29986 10610
rect 30718 10558 30770 10610
rect 31502 10558 31554 10610
rect 33406 10558 33458 10610
rect 33630 10558 33682 10610
rect 33966 10558 34018 10610
rect 34190 10558 34242 10610
rect 34974 10558 35026 10610
rect 35198 10558 35250 10610
rect 35982 10558 36034 10610
rect 41358 10558 41410 10610
rect 42030 10558 42082 10610
rect 42254 10558 42306 10610
rect 46958 10558 47010 10610
rect 47294 10558 47346 10610
rect 47742 10558 47794 10610
rect 48974 10558 49026 10610
rect 50430 10558 50482 10610
rect 50654 10558 50706 10610
rect 52670 10558 52722 10610
rect 54126 10558 54178 10610
rect 54350 10558 54402 10610
rect 11230 10446 11282 10498
rect 13358 10446 13410 10498
rect 13918 10446 13970 10498
rect 16046 10446 16098 10498
rect 20414 10446 20466 10498
rect 21982 10446 22034 10498
rect 24670 10446 24722 10498
rect 25454 10446 25506 10498
rect 28254 10446 28306 10498
rect 31390 10446 31442 10498
rect 39230 10446 39282 10498
rect 40350 10446 40402 10498
rect 46622 10446 46674 10498
rect 7982 10334 8034 10386
rect 12238 10334 12290 10386
rect 14142 10334 14194 10386
rect 14478 10334 14530 10386
rect 18622 10334 18674 10386
rect 19182 10334 19234 10386
rect 22990 10334 23042 10386
rect 23102 10334 23154 10386
rect 31278 10334 31330 10386
rect 39342 10334 39394 10386
rect 40238 10334 40290 10386
rect 41358 10334 41410 10386
rect 42254 10334 42306 10386
rect 48862 10334 48914 10386
rect 52558 10334 52610 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 5630 9998 5682 10050
rect 6302 9998 6354 10050
rect 19742 9998 19794 10050
rect 21758 9998 21810 10050
rect 22878 9998 22930 10050
rect 31054 9998 31106 10050
rect 31726 9998 31778 10050
rect 38222 9998 38274 10050
rect 47406 9998 47458 10050
rect 50430 9998 50482 10050
rect 6302 9886 6354 9938
rect 7534 9886 7586 9938
rect 13806 9886 13858 9938
rect 16046 9886 16098 9938
rect 19182 9886 19234 9938
rect 23998 9886 24050 9938
rect 25006 9886 25058 9938
rect 26238 9886 26290 9938
rect 28030 9886 28082 9938
rect 30494 9886 30546 9938
rect 31390 9886 31442 9938
rect 34078 9886 34130 9938
rect 37886 9886 37938 9938
rect 38446 9886 38498 9938
rect 55582 9886 55634 9938
rect 56366 9886 56418 9938
rect 5966 9774 6018 9826
rect 7086 9774 7138 9826
rect 8318 9774 8370 9826
rect 8990 9774 9042 9826
rect 9774 9774 9826 9826
rect 10222 9774 10274 9826
rect 12014 9774 12066 9826
rect 14030 9774 14082 9826
rect 14702 9774 14754 9826
rect 15038 9774 15090 9826
rect 17054 9774 17106 9826
rect 17950 9774 18002 9826
rect 19294 9774 19346 9826
rect 23214 9774 23266 9826
rect 24222 9774 24274 9826
rect 25118 9774 25170 9826
rect 25566 9774 25618 9826
rect 25902 9774 25954 9826
rect 28142 9774 28194 9826
rect 29374 9774 29426 9826
rect 30270 9774 30322 9826
rect 31950 9774 32002 9826
rect 33966 9774 34018 9826
rect 34526 9774 34578 9826
rect 35422 9774 35474 9826
rect 37214 9774 37266 9826
rect 37662 9774 37714 9826
rect 38782 9774 38834 9826
rect 40126 9774 40178 9826
rect 40350 9774 40402 9826
rect 41582 9774 41634 9826
rect 42702 9774 42754 9826
rect 43598 9774 43650 9826
rect 44270 9774 44322 9826
rect 45166 9774 45218 9826
rect 45390 9774 45442 9826
rect 46398 9774 46450 9826
rect 47518 9774 47570 9826
rect 48414 9774 48466 9826
rect 51998 9774 52050 9826
rect 52782 9774 52834 9826
rect 9662 9662 9714 9714
rect 10558 9662 10610 9714
rect 11678 9662 11730 9714
rect 15262 9662 15314 9714
rect 18174 9662 18226 9714
rect 21422 9662 21474 9714
rect 21982 9662 22034 9714
rect 22542 9662 22594 9714
rect 23438 9662 23490 9714
rect 29822 9662 29874 9714
rect 29934 9662 29986 9714
rect 32958 9662 33010 9714
rect 33406 9662 33458 9714
rect 34974 9662 35026 9714
rect 35982 9662 36034 9714
rect 39118 9662 39170 9714
rect 41022 9662 41074 9714
rect 41358 9662 41410 9714
rect 43486 9662 43538 9714
rect 45726 9662 45778 9714
rect 48862 9662 48914 9714
rect 50654 9662 50706 9714
rect 51214 9662 51266 9714
rect 51662 9662 51714 9714
rect 54014 9662 54066 9714
rect 6862 9550 6914 9602
rect 8654 9550 8706 9602
rect 14366 9550 14418 9602
rect 14814 9550 14866 9602
rect 15710 9550 15762 9602
rect 15934 9550 15986 9602
rect 16158 9550 16210 9602
rect 16942 9550 16994 9602
rect 22990 9550 23042 9602
rect 32510 9550 32562 9602
rect 35534 9550 35586 9602
rect 36094 9550 36146 9602
rect 36990 9550 37042 9602
rect 37102 9550 37154 9602
rect 39678 9550 39730 9602
rect 39790 9550 39842 9602
rect 39902 9550 39954 9602
rect 41918 9550 41970 9602
rect 42478 9550 42530 9602
rect 42590 9550 42642 9602
rect 44158 9550 44210 9602
rect 44830 9550 44882 9602
rect 45838 9550 45890 9602
rect 46062 9550 46114 9602
rect 50094 9550 50146 9602
rect 55022 9550 55074 9602
rect 55918 9550 55970 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 6750 9214 6802 9266
rect 9998 9214 10050 9266
rect 13022 9214 13074 9266
rect 13134 9214 13186 9266
rect 24110 9214 24162 9266
rect 25342 9214 25394 9266
rect 25566 9214 25618 9266
rect 26350 9214 26402 9266
rect 27246 9214 27298 9266
rect 28590 9214 28642 9266
rect 28814 9214 28866 9266
rect 30942 9214 30994 9266
rect 31278 9214 31330 9266
rect 31502 9214 31554 9266
rect 31614 9214 31666 9266
rect 31726 9214 31778 9266
rect 41806 9214 41858 9266
rect 42366 9214 42418 9266
rect 43598 9214 43650 9266
rect 46062 9214 46114 9266
rect 52782 9214 52834 9266
rect 54126 9214 54178 9266
rect 54574 9214 54626 9266
rect 8878 9102 8930 9154
rect 11790 9102 11842 9154
rect 12910 9102 12962 9154
rect 15150 9102 15202 9154
rect 16382 9102 16434 9154
rect 17726 9102 17778 9154
rect 19070 9102 19122 9154
rect 23662 9102 23714 9154
rect 25230 9102 25282 9154
rect 26910 9102 26962 9154
rect 29486 9102 29538 9154
rect 29710 9102 29762 9154
rect 32398 9102 32450 9154
rect 33854 9102 33906 9154
rect 34750 9102 34802 9154
rect 35534 9102 35586 9154
rect 35646 9102 35698 9154
rect 35758 9102 35810 9154
rect 37886 9102 37938 9154
rect 40350 9102 40402 9154
rect 43150 9102 43202 9154
rect 45502 9102 45554 9154
rect 48190 9102 48242 9154
rect 51438 9102 51490 9154
rect 7310 8990 7362 9042
rect 8094 8990 8146 9042
rect 8766 8990 8818 9042
rect 13582 8990 13634 9042
rect 14142 8990 14194 9042
rect 14478 8990 14530 9042
rect 15934 8990 15986 9042
rect 17278 8990 17330 9042
rect 19742 8990 19794 9042
rect 20974 8990 21026 9042
rect 21086 8990 21138 9042
rect 21646 8990 21698 9042
rect 23214 8990 23266 9042
rect 23438 8990 23490 9042
rect 25902 8990 25954 9042
rect 26126 8990 26178 9042
rect 26574 8990 26626 9042
rect 27694 8990 27746 9042
rect 28030 8990 28082 9042
rect 28366 8990 28418 9042
rect 28702 8990 28754 9042
rect 29262 8990 29314 9042
rect 32286 8990 32338 9042
rect 32622 8990 32674 9042
rect 33406 8990 33458 9042
rect 33966 8990 34018 9042
rect 34862 8990 34914 9042
rect 35982 8990 36034 9042
rect 36542 8990 36594 9042
rect 37774 8990 37826 9042
rect 38558 8990 38610 9042
rect 38894 8990 38946 9042
rect 39118 8990 39170 9042
rect 40126 8990 40178 9042
rect 41022 8990 41074 9042
rect 41470 8990 41522 9042
rect 41694 8990 41746 9042
rect 42366 8990 42418 9042
rect 42702 8990 42754 9042
rect 42926 8990 42978 9042
rect 44158 8990 44210 9042
rect 44494 8990 44546 9042
rect 45614 8990 45666 9042
rect 46286 8990 46338 9042
rect 46734 8990 46786 9042
rect 48750 8990 48802 9042
rect 49422 8990 49474 9042
rect 51662 8990 51714 9042
rect 52670 8990 52722 9042
rect 7086 8878 7138 8930
rect 10446 8878 10498 8930
rect 18846 8878 18898 8930
rect 21758 8878 21810 8930
rect 23326 8878 23378 8930
rect 24670 8878 24722 8930
rect 26238 8878 26290 8930
rect 28142 8878 28194 8930
rect 29822 8878 29874 8930
rect 30270 8878 30322 8930
rect 33630 8878 33682 8930
rect 35870 8878 35922 8930
rect 36878 8878 36930 8930
rect 39006 8878 39058 8930
rect 39566 8878 39618 8930
rect 44942 8878 44994 8930
rect 47854 8878 47906 8930
rect 49646 8878 49698 8930
rect 53678 8878 53730 8930
rect 7758 8766 7810 8818
rect 18734 8766 18786 8818
rect 24446 8766 24498 8818
rect 30046 8766 30098 8818
rect 34750 8766 34802 8818
rect 36990 8766 37042 8818
rect 39790 8766 39842 8818
rect 40238 8766 40290 8818
rect 40910 8766 40962 8818
rect 47966 8766 48018 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 18174 8430 18226 8482
rect 47742 8430 47794 8482
rect 8318 8318 8370 8370
rect 20302 8318 20354 8370
rect 22094 8318 22146 8370
rect 24222 8318 24274 8370
rect 29934 8318 29986 8370
rect 32062 8318 32114 8370
rect 37214 8318 37266 8370
rect 37998 8318 38050 8370
rect 39902 8318 39954 8370
rect 43150 8318 43202 8370
rect 51438 8318 51490 8370
rect 51998 8318 52050 8370
rect 52894 8318 52946 8370
rect 53342 8318 53394 8370
rect 53790 8318 53842 8370
rect 7758 8206 7810 8258
rect 8206 8206 8258 8258
rect 11006 8206 11058 8258
rect 12462 8206 12514 8258
rect 12798 8206 12850 8258
rect 16270 8206 16322 8258
rect 17390 8206 17442 8258
rect 19294 8206 19346 8258
rect 19854 8206 19906 8258
rect 20078 8206 20130 8258
rect 20414 8206 20466 8258
rect 21422 8206 21474 8258
rect 24782 8206 24834 8258
rect 27134 8206 27186 8258
rect 27358 8206 27410 8258
rect 28590 8206 28642 8258
rect 29150 8206 29202 8258
rect 33294 8206 33346 8258
rect 33966 8206 34018 8258
rect 34414 8206 34466 8258
rect 35982 8206 36034 8258
rect 36990 8206 37042 8258
rect 37326 8206 37378 8258
rect 38110 8206 38162 8258
rect 39006 8206 39058 8258
rect 40238 8206 40290 8258
rect 42366 8206 42418 8258
rect 43598 8206 43650 8258
rect 45054 8206 45106 8258
rect 46510 8206 46562 8258
rect 46958 8206 47010 8258
rect 48526 8206 48578 8258
rect 48862 8206 48914 8258
rect 49086 8150 49138 8202
rect 8430 8094 8482 8146
rect 9102 8094 9154 8146
rect 11790 8094 11842 8146
rect 12238 8094 12290 8146
rect 18622 8094 18674 8146
rect 32622 8094 32674 8146
rect 32958 8094 33010 8146
rect 34638 8094 34690 8146
rect 35422 8094 35474 8146
rect 35758 8094 35810 8146
rect 39118 8094 39170 8146
rect 39790 8094 39842 8146
rect 41022 8094 41074 8146
rect 42030 8094 42082 8146
rect 45390 8094 45442 8146
rect 14142 7982 14194 8034
rect 15262 7982 15314 8034
rect 15934 7982 15986 8034
rect 26126 7982 26178 8034
rect 27694 7982 27746 8034
rect 28366 7982 28418 8034
rect 28478 7982 28530 8034
rect 33630 7982 33682 8034
rect 34302 7982 34354 8034
rect 36318 7982 36370 8034
rect 41358 7982 41410 8034
rect 49198 7982 49250 8034
rect 49310 7982 49362 8034
rect 50318 7982 50370 8034
rect 54126 7982 54178 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 8318 7646 8370 7698
rect 8542 7646 8594 7698
rect 9998 7646 10050 7698
rect 16046 7646 16098 7698
rect 16718 7646 16770 7698
rect 20414 7646 20466 7698
rect 20638 7646 20690 7698
rect 28030 7646 28082 7698
rect 30046 7646 30098 7698
rect 31166 7646 31218 7698
rect 41358 7646 41410 7698
rect 41470 7646 41522 7698
rect 42366 7646 42418 7698
rect 43710 7646 43762 7698
rect 44382 7646 44434 7698
rect 44606 7646 44658 7698
rect 45166 7646 45218 7698
rect 46734 7646 46786 7698
rect 47182 7646 47234 7698
rect 48078 7646 48130 7698
rect 51662 7646 51714 7698
rect 52110 7646 52162 7698
rect 8206 7534 8258 7586
rect 10894 7534 10946 7586
rect 13470 7534 13522 7586
rect 16606 7534 16658 7586
rect 18734 7534 18786 7586
rect 20078 7534 20130 7586
rect 20302 7534 20354 7586
rect 25678 7534 25730 7586
rect 28478 7534 28530 7586
rect 28814 7534 28866 7586
rect 29150 7534 29202 7586
rect 29934 7534 29986 7586
rect 30830 7534 30882 7586
rect 33182 7534 33234 7586
rect 39230 7534 39282 7586
rect 39342 7534 39394 7586
rect 43374 7534 43426 7586
rect 43486 7534 43538 7586
rect 44158 7534 44210 7586
rect 44494 7534 44546 7586
rect 45838 7534 45890 7586
rect 49982 7534 50034 7586
rect 12686 7422 12738 7474
rect 15934 7422 15986 7474
rect 21646 7422 21698 7474
rect 22430 7422 22482 7474
rect 22878 7422 22930 7474
rect 27806 7422 27858 7474
rect 29374 7422 29426 7474
rect 29710 7422 29762 7474
rect 30494 7422 30546 7474
rect 31054 7422 31106 7474
rect 31502 7422 31554 7474
rect 32510 7422 32562 7474
rect 33518 7422 33570 7474
rect 34078 7422 34130 7474
rect 34526 7422 34578 7474
rect 35534 7422 35586 7474
rect 36318 7422 36370 7474
rect 38110 7422 38162 7474
rect 38782 7422 38834 7474
rect 39566 7422 39618 7474
rect 40798 7422 40850 7474
rect 41246 7422 41298 7474
rect 42926 7422 42978 7474
rect 45614 7422 45666 7474
rect 46398 7422 46450 7474
rect 47406 7422 47458 7474
rect 15598 7310 15650 7362
rect 20302 7310 20354 7362
rect 23214 7310 23266 7362
rect 28926 7310 28978 7362
rect 32062 7310 32114 7362
rect 33182 7310 33234 7362
rect 35422 7310 35474 7362
rect 40350 7310 40402 7362
rect 41918 7310 41970 7362
rect 43374 7310 43426 7362
rect 48190 7310 48242 7362
rect 48862 7310 48914 7362
rect 51102 7310 51154 7362
rect 52446 7310 52498 7362
rect 52894 7310 52946 7362
rect 12238 7198 12290 7250
rect 16718 7198 16770 7250
rect 17502 7198 17554 7250
rect 21086 7198 21138 7250
rect 27470 7198 27522 7250
rect 30270 7198 30322 7250
rect 39790 7198 39842 7250
rect 40126 7198 40178 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 10558 6862 10610 6914
rect 23102 6862 23154 6914
rect 26462 6862 26514 6914
rect 26798 6862 26850 6914
rect 30046 6862 30098 6914
rect 31614 6862 31666 6914
rect 33294 6862 33346 6914
rect 42590 6862 42642 6914
rect 45390 6862 45442 6914
rect 10894 6750 10946 6802
rect 20526 6750 20578 6802
rect 22206 6750 22258 6802
rect 28478 6750 28530 6802
rect 32174 6750 32226 6802
rect 33630 6750 33682 6802
rect 35758 6750 35810 6802
rect 45054 6750 45106 6802
rect 45838 6750 45890 6802
rect 49534 6750 49586 6802
rect 9550 6638 9602 6690
rect 9662 6638 9714 6690
rect 9774 6638 9826 6690
rect 10110 6638 10162 6690
rect 11678 6638 11730 6690
rect 12462 6638 12514 6690
rect 13022 6638 13074 6690
rect 13470 6638 13522 6690
rect 14702 6638 14754 6690
rect 15822 6638 15874 6690
rect 16270 6638 16322 6690
rect 16606 6638 16658 6690
rect 16942 6638 16994 6690
rect 20190 6638 20242 6690
rect 21646 6638 21698 6690
rect 24334 6638 24386 6690
rect 24670 6638 24722 6690
rect 27246 6638 27298 6690
rect 29822 6638 29874 6690
rect 30046 6638 30098 6690
rect 32622 6638 32674 6690
rect 33518 6638 33570 6690
rect 34302 6638 34354 6690
rect 37550 6638 37602 6690
rect 43262 6638 43314 6690
rect 44270 6638 44322 6690
rect 45726 6638 45778 6690
rect 45950 6638 46002 6690
rect 47518 6638 47570 6690
rect 48414 6638 48466 6690
rect 49086 6638 49138 6690
rect 50318 6638 50370 6690
rect 50766 6638 50818 6690
rect 51214 6638 51266 6690
rect 51662 6638 51714 6690
rect 11566 6526 11618 6578
rect 13806 6526 13858 6578
rect 14366 6526 14418 6578
rect 15374 6526 15426 6578
rect 18510 6526 18562 6578
rect 19630 6526 19682 6578
rect 21310 6526 21362 6578
rect 21982 6526 22034 6578
rect 23102 6526 23154 6578
rect 23214 6526 23266 6578
rect 25006 6526 25058 6578
rect 25342 6526 25394 6578
rect 25678 6526 25730 6578
rect 26014 6526 26066 6578
rect 27582 6526 27634 6578
rect 28254 6526 28306 6578
rect 29486 6526 29538 6578
rect 29598 6526 29650 6578
rect 30942 6526 30994 6578
rect 31726 6526 31778 6578
rect 34526 6526 34578 6578
rect 35198 6526 35250 6578
rect 35310 6526 35362 6578
rect 35422 6526 35474 6578
rect 36430 6526 36482 6578
rect 39230 6526 39282 6578
rect 41806 6526 41858 6578
rect 42702 6526 42754 6578
rect 44158 6526 44210 6578
rect 44830 6526 44882 6578
rect 46174 6526 46226 6578
rect 47854 6526 47906 6578
rect 48638 6526 48690 6578
rect 48750 6526 48802 6578
rect 49982 6526 50034 6578
rect 16718 6414 16770 6466
rect 17502 6414 17554 6466
rect 23774 6414 23826 6466
rect 25230 6414 25282 6466
rect 28366 6414 28418 6466
rect 31278 6414 31330 6466
rect 34974 6414 35026 6466
rect 36318 6414 36370 6466
rect 40014 6414 40066 6466
rect 43262 6414 43314 6466
rect 47070 6414 47122 6466
rect 47294 6414 47346 6466
rect 47406 6414 47458 6466
rect 48190 6414 48242 6466
rect 52110 6414 52162 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 12462 6078 12514 6130
rect 13246 6078 13298 6130
rect 13470 6078 13522 6130
rect 14478 6078 14530 6130
rect 14926 6078 14978 6130
rect 15374 6078 15426 6130
rect 15822 6078 15874 6130
rect 16830 6078 16882 6130
rect 17502 6078 17554 6130
rect 18846 6078 18898 6130
rect 20414 6078 20466 6130
rect 20974 6078 21026 6130
rect 21422 6078 21474 6130
rect 21982 6078 22034 6130
rect 22990 6078 23042 6130
rect 23438 6078 23490 6130
rect 24334 6078 24386 6130
rect 24782 6078 24834 6130
rect 25454 6078 25506 6130
rect 26350 6078 26402 6130
rect 29934 6078 29986 6130
rect 31614 6078 31666 6130
rect 35422 6078 35474 6130
rect 39566 6078 39618 6130
rect 39790 6078 39842 6130
rect 42478 6078 42530 6130
rect 44942 6078 44994 6130
rect 45278 6078 45330 6130
rect 47182 6078 47234 6130
rect 47630 6078 47682 6130
rect 48862 6078 48914 6130
rect 49086 6078 49138 6130
rect 49422 6078 49474 6130
rect 49982 6078 50034 6130
rect 50318 6078 50370 6130
rect 13806 5966 13858 6018
rect 28142 5966 28194 6018
rect 31054 5966 31106 6018
rect 34078 5966 34130 6018
rect 35086 5966 35138 6018
rect 35198 5966 35250 6018
rect 41582 5966 41634 6018
rect 43262 5966 43314 6018
rect 46958 5966 47010 6018
rect 47966 5966 48018 6018
rect 48078 5966 48130 6018
rect 48750 5966 48802 6018
rect 19854 5854 19906 5906
rect 22430 5854 22482 5906
rect 27470 5854 27522 5906
rect 28030 5854 28082 5906
rect 28814 5854 28866 5906
rect 30158 5854 30210 5906
rect 31278 5854 31330 5906
rect 32510 5854 32562 5906
rect 33070 5854 33122 5906
rect 33294 5854 33346 5906
rect 34302 5854 34354 5906
rect 35646 5854 35698 5906
rect 38446 5854 38498 5906
rect 38782 5854 38834 5906
rect 40126 5854 40178 5906
rect 41358 5854 41410 5906
rect 41918 5854 41970 5906
rect 42142 5854 42194 5906
rect 45614 5854 45666 5906
rect 45838 5854 45890 5906
rect 46174 5854 46226 5906
rect 46846 5854 46898 5906
rect 16382 5742 16434 5794
rect 29150 5742 29202 5794
rect 32062 5742 32114 5794
rect 34526 5742 34578 5794
rect 36094 5742 36146 5794
rect 38222 5742 38274 5794
rect 39678 5742 39730 5794
rect 46398 5742 46450 5794
rect 50766 5742 50818 5794
rect 22430 5630 22482 5682
rect 23326 5630 23378 5682
rect 24110 5630 24162 5682
rect 24782 5630 24834 5682
rect 30382 5630 30434 5682
rect 30718 5630 30770 5682
rect 49646 5630 49698 5682
rect 50206 5630 50258 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 24110 5294 24162 5346
rect 25118 5294 25170 5346
rect 25678 5294 25730 5346
rect 26798 5294 26850 5346
rect 31390 5294 31442 5346
rect 31726 5294 31778 5346
rect 35646 5294 35698 5346
rect 35982 5294 36034 5346
rect 40574 5294 40626 5346
rect 45726 5294 45778 5346
rect 46062 5294 46114 5346
rect 13806 5182 13858 5234
rect 16046 5182 16098 5234
rect 16382 5182 16434 5234
rect 18846 5182 18898 5234
rect 19406 5182 19458 5234
rect 19966 5182 20018 5234
rect 20302 5182 20354 5234
rect 20862 5182 20914 5234
rect 21870 5182 21922 5234
rect 22430 5182 22482 5234
rect 22990 5182 23042 5234
rect 23662 5182 23714 5234
rect 24110 5182 24162 5234
rect 24670 5182 24722 5234
rect 25006 5182 25058 5234
rect 25678 5182 25730 5234
rect 26574 5182 26626 5234
rect 27134 5182 27186 5234
rect 31614 5182 31666 5234
rect 36990 5182 37042 5234
rect 39118 5182 39170 5234
rect 43038 5182 43090 5234
rect 47518 5182 47570 5234
rect 49646 5182 49698 5234
rect 15486 5070 15538 5122
rect 16942 5070 16994 5122
rect 27694 5070 27746 5122
rect 28254 5070 28306 5122
rect 32062 5070 32114 5122
rect 33070 5070 33122 5122
rect 33966 5070 34018 5122
rect 34974 5070 35026 5122
rect 39902 5070 39954 5122
rect 43374 5070 43426 5122
rect 43822 5070 43874 5122
rect 45054 5070 45106 5122
rect 46846 5070 46898 5122
rect 50206 5070 50258 5122
rect 27358 4958 27410 5010
rect 28030 4958 28082 5010
rect 29598 4958 29650 5010
rect 32174 4958 32226 5010
rect 34862 4958 34914 5010
rect 42030 4958 42082 5010
rect 44158 4958 44210 5010
rect 44942 4958 44994 5010
rect 21534 4846 21586 4898
rect 26126 4846 26178 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 21086 4510 21138 4562
rect 21534 4510 21586 4562
rect 21982 4510 22034 4562
rect 22766 4510 22818 4562
rect 23214 4510 23266 4562
rect 23662 4510 23714 4562
rect 24110 4510 24162 4562
rect 24670 4510 24722 4562
rect 25454 4510 25506 4562
rect 25902 4510 25954 4562
rect 26686 4510 26738 4562
rect 27022 4510 27074 4562
rect 28478 4510 28530 4562
rect 28926 4510 28978 4562
rect 29262 4510 29314 4562
rect 31390 4510 31442 4562
rect 33966 4510 34018 4562
rect 36878 4510 36930 4562
rect 41022 4510 41074 4562
rect 42142 4510 42194 4562
rect 47630 4510 47682 4562
rect 48974 4510 49026 4562
rect 30158 4398 30210 4450
rect 33070 4398 33122 4450
rect 35982 4398 36034 4450
rect 45726 4398 45778 4450
rect 47294 4398 47346 4450
rect 48078 4398 48130 4450
rect 27918 4286 27970 4338
rect 31950 4286 32002 4338
rect 32398 4286 32450 4338
rect 33406 4286 33458 4338
rect 40238 4286 40290 4338
rect 43822 4286 43874 4338
rect 46734 4286 46786 4338
rect 27582 4174 27634 4226
rect 37326 4174 37378 4226
rect 38222 4174 38274 4226
rect 49310 4174 49362 4226
rect 27582 4062 27634 4114
rect 28478 4062 28530 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 36094 3726 36146 3778
rect 38334 3726 38386 3778
rect 45950 3726 46002 3778
rect 46958 3726 47010 3778
rect 23550 3614 23602 3666
rect 24110 3614 24162 3666
rect 24782 3614 24834 3666
rect 25230 3614 25282 3666
rect 26126 3614 26178 3666
rect 27470 3614 27522 3666
rect 27918 3614 27970 3666
rect 28926 3614 28978 3666
rect 29598 3614 29650 3666
rect 31054 3614 31106 3666
rect 33518 3614 33570 3666
rect 39006 3614 39058 3666
rect 40574 3614 40626 3666
rect 42702 3614 42754 3666
rect 43822 3614 43874 3666
rect 45166 3614 45218 3666
rect 45502 3614 45554 3666
rect 46062 3614 46114 3666
rect 46510 3614 46562 3666
rect 46958 3614 47010 3666
rect 47966 3614 48018 3666
rect 48526 3614 48578 3666
rect 25678 3502 25730 3554
rect 30046 3502 30098 3554
rect 31390 3502 31442 3554
rect 33070 3502 33122 3554
rect 33406 3502 33458 3554
rect 33630 3502 33682 3554
rect 33966 3502 34018 3554
rect 34974 3502 35026 3554
rect 38446 3502 38498 3554
rect 39902 3502 39954 3554
rect 44270 3502 44322 3554
rect 47518 3502 47570 3554
rect 26574 3390 26626 3442
rect 27022 3390 27074 3442
rect 29822 3390 29874 3442
rect 31614 3390 31666 3442
rect 32398 3390 32450 3442
rect 32734 3390 32786 3442
rect 34302 3390 34354 3442
rect 34638 3390 34690 3442
rect 35534 3390 35586 3442
rect 37214 3390 37266 3442
rect 38334 3390 38386 3442
rect 44606 3390 44658 3442
rect 7646 3278 7698 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 16128 63200 16240 64000
rect 26208 63200 26320 64000
rect 29568 63200 29680 64000
rect 38304 63200 38416 64000
rect 47712 63200 47824 64000
rect 48384 63200 48496 64000
rect 11452 60564 11508 60574
rect 11340 60508 11452 60564
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 10108 57204 10164 57214
rect 5740 56980 5796 56990
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 1708 55186 1764 55198
rect 1708 55134 1710 55186
rect 1762 55134 1764 55186
rect 1708 55076 1764 55134
rect 1708 54516 1764 55020
rect 1708 54450 1764 54460
rect 2044 55074 2100 55086
rect 2044 55022 2046 55074
rect 2098 55022 2100 55074
rect 1596 53956 1652 53966
rect 1484 53508 1540 53518
rect 1484 50428 1540 53452
rect 1372 50372 1540 50428
rect 1260 48244 1316 48254
rect 1148 45556 1204 45566
rect 1148 38948 1204 45500
rect 1148 38882 1204 38892
rect 1148 30436 1204 30446
rect 924 23716 980 23726
rect 924 17780 980 23660
rect 924 17714 980 17724
rect 1148 16212 1204 30380
rect 1260 28084 1316 48188
rect 1372 33908 1428 50372
rect 1596 49812 1652 53900
rect 2044 51044 2100 55022
rect 2492 55076 2548 55086
rect 2492 54982 2548 55020
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4844 51604 4900 51614
rect 4844 51510 4900 51548
rect 2940 51268 2996 51278
rect 2940 51266 3220 51268
rect 2940 51214 2942 51266
rect 2994 51214 3220 51266
rect 2940 51212 3220 51214
rect 2940 51202 2996 51212
rect 2044 50988 2996 51044
rect 2828 50596 2884 50606
rect 1484 49756 1652 49812
rect 1932 50370 1988 50382
rect 1932 50318 1934 50370
rect 1986 50318 1988 50370
rect 1484 47012 1540 49756
rect 1820 49698 1876 49710
rect 1820 49646 1822 49698
rect 1874 49646 1876 49698
rect 1484 46946 1540 46956
rect 1596 49588 1652 49598
rect 1484 39508 1540 39518
rect 1484 36148 1540 39452
rect 1596 39172 1652 49532
rect 1820 49586 1876 49646
rect 1820 49534 1822 49586
rect 1874 49534 1876 49586
rect 1820 49522 1876 49534
rect 1932 49252 1988 50318
rect 2380 50370 2436 50382
rect 2380 50318 2382 50370
rect 2434 50318 2436 50370
rect 2380 49922 2436 50318
rect 2380 49870 2382 49922
rect 2434 49870 2436 49922
rect 1708 48804 1764 48814
rect 1708 48710 1764 48748
rect 1932 48580 1988 49196
rect 2156 49586 2212 49598
rect 2156 49534 2158 49586
rect 2210 49534 2212 49586
rect 2044 48916 2100 48926
rect 2044 48822 2100 48860
rect 1708 48524 1988 48580
rect 1708 48466 1764 48524
rect 1708 48414 1710 48466
rect 1762 48414 1764 48466
rect 1708 48402 1764 48414
rect 1932 48244 1988 48254
rect 1932 48150 1988 48188
rect 1708 48132 1764 48142
rect 1708 47458 1764 48076
rect 1708 47406 1710 47458
rect 1762 47406 1764 47458
rect 1708 47394 1764 47406
rect 1932 46562 1988 46574
rect 1932 46510 1934 46562
rect 1986 46510 1988 46562
rect 1820 45668 1876 45678
rect 1708 45666 1876 45668
rect 1708 45614 1822 45666
rect 1874 45614 1876 45666
rect 1708 45612 1876 45614
rect 1708 45108 1764 45612
rect 1820 45602 1876 45612
rect 1932 45444 1988 46510
rect 2156 45668 2212 49534
rect 2380 48244 2436 49870
rect 2828 50370 2884 50540
rect 2940 50428 2996 50988
rect 2940 50372 3108 50428
rect 2828 50318 2830 50370
rect 2882 50318 2884 50370
rect 2716 49812 2772 49822
rect 2716 49718 2772 49756
rect 2492 49252 2548 49262
rect 2492 49026 2548 49196
rect 2492 48974 2494 49026
rect 2546 48974 2548 49026
rect 2492 48962 2548 48974
rect 2716 48916 2772 48926
rect 2828 48916 2884 50318
rect 3052 50034 3108 50372
rect 3052 49982 3054 50034
rect 3106 49982 3108 50034
rect 3052 49970 3108 49982
rect 3164 49924 3220 51212
rect 4172 51266 4228 51278
rect 4172 51214 4174 51266
rect 4226 51214 4228 51266
rect 3612 50818 3668 50830
rect 3612 50766 3614 50818
rect 3666 50766 3668 50818
rect 3612 50482 3668 50766
rect 4172 50708 4228 51214
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4172 50642 4228 50652
rect 4508 50818 4564 50830
rect 4508 50766 4510 50818
rect 4562 50766 4564 50818
rect 3612 50430 3614 50482
rect 3666 50430 3668 50482
rect 3612 50418 3668 50430
rect 4396 50484 4452 50522
rect 4396 50418 4452 50428
rect 4508 50428 4564 50766
rect 5180 50596 5236 50606
rect 5180 50502 5236 50540
rect 4060 50370 4116 50382
rect 4508 50372 5012 50428
rect 4060 50318 4062 50370
rect 4114 50318 4116 50370
rect 3388 49924 3444 49934
rect 3164 49922 3444 49924
rect 3164 49870 3390 49922
rect 3442 49870 3444 49922
rect 3164 49868 3444 49870
rect 3388 49812 3444 49868
rect 3388 49746 3444 49756
rect 3948 49698 4004 49710
rect 3948 49646 3950 49698
rect 4002 49646 4004 49698
rect 3948 49588 4004 49646
rect 4060 49588 4116 50318
rect 4508 49698 4564 49710
rect 4956 49700 5012 50372
rect 4508 49646 4510 49698
rect 4562 49646 4564 49698
rect 4508 49588 4564 49646
rect 4060 49532 4564 49588
rect 4844 49698 5012 49700
rect 4844 49646 4958 49698
rect 5010 49646 5012 49698
rect 4844 49644 5012 49646
rect 3836 49140 3892 49150
rect 3724 49084 3836 49140
rect 2772 48860 2884 48916
rect 2716 48822 2772 48860
rect 2380 48178 2436 48188
rect 2492 47346 2548 47358
rect 2492 47294 2494 47346
rect 2546 47294 2548 47346
rect 2492 46900 2548 47294
rect 2492 46834 2548 46844
rect 2268 46788 2324 46798
rect 2268 46694 2324 46732
rect 2492 46676 2548 46686
rect 2380 46674 2548 46676
rect 2380 46622 2494 46674
rect 2546 46622 2548 46674
rect 2380 46620 2548 46622
rect 2380 46004 2436 46620
rect 2492 46610 2548 46620
rect 2716 46674 2772 46686
rect 2716 46622 2718 46674
rect 2770 46622 2772 46674
rect 2156 45612 2324 45668
rect 1932 45388 2212 45444
rect 1708 42756 1764 45052
rect 2044 44996 2100 45006
rect 1932 44994 2100 44996
rect 1932 44942 2046 44994
rect 2098 44942 2100 44994
rect 1932 44940 2100 44942
rect 1820 44324 1876 44334
rect 1820 44230 1876 44268
rect 1820 42756 1876 42766
rect 1708 42754 1876 42756
rect 1708 42702 1822 42754
rect 1874 42702 1876 42754
rect 1708 42700 1876 42702
rect 1820 42690 1876 42700
rect 1932 41860 1988 44940
rect 2044 44930 2100 44940
rect 2044 44212 2100 44222
rect 2044 44118 2100 44156
rect 2156 43876 2212 45388
rect 2268 44324 2324 45612
rect 2380 45106 2436 45948
rect 2604 46562 2660 46574
rect 2604 46510 2606 46562
rect 2658 46510 2660 46562
rect 2604 45780 2660 46510
rect 2716 46116 2772 46622
rect 2716 46050 2772 46060
rect 2604 45714 2660 45724
rect 2716 45444 2772 45454
rect 2380 45054 2382 45106
rect 2434 45054 2436 45106
rect 2380 45042 2436 45054
rect 2604 45218 2660 45230
rect 2604 45166 2606 45218
rect 2658 45166 2660 45218
rect 2268 44258 2324 44268
rect 2604 44324 2660 45166
rect 2716 44546 2772 45388
rect 2716 44494 2718 44546
rect 2770 44494 2772 44546
rect 2716 44482 2772 44494
rect 2380 44212 2436 44222
rect 2380 44118 2436 44156
rect 2604 44210 2660 44268
rect 2604 44158 2606 44210
rect 2658 44158 2660 44210
rect 2604 44146 2660 44158
rect 2044 43820 2212 43876
rect 2044 41972 2100 43820
rect 2156 43650 2212 43662
rect 2828 43652 2884 48860
rect 3500 48916 3556 48926
rect 3500 48822 3556 48860
rect 3164 48804 3220 48814
rect 3052 48802 3220 48804
rect 3052 48750 3166 48802
rect 3218 48750 3220 48802
rect 3052 48748 3220 48750
rect 3052 48354 3108 48748
rect 3164 48738 3220 48748
rect 3052 48302 3054 48354
rect 3106 48302 3108 48354
rect 3052 45778 3108 48302
rect 3612 46900 3668 46910
rect 3612 46786 3668 46844
rect 3612 46734 3614 46786
rect 3666 46734 3668 46786
rect 3612 46722 3668 46734
rect 3164 46452 3220 46462
rect 3164 46450 3332 46452
rect 3164 46398 3166 46450
rect 3218 46398 3332 46450
rect 3164 46396 3332 46398
rect 3164 46386 3220 46396
rect 3052 45726 3054 45778
rect 3106 45726 3108 45778
rect 3052 45714 3108 45726
rect 3164 45220 3220 45230
rect 3164 45126 3220 45164
rect 3052 45108 3108 45118
rect 3052 45014 3108 45052
rect 3052 44212 3108 44222
rect 3052 44118 3108 44156
rect 2156 43598 2158 43650
rect 2210 43598 2212 43650
rect 2156 42980 2212 43598
rect 2156 42914 2212 42924
rect 2268 43596 2884 43652
rect 3164 44098 3220 44110
rect 3164 44046 3166 44098
rect 3218 44046 3220 44098
rect 2156 42644 2212 42654
rect 2156 42550 2212 42588
rect 2044 41906 2100 41916
rect 1596 39106 1652 39116
rect 1708 41804 1988 41860
rect 2156 41860 2212 41870
rect 1596 38948 1652 38958
rect 1596 37940 1652 38892
rect 1596 37874 1652 37884
rect 1484 36082 1540 36092
rect 1708 36036 1764 41804
rect 2156 41766 2212 41804
rect 2268 41186 2324 43596
rect 3164 43428 3220 44046
rect 3276 44100 3332 46396
rect 3388 46450 3444 46462
rect 3388 46398 3390 46450
rect 3442 46398 3444 46450
rect 3388 45108 3444 46398
rect 3612 46116 3668 46126
rect 3612 45892 3668 46060
rect 3612 45826 3668 45836
rect 3724 45108 3780 49084
rect 3836 49074 3892 49084
rect 3948 48804 4004 49532
rect 3948 48738 4004 48748
rect 4060 49028 4116 49038
rect 4060 48468 4116 48972
rect 4172 48802 4228 48814
rect 4172 48750 4174 48802
rect 4226 48750 4228 48802
rect 4172 48692 4228 48750
rect 4172 48626 4228 48636
rect 4172 48468 4228 48478
rect 4060 48466 4228 48468
rect 4060 48414 4174 48466
rect 4226 48414 4228 48466
rect 4060 48412 4228 48414
rect 4172 48402 4228 48412
rect 4284 48244 4340 49532
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4508 49140 4564 49150
rect 4508 49046 4564 49084
rect 4732 49028 4788 49038
rect 4732 48934 4788 48972
rect 4620 48356 4676 48366
rect 4060 48188 4340 48244
rect 4396 48354 4676 48356
rect 4396 48302 4622 48354
rect 4674 48302 4676 48354
rect 4396 48300 4676 48302
rect 3948 47012 4004 47022
rect 3948 46786 4004 46956
rect 3948 46734 3950 46786
rect 4002 46734 4004 46786
rect 3948 46722 4004 46734
rect 3836 46676 3892 46686
rect 3836 46582 3892 46620
rect 4060 46676 4116 48188
rect 4396 48020 4452 48300
rect 4620 48290 4676 48300
rect 4060 46610 4116 46620
rect 4284 47964 4452 48020
rect 4284 46340 4340 47964
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4732 47684 4788 47694
rect 4620 47628 4732 47684
rect 4620 47570 4676 47628
rect 4732 47618 4788 47628
rect 4620 47518 4622 47570
rect 4674 47518 4676 47570
rect 4620 47506 4676 47518
rect 4844 47124 4900 49644
rect 4956 49634 5012 49644
rect 5516 49698 5572 49710
rect 5516 49646 5518 49698
rect 5570 49646 5572 49698
rect 5516 49588 5572 49646
rect 5516 49522 5572 49532
rect 5628 49140 5684 49150
rect 5628 49046 5684 49084
rect 4956 48916 5012 48926
rect 4956 48466 5012 48860
rect 4956 48414 4958 48466
rect 5010 48414 5012 48466
rect 4956 47796 5012 48414
rect 5068 48802 5124 48814
rect 5068 48750 5070 48802
rect 5122 48750 5124 48802
rect 5068 48244 5124 48750
rect 5740 48354 5796 56924
rect 8652 55076 8708 55086
rect 8652 53508 8708 55020
rect 9996 55074 10052 55086
rect 9996 55022 9998 55074
rect 10050 55022 10052 55074
rect 9548 54852 9604 54862
rect 8652 53414 8708 53452
rect 9100 53508 9156 53518
rect 9100 53414 9156 53452
rect 8540 53284 8596 53294
rect 8428 53228 8540 53284
rect 6860 52948 6916 52958
rect 6860 52274 6916 52892
rect 7756 52948 7812 52958
rect 7756 52854 7812 52892
rect 8092 52836 8148 52846
rect 7980 52834 8148 52836
rect 7980 52782 8094 52834
rect 8146 52782 8148 52834
rect 7980 52780 8148 52782
rect 6860 52222 6862 52274
rect 6914 52222 6916 52274
rect 6188 52164 6244 52174
rect 5852 51604 5908 51614
rect 5852 51510 5908 51548
rect 6188 50708 6244 52108
rect 6524 51716 6580 51726
rect 6412 51266 6468 51278
rect 6412 51214 6414 51266
rect 6466 51214 6468 51266
rect 6412 51156 6468 51214
rect 6412 51090 6468 51100
rect 6188 50706 6356 50708
rect 6188 50654 6190 50706
rect 6242 50654 6356 50706
rect 6188 50652 6356 50654
rect 6188 50642 6244 50652
rect 5964 50036 6020 50046
rect 5964 49942 6020 49980
rect 5852 49028 5908 49038
rect 5852 48934 5908 48972
rect 6188 48802 6244 48814
rect 6188 48750 6190 48802
rect 6242 48750 6244 48802
rect 5740 48302 5742 48354
rect 5794 48302 5796 48354
rect 5740 48290 5796 48302
rect 6076 48692 6132 48702
rect 5292 48244 5348 48254
rect 5068 48242 5348 48244
rect 5068 48190 5294 48242
rect 5346 48190 5348 48242
rect 5068 48188 5348 48190
rect 5292 48178 5348 48188
rect 4956 47730 5012 47740
rect 4956 47348 5012 47358
rect 4956 47254 5012 47292
rect 5404 47348 5460 47358
rect 5068 47236 5124 47246
rect 5068 47142 5124 47180
rect 4844 47068 5012 47124
rect 4508 46562 4564 46574
rect 4508 46510 4510 46562
rect 4562 46510 4564 46562
rect 4508 46452 4564 46510
rect 4508 46386 4564 46396
rect 4844 46562 4900 46574
rect 4844 46510 4846 46562
rect 4898 46510 4900 46562
rect 4060 46284 4340 46340
rect 4476 46284 4740 46294
rect 4060 45220 4116 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4844 46004 4900 46510
rect 4620 45948 4900 46004
rect 4172 45892 4228 45902
rect 4172 45330 4228 45836
rect 4508 45778 4564 45790
rect 4508 45726 4510 45778
rect 4562 45726 4564 45778
rect 4284 45666 4340 45678
rect 4284 45614 4286 45666
rect 4338 45614 4340 45666
rect 4284 45556 4340 45614
rect 4284 45490 4340 45500
rect 4508 45444 4564 45726
rect 4508 45378 4564 45388
rect 4172 45278 4174 45330
rect 4226 45278 4228 45330
rect 4172 45266 4228 45278
rect 4060 45154 4116 45164
rect 4172 45108 4228 45118
rect 3724 45052 4004 45108
rect 3388 45042 3444 45052
rect 3836 44882 3892 44894
rect 3836 44830 3838 44882
rect 3890 44830 3892 44882
rect 3500 44436 3556 44446
rect 3500 44342 3556 44380
rect 3388 44324 3444 44334
rect 3388 44230 3444 44268
rect 3612 44322 3668 44334
rect 3612 44270 3614 44322
rect 3666 44270 3668 44322
rect 3276 44034 3332 44044
rect 2828 43372 3220 43428
rect 2492 42980 2548 42990
rect 2492 42886 2548 42924
rect 2268 41134 2270 41186
rect 2322 41134 2324 41186
rect 1932 40964 1988 40974
rect 1932 40870 1988 40908
rect 2268 40740 2324 41134
rect 2268 40674 2324 40684
rect 2492 42644 2548 42654
rect 2492 40404 2548 42588
rect 2828 42642 2884 43372
rect 3612 43316 3668 44270
rect 3836 43876 3892 44830
rect 3836 43810 3892 43820
rect 3948 43762 4004 45052
rect 4172 44436 4228 45052
rect 4620 45108 4676 45948
rect 4620 45042 4676 45052
rect 4732 45778 4788 45790
rect 4732 45726 4734 45778
rect 4786 45726 4788 45778
rect 4732 44884 4788 45726
rect 4844 45668 4900 45678
rect 4844 45574 4900 45612
rect 4844 44996 4900 45006
rect 4844 44902 4900 44940
rect 4284 44828 4788 44884
rect 4284 44548 4340 44828
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4284 44492 4452 44548
rect 4172 44380 4340 44436
rect 4284 44322 4340 44380
rect 4284 44270 4286 44322
rect 4338 44270 4340 44322
rect 4284 44258 4340 44270
rect 4396 44324 4452 44492
rect 4620 44436 4676 44446
rect 4620 44342 4676 44380
rect 4396 44230 4452 44268
rect 4732 44322 4788 44334
rect 4732 44270 4734 44322
rect 4786 44270 4788 44322
rect 4172 44212 4228 44222
rect 4172 44118 4228 44156
rect 4060 44100 4116 44110
rect 4060 43876 4116 44044
rect 4060 43820 4340 43876
rect 3948 43710 3950 43762
rect 4002 43710 4004 43762
rect 3388 43260 3668 43316
rect 3724 43316 3780 43326
rect 3276 42868 3332 42878
rect 2828 42590 2830 42642
rect 2882 42590 2884 42642
rect 2828 42578 2884 42590
rect 3052 42866 3332 42868
rect 3052 42814 3278 42866
rect 3330 42814 3332 42866
rect 3052 42812 3332 42814
rect 2604 42532 2660 42542
rect 2604 42530 2772 42532
rect 2604 42478 2606 42530
rect 2658 42478 2772 42530
rect 2604 42476 2772 42478
rect 2604 42466 2660 42476
rect 2716 42420 2772 42476
rect 3052 42420 3108 42812
rect 3276 42802 3332 42812
rect 2716 42364 3108 42420
rect 3164 42642 3220 42654
rect 3164 42590 3166 42642
rect 3218 42590 3220 42642
rect 3164 42308 3220 42590
rect 3388 42644 3444 43260
rect 3724 43204 3780 43260
rect 3388 42578 3444 42588
rect 3500 43148 3780 43204
rect 3500 42642 3556 43148
rect 3724 42980 3780 42990
rect 3724 42754 3780 42924
rect 3724 42702 3726 42754
rect 3778 42702 3780 42754
rect 3724 42690 3780 42702
rect 3500 42590 3502 42642
rect 3554 42590 3556 42642
rect 3164 42242 3220 42252
rect 3276 42532 3332 42542
rect 3276 42082 3332 42476
rect 3276 42030 3278 42082
rect 3330 42030 3332 42082
rect 3276 42018 3332 42030
rect 3388 42420 3444 42430
rect 3388 42194 3444 42364
rect 3388 42142 3390 42194
rect 3442 42142 3444 42194
rect 2940 41972 2996 41982
rect 2604 41860 2660 41870
rect 2604 41858 2884 41860
rect 2604 41806 2606 41858
rect 2658 41806 2884 41858
rect 2604 41804 2884 41806
rect 2604 41794 2660 41804
rect 2716 40516 2772 40526
rect 2716 40422 2772 40460
rect 2604 40404 2660 40414
rect 2492 40402 2660 40404
rect 2492 40350 2606 40402
rect 2658 40350 2660 40402
rect 2492 40348 2660 40350
rect 2604 40338 2660 40348
rect 2268 40290 2324 40302
rect 2268 40238 2270 40290
rect 2322 40238 2324 40290
rect 2268 39508 2324 40238
rect 2268 39442 2324 39452
rect 2380 40292 2436 40302
rect 2380 39506 2436 40236
rect 2380 39454 2382 39506
rect 2434 39454 2436 39506
rect 2380 39442 2436 39454
rect 2156 38946 2212 38958
rect 2156 38894 2158 38946
rect 2210 38894 2212 38946
rect 2156 38668 2212 38894
rect 2828 38668 2884 41804
rect 2940 41524 2996 41916
rect 2940 41458 2996 41468
rect 3164 41972 3220 41982
rect 2940 41300 2996 41310
rect 2940 41206 2996 41244
rect 3164 40516 3220 41916
rect 3164 40450 3220 40460
rect 3388 40292 3444 42142
rect 3388 40198 3444 40236
rect 2044 38612 2100 38622
rect 2156 38612 2436 38668
rect 2828 38612 2996 38668
rect 2044 38162 2100 38556
rect 2268 38276 2324 38286
rect 2044 38110 2046 38162
rect 2098 38110 2100 38162
rect 2044 38098 2100 38110
rect 2156 38220 2268 38276
rect 2044 37492 2100 37502
rect 2156 37492 2212 38220
rect 2268 38210 2324 38220
rect 2380 38162 2436 38612
rect 2380 38110 2382 38162
rect 2434 38110 2436 38162
rect 2380 38098 2436 38110
rect 2604 37938 2660 37950
rect 2604 37886 2606 37938
rect 2658 37886 2660 37938
rect 2044 37490 2212 37492
rect 2044 37438 2046 37490
rect 2098 37438 2212 37490
rect 2044 37436 2212 37438
rect 2268 37826 2324 37838
rect 2268 37774 2270 37826
rect 2322 37774 2324 37826
rect 2044 37426 2100 37436
rect 2268 36596 2324 37774
rect 2492 37826 2548 37838
rect 2492 37774 2494 37826
rect 2546 37774 2548 37826
rect 2492 37492 2548 37774
rect 2492 37378 2548 37436
rect 2492 37326 2494 37378
rect 2546 37326 2548 37378
rect 2492 37314 2548 37326
rect 2604 37156 2660 37886
rect 2716 37940 2772 37978
rect 2716 37874 2772 37884
rect 2716 37716 2772 37726
rect 2716 37378 2772 37660
rect 2716 37326 2718 37378
rect 2770 37326 2772 37378
rect 2716 37314 2772 37326
rect 2828 37380 2884 37390
rect 2828 37286 2884 37324
rect 2716 37156 2772 37166
rect 2604 37154 2772 37156
rect 2604 37102 2718 37154
rect 2770 37102 2772 37154
rect 2604 37100 2772 37102
rect 2716 37090 2772 37100
rect 2492 36596 2548 36606
rect 2268 36594 2548 36596
rect 2268 36542 2494 36594
rect 2546 36542 2548 36594
rect 2268 36540 2548 36542
rect 2940 36596 2996 38612
rect 3052 38164 3108 38174
rect 3500 38164 3556 42590
rect 3948 42532 4004 43710
rect 4284 43650 4340 43820
rect 4732 43764 4788 44270
rect 4284 43598 4286 43650
rect 4338 43598 4340 43650
rect 4284 43586 4340 43598
rect 4396 43708 4788 43764
rect 4172 43538 4228 43550
rect 4172 43486 4174 43538
rect 4226 43486 4228 43538
rect 4172 43428 4228 43486
rect 4172 43362 4228 43372
rect 4396 43316 4452 43708
rect 4284 43260 4452 43316
rect 4508 43538 4564 43550
rect 4508 43486 4510 43538
rect 4562 43486 4564 43538
rect 4508 43316 4564 43486
rect 4732 43540 4788 43550
rect 4732 43538 4900 43540
rect 4732 43486 4734 43538
rect 4786 43486 4900 43538
rect 4732 43484 4900 43486
rect 4732 43474 4788 43484
rect 4172 42980 4228 42990
rect 4284 42980 4340 43260
rect 4508 43250 4564 43260
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4228 42924 4340 42980
rect 4172 42886 4228 42924
rect 4620 42868 4676 42878
rect 4620 42774 4676 42812
rect 4060 42644 4116 42682
rect 4060 42578 4116 42588
rect 4844 42644 4900 43484
rect 4844 42578 4900 42588
rect 3836 42476 4004 42532
rect 3836 42308 3892 42476
rect 4284 42308 4340 42318
rect 3836 42252 4228 42308
rect 3948 42084 4004 42094
rect 3948 41990 4004 42028
rect 3612 41972 3668 41982
rect 3836 41972 3892 41982
rect 3612 41970 3892 41972
rect 3612 41918 3614 41970
rect 3666 41918 3838 41970
rect 3890 41918 3892 41970
rect 3612 41916 3892 41918
rect 3612 41906 3668 41916
rect 3836 41906 3892 41916
rect 3948 41746 4004 41758
rect 3948 41694 3950 41746
rect 4002 41694 4004 41746
rect 3948 41300 4004 41694
rect 3948 41234 4004 41244
rect 3724 40684 4116 40740
rect 3724 40626 3780 40684
rect 3724 40574 3726 40626
rect 3778 40574 3780 40626
rect 3724 40562 3780 40574
rect 3836 40516 3892 40526
rect 3724 39396 3780 39406
rect 3612 38164 3668 38174
rect 3500 38162 3668 38164
rect 3500 38110 3614 38162
rect 3666 38110 3668 38162
rect 3500 38108 3668 38110
rect 3052 37490 3108 38108
rect 3612 38098 3668 38108
rect 3724 38050 3780 39340
rect 3836 39058 3892 40460
rect 3836 39006 3838 39058
rect 3890 39006 3892 39058
rect 3836 38994 3892 39006
rect 3724 37998 3726 38050
rect 3778 37998 3780 38050
rect 3724 37986 3780 37998
rect 4060 38834 4116 40684
rect 4172 39732 4228 42252
rect 4172 39638 4228 39676
rect 4284 39508 4340 42252
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4060 38782 4062 38834
rect 4114 38782 4116 38834
rect 3388 37938 3444 37950
rect 3388 37886 3390 37938
rect 3442 37886 3444 37938
rect 3388 37716 3444 37886
rect 3388 37650 3444 37660
rect 3052 37438 3054 37490
rect 3106 37438 3108 37490
rect 3052 37426 3108 37438
rect 3276 37492 3332 37502
rect 4060 37492 4116 38782
rect 3052 36596 3108 36606
rect 2940 36540 3052 36596
rect 2492 36530 2548 36540
rect 3052 36530 3108 36540
rect 2156 36484 2212 36494
rect 2156 36372 2212 36428
rect 2828 36484 2884 36494
rect 2884 36428 2996 36484
rect 2828 36418 2884 36428
rect 1708 35970 1764 35980
rect 2044 36370 2212 36372
rect 2044 36318 2158 36370
rect 2210 36318 2212 36370
rect 2044 36316 2212 36318
rect 2044 35922 2100 36316
rect 2156 36306 2212 36316
rect 2940 36370 2996 36428
rect 3276 36482 3332 37436
rect 3276 36430 3278 36482
rect 3330 36430 3332 36482
rect 3276 36418 3332 36430
rect 3500 37436 4116 37492
rect 4172 39452 4340 39508
rect 4396 39618 4452 39630
rect 4396 39566 4398 39618
rect 4450 39566 4452 39618
rect 3500 37154 3556 37436
rect 3500 37102 3502 37154
rect 3554 37102 3556 37154
rect 2940 36318 2942 36370
rect 2994 36318 2996 36370
rect 2940 36306 2996 36318
rect 2044 35870 2046 35922
rect 2098 35870 2100 35922
rect 2044 35858 2100 35870
rect 2380 36260 2436 36270
rect 2380 35812 2436 36204
rect 2604 36260 2660 36270
rect 2604 36166 2660 36204
rect 2268 35810 2436 35812
rect 2268 35758 2382 35810
rect 2434 35758 2436 35810
rect 2268 35756 2436 35758
rect 1932 35700 1988 35710
rect 1932 35698 2100 35700
rect 1932 35646 1934 35698
rect 1986 35646 2100 35698
rect 1932 35644 2100 35646
rect 1932 35634 1988 35644
rect 1372 33842 1428 33852
rect 1932 34690 1988 34702
rect 1932 34638 1934 34690
rect 1986 34638 1988 34690
rect 1932 34468 1988 34638
rect 1932 33796 1988 34412
rect 2044 34020 2100 35644
rect 2156 35698 2212 35710
rect 2156 35646 2158 35698
rect 2210 35646 2212 35698
rect 2156 35028 2212 35646
rect 2156 34962 2212 34972
rect 2156 34580 2212 34590
rect 2156 34130 2212 34524
rect 2156 34078 2158 34130
rect 2210 34078 2212 34130
rect 2156 34066 2212 34078
rect 2044 33954 2100 33964
rect 1708 33740 1988 33796
rect 1708 33124 1764 33740
rect 1932 33572 1988 33582
rect 1932 33478 1988 33516
rect 2156 33572 2212 33582
rect 2268 33572 2324 35756
rect 2380 35746 2436 35756
rect 3388 35810 3444 35822
rect 3388 35758 3390 35810
rect 3442 35758 3444 35810
rect 3052 35476 3108 35486
rect 3388 35476 3444 35758
rect 3500 35698 3556 37102
rect 3500 35646 3502 35698
rect 3554 35646 3556 35698
rect 3500 35634 3556 35646
rect 3612 37266 3668 37278
rect 3612 37214 3614 37266
rect 3666 37214 3668 37266
rect 3612 37044 3668 37214
rect 3612 35476 3668 36988
rect 4172 36706 4228 39452
rect 4396 39396 4452 39566
rect 4396 38836 4452 39340
rect 4732 39396 4788 39406
rect 4732 39302 4788 39340
rect 4732 38948 4788 38958
rect 4732 38854 4788 38892
rect 4396 38770 4452 38780
rect 4508 38834 4564 38846
rect 4508 38782 4510 38834
rect 4562 38782 4564 38834
rect 4172 36654 4174 36706
rect 4226 36654 4228 36706
rect 4172 36642 4228 36654
rect 4284 38722 4340 38734
rect 4284 38670 4286 38722
rect 4338 38670 4340 38722
rect 3388 35420 3668 35476
rect 3948 36594 4004 36606
rect 3948 36542 3950 36594
rect 4002 36542 4004 36594
rect 3948 36260 4004 36542
rect 3052 35138 3108 35420
rect 3052 35086 3054 35138
rect 3106 35086 3108 35138
rect 3052 35074 3108 35086
rect 2492 34916 2548 34926
rect 2380 34802 2436 34814
rect 2380 34750 2382 34802
rect 2434 34750 2436 34802
rect 2380 34356 2436 34750
rect 2380 34290 2436 34300
rect 2492 34354 2548 34860
rect 2492 34302 2494 34354
rect 2546 34302 2548 34354
rect 2492 34290 2548 34302
rect 2604 34914 2660 34926
rect 2604 34862 2606 34914
rect 2658 34862 2660 34914
rect 2604 34804 2660 34862
rect 2212 33516 2324 33572
rect 2380 34130 2436 34142
rect 2380 34078 2382 34130
rect 2434 34078 2436 34130
rect 2156 33506 2212 33516
rect 2156 33124 2212 33134
rect 1708 33068 1988 33124
rect 1820 32676 1876 32686
rect 1708 32620 1820 32676
rect 1708 31220 1764 32620
rect 1820 32610 1876 32620
rect 1820 32452 1876 32462
rect 1820 31332 1876 32396
rect 1932 31890 1988 33068
rect 1932 31838 1934 31890
rect 1986 31838 1988 31890
rect 1932 31826 1988 31838
rect 2044 32562 2100 32574
rect 2044 32510 2046 32562
rect 2098 32510 2100 32562
rect 2044 31556 2100 32510
rect 2156 32228 2212 33068
rect 2380 33124 2436 34078
rect 2380 33058 2436 33068
rect 2492 34020 2548 34030
rect 2492 32900 2548 33964
rect 2268 32844 2548 32900
rect 2268 32676 2324 32844
rect 2268 32450 2324 32620
rect 2492 32676 2548 32686
rect 2268 32398 2270 32450
rect 2322 32398 2324 32450
rect 2268 32386 2324 32398
rect 2380 32562 2436 32574
rect 2380 32510 2382 32562
rect 2434 32510 2436 32562
rect 2380 32452 2436 32510
rect 2380 32386 2436 32396
rect 2156 32172 2436 32228
rect 2156 31780 2212 31818
rect 2156 31714 2212 31724
rect 2380 31778 2436 32172
rect 2380 31726 2382 31778
rect 2434 31726 2436 31778
rect 2380 31714 2436 31726
rect 2044 31500 2436 31556
rect 1820 31276 2324 31332
rect 1708 31164 2100 31220
rect 2044 31106 2100 31164
rect 2268 31218 2324 31276
rect 2268 31166 2270 31218
rect 2322 31166 2324 31218
rect 2268 31154 2324 31166
rect 2044 31054 2046 31106
rect 2098 31054 2100 31106
rect 2044 31042 2100 31054
rect 2156 31108 2212 31118
rect 2156 31014 2212 31052
rect 1260 28018 1316 28028
rect 1596 30996 1652 31006
rect 1148 16146 1204 16156
rect 1260 27636 1316 27646
rect 1260 15540 1316 27580
rect 1596 26852 1652 30940
rect 2268 30098 2324 30110
rect 2268 30046 2270 30098
rect 2322 30046 2324 30098
rect 2044 29652 2100 29662
rect 1708 29314 1764 29326
rect 1708 29262 1710 29314
rect 1762 29262 1764 29314
rect 1708 28868 1764 29262
rect 1708 28754 1764 28812
rect 1708 28702 1710 28754
rect 1762 28702 1764 28754
rect 1708 28690 1764 28702
rect 1932 28756 1988 28766
rect 1820 28644 1876 28654
rect 1820 28550 1876 28588
rect 1932 27972 1988 28700
rect 1932 27858 1988 27916
rect 1932 27806 1934 27858
rect 1986 27806 1988 27858
rect 1932 27794 1988 27806
rect 1932 27188 1988 27198
rect 1932 27074 1988 27132
rect 1932 27022 1934 27074
rect 1986 27022 1988 27074
rect 1932 27010 1988 27022
rect 1596 26796 1764 26852
rect 1708 26404 1764 26796
rect 2044 26514 2100 29596
rect 2268 28868 2324 30046
rect 2268 28802 2324 28812
rect 2380 28866 2436 31500
rect 2380 28814 2382 28866
rect 2434 28814 2436 28866
rect 2380 28756 2436 28814
rect 2380 28690 2436 28700
rect 2492 31218 2548 32620
rect 2492 31166 2494 31218
rect 2546 31166 2548 31218
rect 2268 28420 2324 28430
rect 2268 28082 2324 28364
rect 2492 28196 2548 31166
rect 2604 28420 2660 34748
rect 3612 34804 3668 34814
rect 3388 34692 3444 34702
rect 3388 34690 3556 34692
rect 3388 34638 3390 34690
rect 3442 34638 3556 34690
rect 3388 34636 3556 34638
rect 3388 34626 3444 34636
rect 2940 34356 2996 34366
rect 2716 34132 2772 34142
rect 2940 34132 2996 34300
rect 3388 34244 3444 34254
rect 3388 34150 3444 34188
rect 3164 34132 3220 34142
rect 2716 34130 2884 34132
rect 2716 34078 2718 34130
rect 2770 34078 2884 34130
rect 2716 34076 2884 34078
rect 2716 34066 2772 34076
rect 2716 33572 2772 33582
rect 2716 32002 2772 33516
rect 2716 31950 2718 32002
rect 2770 31950 2772 32002
rect 2716 31938 2772 31950
rect 2828 32004 2884 34076
rect 2940 34130 3220 34132
rect 2940 34078 3166 34130
rect 3218 34078 3220 34130
rect 2940 34076 3220 34078
rect 2940 32452 2996 34076
rect 3164 34066 3220 34076
rect 3052 32676 3108 32686
rect 3052 32674 3332 32676
rect 3052 32622 3054 32674
rect 3106 32622 3332 32674
rect 3052 32620 3332 32622
rect 3052 32610 3108 32620
rect 2940 32396 3108 32452
rect 2828 31938 2884 31948
rect 2940 31892 2996 31902
rect 2604 28354 2660 28364
rect 2716 31778 2772 31790
rect 2716 31726 2718 31778
rect 2770 31726 2772 31778
rect 2716 30996 2772 31726
rect 2492 28140 2660 28196
rect 2268 28030 2270 28082
rect 2322 28030 2324 28082
rect 2268 28018 2324 28030
rect 2268 27860 2324 27870
rect 2156 26964 2212 26974
rect 2268 26964 2324 27804
rect 2604 27858 2660 28140
rect 2604 27806 2606 27858
rect 2658 27806 2660 27858
rect 2604 27794 2660 27806
rect 2716 27524 2772 30940
rect 2604 27468 2772 27524
rect 2828 31780 2884 31790
rect 2828 31332 2884 31724
rect 2940 31554 2996 31836
rect 2940 31502 2942 31554
rect 2994 31502 2996 31554
rect 2940 31490 2996 31502
rect 3052 31332 3108 32396
rect 2828 31276 3108 31332
rect 3164 32116 3220 32126
rect 2604 27186 2660 27468
rect 2604 27134 2606 27186
rect 2658 27134 2660 27186
rect 2604 27122 2660 27134
rect 2716 27188 2772 27198
rect 2156 26962 2324 26964
rect 2156 26910 2158 26962
rect 2210 26910 2324 26962
rect 2156 26908 2324 26910
rect 2156 26898 2212 26908
rect 2044 26462 2046 26514
rect 2098 26462 2100 26514
rect 2044 26450 2100 26462
rect 2156 26404 2212 26414
rect 1708 26402 1876 26404
rect 1708 26350 1710 26402
rect 1762 26350 1876 26402
rect 1708 26348 1876 26350
rect 1708 26338 1764 26348
rect 1708 24948 1764 24958
rect 1372 24612 1428 24622
rect 1372 16772 1428 24556
rect 1484 23828 1540 23838
rect 1484 18452 1540 23772
rect 1708 23266 1764 24892
rect 1708 23214 1710 23266
rect 1762 23214 1764 23266
rect 1708 22820 1764 23214
rect 1820 23156 1876 26348
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 2044 23380 2100 23390
rect 2044 23286 2100 23324
rect 1820 23100 2100 23156
rect 1708 22754 1764 22764
rect 1708 22596 1764 22606
rect 1708 22146 1764 22540
rect 1708 22094 1710 22146
rect 1762 22094 1764 22146
rect 1708 22082 1764 22094
rect 1708 21924 1764 21934
rect 1708 20018 1764 21868
rect 1820 21812 1876 21822
rect 1820 20802 1876 21756
rect 1820 20750 1822 20802
rect 1874 20750 1876 20802
rect 1820 20738 1876 20750
rect 1932 20578 1988 20590
rect 1932 20526 1934 20578
rect 1986 20526 1988 20578
rect 1932 20132 1988 20526
rect 1932 20066 1988 20076
rect 1708 19966 1710 20018
rect 1762 19966 1764 20018
rect 1708 19954 1764 19966
rect 2044 19236 2100 23100
rect 2156 21924 2212 26348
rect 2156 21858 2212 21868
rect 2156 20578 2212 20590
rect 2156 20526 2158 20578
rect 2210 20526 2212 20578
rect 2156 20356 2212 20526
rect 2156 20290 2212 20300
rect 2268 20188 2324 26908
rect 2380 25396 2436 25406
rect 2380 23826 2436 25340
rect 2604 25060 2660 25070
rect 2380 23774 2382 23826
rect 2434 23774 2436 23826
rect 2380 23762 2436 23774
rect 2492 24948 2548 24958
rect 2380 21812 2436 21822
rect 2492 21812 2548 24892
rect 2604 24164 2660 25004
rect 2716 24276 2772 27132
rect 2828 24500 2884 31276
rect 3164 30994 3220 32060
rect 3276 31892 3332 32620
rect 3500 32116 3556 34636
rect 3612 34244 3668 34748
rect 3612 34178 3668 34188
rect 3612 32676 3668 32686
rect 3612 32562 3668 32620
rect 3612 32510 3614 32562
rect 3666 32510 3668 32562
rect 3612 32498 3668 32510
rect 3500 32002 3556 32060
rect 3500 31950 3502 32002
rect 3554 31950 3556 32002
rect 3500 31938 3556 31950
rect 3724 31892 3780 31902
rect 3276 31836 3444 31892
rect 3276 31668 3332 31678
rect 3276 31574 3332 31612
rect 3164 30942 3166 30994
rect 3218 30942 3220 30994
rect 3164 30930 3220 30942
rect 3052 29988 3108 29998
rect 2940 28084 2996 28094
rect 2940 26628 2996 28028
rect 3052 27074 3108 29932
rect 3164 29316 3220 29326
rect 3164 28082 3220 29260
rect 3164 28030 3166 28082
rect 3218 28030 3220 28082
rect 3164 28018 3220 28030
rect 3388 28196 3444 31836
rect 3724 31890 3892 31892
rect 3724 31838 3726 31890
rect 3778 31838 3892 31890
rect 3724 31836 3892 31838
rect 3724 31826 3780 31836
rect 3724 30996 3780 31006
rect 3724 30902 3780 30940
rect 3836 30882 3892 31836
rect 3948 31780 4004 36204
rect 4284 35812 4340 38670
rect 4508 38668 4564 38782
rect 4508 38612 4900 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4732 38050 4788 38062
rect 4732 37998 4734 38050
rect 4786 37998 4788 38050
rect 4732 37604 4788 37998
rect 4844 37828 4900 38612
rect 4956 38164 5012 47068
rect 5292 46900 5348 46910
rect 5180 45890 5236 45902
rect 5180 45838 5182 45890
rect 5234 45838 5236 45890
rect 5180 43650 5236 45838
rect 5292 45106 5348 46844
rect 5292 45054 5294 45106
rect 5346 45054 5348 45106
rect 5292 45042 5348 45054
rect 5180 43598 5182 43650
rect 5234 43598 5236 43650
rect 5180 43586 5236 43598
rect 5404 43428 5460 47292
rect 5628 47236 5684 47246
rect 5516 44548 5572 44558
rect 5516 43538 5572 44492
rect 5516 43486 5518 43538
rect 5570 43486 5572 43538
rect 5516 43474 5572 43486
rect 5180 43372 5460 43428
rect 5068 42530 5124 42542
rect 5068 42478 5070 42530
rect 5122 42478 5124 42530
rect 5068 41972 5124 42478
rect 5068 41906 5124 41916
rect 5180 42194 5236 43372
rect 5628 42754 5684 47180
rect 6076 46674 6132 48636
rect 6188 46788 6244 48750
rect 6300 48468 6356 50652
rect 6412 50036 6468 50046
rect 6524 50036 6580 51660
rect 6860 51604 6916 52222
rect 7868 52386 7924 52398
rect 7868 52334 7870 52386
rect 7922 52334 7924 52386
rect 7420 52164 7476 52174
rect 7420 52070 7476 52108
rect 7196 51940 7252 51950
rect 6916 51548 7028 51604
rect 6860 51538 6916 51548
rect 6860 51268 6916 51278
rect 6860 51174 6916 51212
rect 6860 50596 6916 50606
rect 6636 50540 6804 50596
rect 6636 50482 6692 50540
rect 6636 50430 6638 50482
rect 6690 50430 6692 50482
rect 6636 50418 6692 50430
rect 6748 50372 6804 50540
rect 6412 50034 6580 50036
rect 6412 49982 6414 50034
rect 6466 49982 6580 50034
rect 6412 49980 6580 49982
rect 6636 50036 6692 50046
rect 6412 49970 6468 49980
rect 6636 48804 6692 49980
rect 6748 50034 6804 50316
rect 6748 49982 6750 50034
rect 6802 49982 6804 50034
rect 6748 49970 6804 49982
rect 6860 49138 6916 50540
rect 6860 49086 6862 49138
rect 6914 49086 6916 49138
rect 6860 49074 6916 49086
rect 6972 49028 7028 51548
rect 7196 51602 7252 51884
rect 7196 51550 7198 51602
rect 7250 51550 7252 51602
rect 7084 50596 7140 50634
rect 7084 50530 7140 50540
rect 7196 50428 7252 51550
rect 7868 51938 7924 52334
rect 7868 51886 7870 51938
rect 7922 51886 7924 51938
rect 7084 50372 7252 50428
rect 7644 51268 7700 51278
rect 7868 51268 7924 51886
rect 7644 51266 7924 51268
rect 7644 51214 7646 51266
rect 7698 51214 7924 51266
rect 7644 51212 7924 51214
rect 7084 50036 7140 50372
rect 7532 50370 7588 50382
rect 7532 50318 7534 50370
rect 7586 50318 7588 50370
rect 7084 49970 7140 49980
rect 7308 50036 7364 50046
rect 7308 49942 7364 49980
rect 7196 49028 7252 49038
rect 6972 49026 7252 49028
rect 6972 48974 7198 49026
rect 7250 48974 7252 49026
rect 6972 48972 7252 48974
rect 6636 48748 7028 48804
rect 6300 48412 6468 48468
rect 6188 46722 6244 46732
rect 6300 48242 6356 48254
rect 6300 48190 6302 48242
rect 6354 48190 6356 48242
rect 6076 46622 6078 46674
rect 6130 46622 6132 46674
rect 5740 46004 5796 46014
rect 5740 45910 5796 45948
rect 6076 45890 6132 46622
rect 6076 45838 6078 45890
rect 6130 45838 6132 45890
rect 6076 45826 6132 45838
rect 6300 46562 6356 48190
rect 6300 46510 6302 46562
rect 6354 46510 6356 46562
rect 6300 45892 6356 46510
rect 6300 45826 6356 45836
rect 5964 45108 6020 45118
rect 5740 44994 5796 45006
rect 5740 44942 5742 44994
rect 5794 44942 5796 44994
rect 5740 44884 5796 44942
rect 5740 44818 5796 44828
rect 5740 44436 5796 44446
rect 5740 44342 5796 44380
rect 5964 44210 6020 45052
rect 6300 45106 6356 45118
rect 6300 45054 6302 45106
rect 6354 45054 6356 45106
rect 6076 44548 6132 44558
rect 6076 44322 6132 44492
rect 6300 44436 6356 45054
rect 6300 44370 6356 44380
rect 6076 44270 6078 44322
rect 6130 44270 6132 44322
rect 6076 44258 6132 44270
rect 5964 44158 5966 44210
rect 6018 44158 6020 44210
rect 5964 43538 6020 44158
rect 5964 43486 5966 43538
rect 6018 43486 6020 43538
rect 5964 43474 6020 43486
rect 6300 43650 6356 43662
rect 6300 43598 6302 43650
rect 6354 43598 6356 43650
rect 6300 43316 6356 43598
rect 6412 43652 6468 48412
rect 6748 48242 6804 48254
rect 6748 48190 6750 48242
rect 6802 48190 6804 48242
rect 6524 47348 6580 47358
rect 6524 47254 6580 47292
rect 6636 46786 6692 46798
rect 6636 46734 6638 46786
rect 6690 46734 6692 46786
rect 6636 45220 6692 46734
rect 6748 46004 6804 48190
rect 6860 46788 6916 46798
rect 6860 46694 6916 46732
rect 6804 45948 6916 46004
rect 6748 45938 6804 45948
rect 6748 45780 6804 45790
rect 6748 45686 6804 45724
rect 6636 45126 6692 45164
rect 6524 45108 6580 45118
rect 6524 44994 6580 45052
rect 6524 44942 6526 44994
rect 6578 44942 6580 44994
rect 6524 44930 6580 44942
rect 6860 44322 6916 45948
rect 6860 44270 6862 44322
rect 6914 44270 6916 44322
rect 6860 44258 6916 44270
rect 6972 43876 7028 48748
rect 7084 48132 7140 48972
rect 7196 48962 7252 48972
rect 7532 48356 7588 50318
rect 7532 48290 7588 48300
rect 7084 48066 7140 48076
rect 7420 47460 7476 47470
rect 7308 46900 7364 46910
rect 7308 46674 7364 46844
rect 7308 46622 7310 46674
rect 7362 46622 7364 46674
rect 7196 45780 7252 45790
rect 7308 45780 7364 46622
rect 7196 45778 7364 45780
rect 7196 45726 7198 45778
rect 7250 45726 7364 45778
rect 7196 45724 7364 45726
rect 7420 46114 7476 47404
rect 7420 46062 7422 46114
rect 7474 46062 7476 46114
rect 7196 45714 7252 45724
rect 7420 45556 7476 46062
rect 7644 45780 7700 51212
rect 7868 50708 7924 50718
rect 7868 50614 7924 50652
rect 7980 50428 8036 52780
rect 8092 52770 8148 52780
rect 8316 52724 8372 52734
rect 8204 52668 8316 52724
rect 8204 52164 8260 52668
rect 8316 52658 8372 52668
rect 8316 52386 8372 52398
rect 8316 52334 8318 52386
rect 8370 52334 8372 52386
rect 8316 52274 8372 52334
rect 8316 52222 8318 52274
rect 8370 52222 8372 52274
rect 8316 52210 8372 52222
rect 7868 50372 8036 50428
rect 8092 52108 8260 52164
rect 8092 50708 8148 52108
rect 8204 51604 8260 51614
rect 8428 51604 8484 53228
rect 8540 53218 8596 53228
rect 9100 53172 9156 53182
rect 9100 53078 9156 53116
rect 8204 51602 8484 51604
rect 8204 51550 8206 51602
rect 8258 51550 8484 51602
rect 8204 51548 8484 51550
rect 8540 52834 8596 52846
rect 8540 52782 8542 52834
rect 8594 52782 8596 52834
rect 8204 51538 8260 51548
rect 7756 49700 7812 49710
rect 7756 49606 7812 49644
rect 7084 45500 7476 45556
rect 7532 45724 7700 45780
rect 7084 45330 7140 45500
rect 7084 45278 7086 45330
rect 7138 45278 7140 45330
rect 7084 44884 7140 45278
rect 7308 45332 7364 45342
rect 7308 45238 7364 45276
rect 7420 45220 7476 45230
rect 7420 45126 7476 45164
rect 7084 44818 7140 44828
rect 7308 44994 7364 45006
rect 7308 44942 7310 44994
rect 7362 44942 7364 44994
rect 7196 44324 7252 44334
rect 7196 44230 7252 44268
rect 6972 43820 7252 43876
rect 7084 43652 7140 43662
rect 6468 43596 6580 43652
rect 6412 43586 6468 43596
rect 6300 43250 6356 43260
rect 5628 42702 5630 42754
rect 5682 42702 5684 42754
rect 5628 42690 5684 42702
rect 5740 42868 5796 42878
rect 5740 42642 5796 42812
rect 5964 42756 6020 42766
rect 5964 42662 6020 42700
rect 5740 42590 5742 42642
rect 5794 42590 5796 42642
rect 5740 42578 5796 42590
rect 6300 42642 6356 42654
rect 6300 42590 6302 42642
rect 6354 42590 6356 42642
rect 6188 42532 6244 42542
rect 5180 42142 5182 42194
rect 5234 42142 5236 42194
rect 5068 41300 5124 41310
rect 5180 41300 5236 42142
rect 5740 42420 5796 42430
rect 5068 41298 5236 41300
rect 5068 41246 5070 41298
rect 5122 41246 5236 41298
rect 5068 41244 5236 41246
rect 5068 41234 5124 41244
rect 5180 40626 5236 41244
rect 5180 40574 5182 40626
rect 5234 40574 5236 40626
rect 5180 40562 5236 40574
rect 5516 41860 5572 41870
rect 5292 39396 5348 39406
rect 5068 38948 5124 38958
rect 5068 38668 5124 38892
rect 5068 38612 5236 38668
rect 4956 38070 5012 38108
rect 4844 37762 4900 37772
rect 5068 37604 5124 37614
rect 4732 37548 5068 37604
rect 4732 37380 4788 37548
rect 5068 37538 5124 37548
rect 4732 37314 4788 37324
rect 5068 36932 5124 36942
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 5068 36594 5124 36876
rect 5068 36542 5070 36594
rect 5122 36542 5124 36594
rect 5068 36530 5124 36542
rect 4396 36482 4452 36494
rect 4396 36430 4398 36482
rect 4450 36430 4452 36482
rect 4396 36372 4452 36430
rect 4396 36306 4452 36316
rect 4284 35746 4340 35756
rect 4732 35700 4788 35710
rect 5180 35700 5236 38612
rect 5292 37266 5348 39340
rect 5404 38836 5460 38846
rect 5404 38742 5460 38780
rect 5292 37214 5294 37266
rect 5346 37214 5348 37266
rect 5292 37202 5348 37214
rect 5516 36932 5572 41804
rect 5740 41298 5796 42364
rect 5740 41246 5742 41298
rect 5794 41246 5796 41298
rect 5740 41234 5796 41246
rect 6188 41186 6244 42476
rect 6300 42420 6356 42590
rect 6300 42354 6356 42364
rect 6300 41972 6356 41982
rect 6300 41878 6356 41916
rect 6524 41298 6580 43596
rect 6636 43540 6692 43550
rect 6636 42754 6692 43484
rect 6636 42702 6638 42754
rect 6690 42702 6692 42754
rect 6636 42690 6692 42702
rect 6972 43538 7028 43550
rect 6972 43486 6974 43538
rect 7026 43486 7028 43538
rect 6972 42308 7028 43486
rect 7084 43428 7140 43596
rect 7084 42754 7140 43372
rect 7196 43204 7252 43820
rect 7196 43138 7252 43148
rect 7084 42702 7086 42754
rect 7138 42702 7140 42754
rect 7084 42690 7140 42702
rect 7196 42530 7252 42542
rect 7196 42478 7198 42530
rect 7250 42478 7252 42530
rect 6972 42252 7140 42308
rect 6860 42196 6916 42206
rect 6748 42140 6860 42196
rect 6636 42084 6692 42094
rect 6636 41990 6692 42028
rect 6748 42082 6804 42140
rect 6860 42130 6916 42140
rect 6748 42030 6750 42082
rect 6802 42030 6804 42082
rect 6748 42018 6804 42030
rect 6972 42084 7028 42094
rect 6972 41990 7028 42028
rect 6972 41748 7028 41758
rect 6524 41246 6526 41298
rect 6578 41246 6580 41298
rect 6524 41234 6580 41246
rect 6860 41300 6916 41310
rect 6188 41134 6190 41186
rect 6242 41134 6244 41186
rect 6188 41122 6244 41134
rect 6076 40964 6132 40974
rect 6076 39956 6132 40908
rect 6076 39890 6132 39900
rect 6188 40628 6244 40638
rect 5628 39732 5684 39742
rect 5628 38834 5684 39676
rect 6076 39732 6132 39742
rect 6076 39638 6132 39676
rect 5628 38782 5630 38834
rect 5682 38782 5684 38834
rect 5628 38770 5684 38782
rect 5964 38836 6020 38846
rect 5964 38742 6020 38780
rect 6076 37938 6132 37950
rect 6076 37886 6078 37938
rect 6130 37886 6132 37938
rect 6076 37492 6132 37886
rect 6076 37426 6132 37436
rect 5740 37156 5796 37166
rect 5740 37062 5796 37100
rect 5516 36866 5572 36876
rect 5628 36372 5684 36382
rect 5628 36278 5684 36316
rect 5852 36260 5908 36270
rect 4732 35698 5236 35700
rect 4732 35646 4734 35698
rect 4786 35646 5236 35698
rect 4732 35644 5236 35646
rect 5404 36036 5460 36046
rect 4732 35634 4788 35644
rect 4284 35586 4340 35598
rect 4284 35534 4286 35586
rect 4338 35534 4340 35586
rect 4060 35026 4116 35038
rect 4060 34974 4062 35026
rect 4114 34974 4116 35026
rect 4060 34020 4116 34974
rect 4060 33926 4116 33964
rect 4172 35028 4228 35038
rect 4172 34914 4228 34972
rect 4172 34862 4174 34914
rect 4226 34862 4228 34914
rect 4060 33460 4116 33470
rect 4060 33346 4116 33404
rect 4060 33294 4062 33346
rect 4114 33294 4116 33346
rect 4060 33282 4116 33294
rect 4060 33124 4116 33134
rect 4060 32564 4116 33068
rect 4060 32470 4116 32508
rect 4172 32452 4228 34862
rect 4284 34132 4340 35534
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4508 34916 4564 34926
rect 4508 34914 4676 34916
rect 4508 34862 4510 34914
rect 4562 34862 4676 34914
rect 4508 34860 4676 34862
rect 4508 34850 4564 34860
rect 4620 34356 4676 34860
rect 4732 34690 4788 34702
rect 4732 34638 4734 34690
rect 4786 34638 4788 34690
rect 4732 34580 4788 34638
rect 4844 34580 4900 34590
rect 4732 34524 4844 34580
rect 4844 34514 4900 34524
rect 4620 34300 4900 34356
rect 4732 34132 4788 34142
rect 4284 34130 4788 34132
rect 4284 34078 4734 34130
rect 4786 34078 4788 34130
rect 4284 34076 4788 34078
rect 4284 33572 4340 34076
rect 4732 34066 4788 34076
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4284 33506 4340 33516
rect 4844 32676 4900 34300
rect 4844 32582 4900 32620
rect 4956 33348 5012 33358
rect 4172 32386 4228 32396
rect 4508 32452 4564 32462
rect 4956 32452 5012 33292
rect 4508 32358 4564 32396
rect 4844 32396 5012 32452
rect 5180 33122 5236 33134
rect 5180 33070 5182 33122
rect 5234 33070 5236 33122
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4732 32004 4788 32014
rect 4844 32004 4900 32396
rect 5180 32116 5236 33070
rect 5180 32050 5236 32060
rect 5404 32900 5460 35980
rect 5852 35138 5908 36204
rect 5852 35086 5854 35138
rect 5906 35086 5908 35138
rect 5852 35074 5908 35086
rect 5964 36258 6020 36270
rect 5964 36206 5966 36258
rect 6018 36206 6020 36258
rect 5964 35698 6020 36206
rect 5964 35646 5966 35698
rect 6018 35646 6020 35698
rect 5964 34804 6020 35646
rect 6188 35140 6244 40572
rect 6300 40404 6356 40414
rect 6748 40404 6804 40414
rect 6300 40402 6804 40404
rect 6300 40350 6302 40402
rect 6354 40350 6750 40402
rect 6802 40350 6804 40402
rect 6300 40348 6804 40350
rect 6300 40338 6356 40348
rect 6748 40338 6804 40348
rect 6860 40180 6916 41244
rect 6748 40124 6916 40180
rect 6412 39620 6468 39630
rect 6412 39526 6468 39564
rect 6300 39508 6356 39518
rect 6300 39414 6356 39452
rect 6300 38722 6356 38734
rect 6300 38670 6302 38722
rect 6354 38670 6356 38722
rect 6300 38668 6356 38670
rect 6300 38612 6692 38668
rect 6412 37828 6468 37838
rect 6412 37490 6468 37772
rect 6412 37438 6414 37490
rect 6466 37438 6468 37490
rect 6412 37426 6468 37438
rect 6636 37266 6692 38612
rect 6636 37214 6638 37266
rect 6690 37214 6692 37266
rect 6636 37044 6692 37214
rect 6636 36978 6692 36988
rect 6524 36708 6580 36718
rect 6524 36614 6580 36652
rect 6748 35252 6804 40124
rect 6972 39732 7028 41692
rect 7084 41188 7140 42252
rect 7196 41860 7252 42478
rect 7308 42196 7364 44942
rect 7420 43428 7476 43438
rect 7532 43428 7588 45724
rect 7756 45668 7812 45678
rect 7420 43426 7588 43428
rect 7420 43374 7422 43426
rect 7474 43374 7588 43426
rect 7420 43372 7588 43374
rect 7644 45666 7812 45668
rect 7644 45614 7758 45666
rect 7810 45614 7812 45666
rect 7644 45612 7812 45614
rect 7644 44322 7700 45612
rect 7756 45602 7812 45612
rect 7868 45444 7924 50372
rect 8092 50034 8148 50652
rect 8092 49982 8094 50034
rect 8146 49982 8148 50034
rect 8092 49970 8148 49982
rect 8204 51156 8260 51166
rect 7980 48914 8036 48926
rect 7980 48862 7982 48914
rect 8034 48862 8036 48914
rect 7980 46900 8036 48862
rect 8092 48468 8148 48478
rect 8204 48468 8260 51100
rect 8428 50482 8484 50494
rect 8428 50430 8430 50482
rect 8482 50430 8484 50482
rect 8428 50428 8484 50430
rect 8316 50372 8484 50428
rect 8316 49364 8372 50316
rect 8540 49924 8596 52782
rect 9100 52276 9156 52286
rect 9548 52276 9604 54796
rect 9996 54628 10052 55022
rect 9996 54562 10052 54572
rect 9660 54404 9716 54414
rect 9660 54310 9716 54348
rect 10108 53730 10164 57148
rect 11228 55970 11284 55982
rect 11228 55918 11230 55970
rect 11282 55918 11284 55970
rect 10556 55076 10612 55086
rect 10556 54982 10612 55020
rect 11004 55076 11060 55086
rect 11004 54982 11060 55020
rect 11228 54852 11284 55918
rect 11228 54786 11284 54796
rect 10108 53678 10110 53730
rect 10162 53678 10164 53730
rect 10108 53666 10164 53678
rect 10220 54402 10276 54414
rect 10220 54350 10222 54402
rect 10274 54350 10276 54402
rect 9660 53620 9716 53630
rect 9660 53526 9716 53564
rect 10220 53508 10276 54350
rect 10668 54402 10724 54414
rect 10668 54350 10670 54402
rect 10722 54350 10724 54402
rect 10668 53954 10724 54350
rect 10668 53902 10670 53954
rect 10722 53902 10724 53954
rect 10668 53890 10724 53902
rect 10892 54404 10948 54414
rect 10892 54180 10948 54348
rect 11004 54402 11060 54414
rect 11004 54350 11006 54402
rect 11058 54350 11060 54402
rect 11004 54292 11060 54350
rect 11004 54226 11060 54236
rect 10892 53730 10948 54124
rect 10892 53678 10894 53730
rect 10946 53678 10948 53730
rect 10892 53666 10948 53678
rect 11340 53620 11396 60508
rect 11452 60498 11508 60508
rect 16156 60228 16212 63200
rect 25340 60564 25396 60574
rect 25396 60508 25508 60564
rect 25340 60498 25396 60508
rect 16156 60162 16212 60172
rect 17948 60228 18004 60238
rect 17948 60134 18004 60172
rect 15372 60004 15428 60014
rect 15260 60002 15428 60004
rect 15260 59950 15374 60002
rect 15426 59950 15428 60002
rect 15260 59948 15428 59950
rect 13580 59892 13636 59902
rect 13580 59798 13636 59836
rect 13804 59890 13860 59902
rect 13804 59838 13806 59890
rect 13858 59838 13860 59890
rect 12908 58996 12964 59006
rect 12684 57538 12740 57550
rect 12684 57486 12686 57538
rect 12738 57486 12740 57538
rect 12124 57428 12180 57438
rect 12124 56978 12180 57372
rect 12684 57428 12740 57486
rect 12684 57362 12740 57372
rect 12124 56926 12126 56978
rect 12178 56926 12180 56978
rect 12124 56914 12180 56926
rect 11676 56644 11732 56654
rect 11564 56642 11732 56644
rect 11564 56590 11678 56642
rect 11730 56590 11732 56642
rect 11564 56588 11732 56590
rect 11452 55074 11508 55086
rect 11452 55022 11454 55074
rect 11506 55022 11508 55074
rect 11452 53844 11508 55022
rect 11564 54628 11620 56588
rect 11676 56578 11732 56588
rect 12572 56642 12628 56654
rect 12572 56590 12574 56642
rect 12626 56590 12628 56642
rect 12572 56196 12628 56590
rect 12572 56130 12628 56140
rect 11676 55970 11732 55982
rect 11676 55918 11678 55970
rect 11730 55918 11732 55970
rect 11676 55524 11732 55918
rect 12124 55972 12180 55982
rect 12572 55972 12628 55982
rect 12124 55970 12572 55972
rect 12124 55918 12126 55970
rect 12178 55918 12572 55970
rect 12124 55916 12572 55918
rect 12124 55906 12180 55916
rect 12572 55878 12628 55916
rect 11676 55458 11732 55468
rect 12684 55188 12740 55198
rect 11788 55076 11844 55086
rect 11676 54628 11732 54638
rect 11564 54572 11676 54628
rect 11676 54562 11732 54572
rect 11788 54402 11844 55020
rect 11788 54350 11790 54402
rect 11842 54350 11844 54402
rect 11788 54292 11844 54350
rect 11788 54226 11844 54236
rect 11900 55074 11956 55086
rect 11900 55022 11902 55074
rect 11954 55022 11956 55074
rect 11452 53778 11508 53788
rect 11676 53842 11732 53854
rect 11676 53790 11678 53842
rect 11730 53790 11732 53842
rect 11564 53732 11620 53742
rect 11452 53620 11508 53630
rect 11340 53618 11508 53620
rect 11340 53566 11454 53618
rect 11506 53566 11508 53618
rect 11340 53564 11508 53566
rect 11452 53554 11508 53564
rect 9884 53284 9940 53294
rect 9884 53170 9940 53228
rect 9884 53118 9886 53170
rect 9938 53118 9940 53170
rect 9884 53106 9940 53118
rect 9156 52274 9604 52276
rect 9156 52222 9550 52274
rect 9602 52222 9604 52274
rect 9156 52220 9604 52222
rect 9100 52182 9156 52220
rect 9548 52210 9604 52220
rect 10108 52722 10164 52734
rect 10108 52670 10110 52722
rect 10162 52670 10164 52722
rect 10108 52162 10164 52670
rect 10220 52276 10276 53452
rect 10556 53508 10612 53518
rect 10556 53414 10612 53452
rect 11228 53508 11284 53518
rect 10444 52836 10500 52846
rect 10892 52836 10948 52846
rect 10444 52834 10948 52836
rect 10444 52782 10446 52834
rect 10498 52782 10894 52834
rect 10946 52782 10948 52834
rect 10444 52780 10948 52782
rect 10444 52770 10500 52780
rect 10220 52210 10276 52220
rect 10108 52110 10110 52162
rect 10162 52110 10164 52162
rect 10108 52098 10164 52110
rect 8764 51940 8820 51950
rect 8764 51846 8820 51884
rect 10220 51940 10276 51950
rect 10444 51940 10500 51950
rect 10108 51828 10164 51838
rect 9996 51772 10108 51828
rect 8652 51604 8708 51614
rect 8652 51510 8708 51548
rect 9100 51266 9156 51278
rect 9100 51214 9102 51266
rect 9154 51214 9156 51266
rect 9100 51044 9156 51214
rect 8652 50482 8708 50494
rect 8652 50430 8654 50482
rect 8706 50430 8708 50482
rect 8652 50148 8708 50430
rect 8652 50082 8708 50092
rect 8764 50482 8820 50494
rect 8764 50430 8766 50482
rect 8818 50430 8820 50482
rect 8540 49858 8596 49868
rect 8316 49298 8372 49308
rect 8428 49810 8484 49822
rect 8428 49758 8430 49810
rect 8482 49758 8484 49810
rect 8092 48466 8260 48468
rect 8092 48414 8094 48466
rect 8146 48414 8260 48466
rect 8092 48412 8260 48414
rect 8092 48402 8148 48412
rect 8316 48244 8372 48254
rect 8316 48150 8372 48188
rect 8316 47684 8372 47694
rect 8316 47236 8372 47628
rect 8316 47012 8372 47180
rect 8428 47572 8484 49758
rect 8652 49810 8708 49822
rect 8652 49758 8654 49810
rect 8706 49758 8708 49810
rect 8540 47684 8596 47694
rect 8652 47684 8708 49758
rect 8764 48692 8820 50430
rect 8988 50484 9044 50522
rect 8988 50418 9044 50428
rect 9100 50036 9156 50988
rect 9548 50820 9604 50830
rect 9324 50708 9380 50718
rect 9324 50594 9380 50652
rect 9324 50542 9326 50594
rect 9378 50542 9380 50594
rect 9324 50530 9380 50542
rect 9436 50596 9492 50606
rect 9100 49970 9156 49980
rect 9100 49812 9156 49822
rect 9100 49810 9380 49812
rect 9100 49758 9102 49810
rect 9154 49758 9380 49810
rect 9100 49756 9380 49758
rect 9100 49746 9156 49756
rect 8876 49700 8932 49710
rect 8876 49606 8932 49644
rect 8764 48626 8820 48636
rect 8764 48468 8820 48478
rect 8764 48466 9268 48468
rect 8764 48414 8766 48466
rect 8818 48414 9268 48466
rect 8764 48412 9268 48414
rect 8764 48402 8820 48412
rect 8988 48242 9044 48254
rect 8988 48190 8990 48242
rect 9042 48190 9044 48242
rect 8540 47682 8708 47684
rect 8540 47630 8542 47682
rect 8594 47630 8708 47682
rect 8540 47628 8708 47630
rect 8540 47618 8596 47628
rect 8428 47124 8484 47516
rect 8652 47348 8708 47628
rect 8652 47282 8708 47292
rect 8876 48130 8932 48142
rect 8876 48078 8878 48130
rect 8930 48078 8932 48130
rect 8428 47068 8708 47124
rect 8316 46956 8596 47012
rect 7980 46844 8484 46900
rect 8428 46786 8484 46844
rect 8540 46898 8596 46956
rect 8540 46846 8542 46898
rect 8594 46846 8596 46898
rect 8540 46834 8596 46846
rect 8428 46734 8430 46786
rect 8482 46734 8484 46786
rect 8428 46722 8484 46734
rect 8316 46674 8372 46686
rect 8316 46622 8318 46674
rect 8370 46622 8372 46674
rect 8316 45556 8372 46622
rect 8652 46002 8708 47068
rect 8876 46788 8932 48078
rect 8988 47124 9044 48190
rect 9212 47796 9268 48412
rect 9212 47570 9268 47740
rect 9212 47518 9214 47570
rect 9266 47518 9268 47570
rect 9212 47506 9268 47518
rect 9324 47458 9380 49756
rect 9324 47406 9326 47458
rect 9378 47406 9380 47458
rect 8988 47058 9044 47068
rect 9212 47348 9268 47358
rect 8876 46722 8932 46732
rect 8652 45950 8654 46002
rect 8706 45950 8708 46002
rect 8652 45938 8708 45950
rect 8764 46562 8820 46574
rect 8764 46510 8766 46562
rect 8818 46510 8820 46562
rect 8764 46004 8820 46510
rect 8764 45938 8820 45948
rect 8988 46450 9044 46462
rect 8988 46398 8990 46450
rect 9042 46398 9044 46450
rect 8092 45500 8372 45556
rect 8540 45890 8596 45902
rect 8540 45838 8542 45890
rect 8594 45838 8596 45890
rect 8540 45556 8596 45838
rect 8652 45780 8708 45790
rect 8652 45778 8820 45780
rect 8652 45726 8654 45778
rect 8706 45726 8820 45778
rect 8652 45724 8820 45726
rect 8652 45714 8708 45724
rect 8540 45500 8708 45556
rect 8092 45444 8148 45500
rect 7644 44270 7646 44322
rect 7698 44270 7700 44322
rect 7420 42308 7476 43372
rect 7420 42242 7476 42252
rect 7532 43204 7588 43214
rect 7308 42130 7364 42140
rect 7532 42084 7588 43148
rect 7644 42754 7700 44270
rect 7644 42702 7646 42754
rect 7698 42702 7700 42754
rect 7644 42690 7700 42702
rect 7756 45388 8148 45444
rect 7532 42018 7588 42028
rect 7308 41970 7364 41982
rect 7308 41918 7310 41970
rect 7362 41918 7364 41970
rect 7308 41860 7364 41918
rect 7532 41860 7588 41870
rect 7308 41858 7588 41860
rect 7308 41806 7534 41858
rect 7586 41806 7588 41858
rect 7308 41804 7588 41806
rect 7196 41794 7252 41804
rect 7532 41794 7588 41804
rect 7084 40514 7140 41132
rect 7420 41412 7476 41422
rect 7084 40462 7086 40514
rect 7138 40462 7140 40514
rect 7084 40292 7140 40462
rect 7084 40226 7140 40236
rect 7196 40740 7252 40750
rect 6972 39666 7028 39676
rect 6860 39620 6916 39630
rect 6860 39526 6916 39564
rect 6748 35186 6804 35196
rect 6972 38946 7028 38958
rect 6972 38894 6974 38946
rect 7026 38894 7028 38946
rect 6188 35084 6468 35140
rect 6188 34916 6244 34926
rect 6188 34822 6244 34860
rect 5964 34738 6020 34748
rect 6300 34804 6356 34814
rect 5628 34580 5684 34590
rect 5628 33346 5684 34524
rect 6076 34130 6132 34142
rect 6076 34078 6078 34130
rect 6130 34078 6132 34130
rect 5628 33294 5630 33346
rect 5682 33294 5684 33346
rect 5628 33282 5684 33294
rect 5964 33572 6020 33582
rect 5068 32004 5124 32014
rect 4788 31948 4900 32004
rect 4956 31948 5068 32004
rect 4732 31890 4788 31948
rect 4732 31838 4734 31890
rect 4786 31838 4788 31890
rect 4732 31826 4788 31838
rect 3948 31714 4004 31724
rect 4284 31780 4340 31790
rect 3836 30830 3838 30882
rect 3890 30830 3892 30882
rect 3836 30212 3892 30830
rect 3836 30146 3892 30156
rect 3948 31556 4004 31566
rect 3500 29988 3556 29998
rect 3500 29894 3556 29932
rect 3836 29540 3892 29550
rect 3948 29540 4004 31500
rect 3836 29538 4004 29540
rect 3836 29486 3838 29538
rect 3890 29486 4004 29538
rect 3836 29484 4004 29486
rect 3836 29474 3892 29484
rect 3052 27022 3054 27074
rect 3106 27022 3108 27074
rect 3052 27010 3108 27022
rect 3388 27074 3444 28140
rect 3388 27022 3390 27074
rect 3442 27022 3444 27074
rect 3388 27010 3444 27022
rect 3500 29204 3556 29214
rect 3500 27970 3556 29148
rect 4284 28084 4340 31724
rect 4844 31778 4900 31790
rect 4844 31726 4846 31778
rect 4898 31726 4900 31778
rect 4844 31332 4900 31726
rect 4844 31266 4900 31276
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4956 30434 5012 31948
rect 5068 31938 5124 31948
rect 4956 30382 4958 30434
rect 5010 30382 5012 30434
rect 4956 30370 5012 30382
rect 4620 30322 4676 30334
rect 4620 30270 4622 30322
rect 4674 30270 4676 30322
rect 4508 29426 4564 29438
rect 4508 29374 4510 29426
rect 4562 29374 4564 29426
rect 4508 29204 4564 29374
rect 4620 29316 4676 30270
rect 4732 30210 4788 30222
rect 4732 30158 4734 30210
rect 4786 30158 4788 30210
rect 4732 30100 4788 30158
rect 4732 29652 4788 30044
rect 4732 29586 4788 29596
rect 4620 29250 4676 29260
rect 4508 29138 4564 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4396 28868 4452 28878
rect 4396 28530 4452 28812
rect 4396 28478 4398 28530
rect 4450 28478 4452 28530
rect 4396 28466 4452 28478
rect 5404 28308 5460 32844
rect 5852 32676 5908 32686
rect 5852 32564 5908 32620
rect 5628 32562 5908 32564
rect 5628 32510 5854 32562
rect 5906 32510 5908 32562
rect 5628 32508 5908 32510
rect 5516 31780 5572 31790
rect 5516 31108 5572 31724
rect 5628 31778 5684 32508
rect 5852 32498 5908 32508
rect 5964 32564 6020 33516
rect 5628 31726 5630 31778
rect 5682 31726 5684 31778
rect 5628 31714 5684 31726
rect 5964 31778 6020 32508
rect 5964 31726 5966 31778
rect 6018 31726 6020 31778
rect 5964 31714 6020 31726
rect 6076 31780 6132 34078
rect 6188 33348 6244 33358
rect 6300 33348 6356 34748
rect 6412 34020 6468 35084
rect 6748 35028 6804 35038
rect 6748 34802 6804 34972
rect 6748 34750 6750 34802
rect 6802 34750 6804 34802
rect 6748 34738 6804 34750
rect 6860 34914 6916 34926
rect 6860 34862 6862 34914
rect 6914 34862 6916 34914
rect 6860 34804 6916 34862
rect 6860 34738 6916 34748
rect 6860 34132 6916 34142
rect 6412 33954 6468 33964
rect 6636 34130 6916 34132
rect 6636 34078 6862 34130
rect 6914 34078 6916 34130
rect 6636 34076 6916 34078
rect 6188 33346 6356 33348
rect 6188 33294 6190 33346
rect 6242 33294 6356 33346
rect 6188 33292 6356 33294
rect 6188 33282 6244 33292
rect 6524 32676 6580 32686
rect 6188 32562 6244 32574
rect 6188 32510 6190 32562
rect 6242 32510 6244 32562
rect 6188 32004 6244 32510
rect 6188 31938 6244 31948
rect 6188 31780 6244 31790
rect 6076 31778 6244 31780
rect 6076 31726 6190 31778
rect 6242 31726 6244 31778
rect 6076 31724 6244 31726
rect 6188 31668 6244 31724
rect 6188 31444 6244 31612
rect 6412 31780 6468 31790
rect 6412 31554 6468 31724
rect 6412 31502 6414 31554
rect 6466 31502 6468 31554
rect 6412 31490 6468 31502
rect 6188 31378 6244 31388
rect 5628 31108 5684 31118
rect 5516 31106 5684 31108
rect 5516 31054 5630 31106
rect 5682 31054 5684 31106
rect 5516 31052 5684 31054
rect 5628 31042 5684 31052
rect 5852 30996 5908 31006
rect 5628 30324 5684 30334
rect 5516 29538 5572 29550
rect 5516 29486 5518 29538
rect 5570 29486 5572 29538
rect 5516 28868 5572 29486
rect 5516 28802 5572 28812
rect 5628 28644 5684 30268
rect 5740 30212 5796 30222
rect 5740 30118 5796 30156
rect 5628 28530 5684 28588
rect 5628 28478 5630 28530
rect 5682 28478 5684 28530
rect 5628 28466 5684 28478
rect 5740 28532 5796 28542
rect 5852 28532 5908 30940
rect 5964 30994 6020 31006
rect 5964 30942 5966 30994
rect 6018 30942 6020 30994
rect 5964 28642 6020 30942
rect 6076 30212 6132 30222
rect 6076 30118 6132 30156
rect 6300 30098 6356 30110
rect 6300 30046 6302 30098
rect 6354 30046 6356 30098
rect 6300 29316 6356 30046
rect 6524 30100 6580 32620
rect 6636 31220 6692 34076
rect 6860 34066 6916 34076
rect 6860 33572 6916 33582
rect 6860 33234 6916 33516
rect 6860 33182 6862 33234
rect 6914 33182 6916 33234
rect 6860 33170 6916 33182
rect 6972 32004 7028 38894
rect 7196 37492 7252 40684
rect 7420 40402 7476 41356
rect 7644 41300 7700 41310
rect 7756 41300 7812 45388
rect 8204 45332 8260 45342
rect 8204 45218 8260 45276
rect 8204 45166 8206 45218
rect 8258 45166 8260 45218
rect 8204 45154 8260 45166
rect 8540 45330 8596 45342
rect 8540 45278 8542 45330
rect 8594 45278 8596 45330
rect 7868 45108 7924 45118
rect 7868 45106 8036 45108
rect 7868 45054 7870 45106
rect 7922 45054 8036 45106
rect 7868 45052 8036 45054
rect 7868 45042 7924 45052
rect 7868 44436 7924 44446
rect 7868 42082 7924 44380
rect 7980 43538 8036 45052
rect 8428 45106 8484 45118
rect 8428 45054 8430 45106
rect 8482 45054 8484 45106
rect 8316 44436 8372 44446
rect 8316 44322 8372 44380
rect 8316 44270 8318 44322
rect 8370 44270 8372 44322
rect 8316 44258 8372 44270
rect 8428 43876 8484 45054
rect 8540 44324 8596 45278
rect 8652 44660 8708 45500
rect 8764 45444 8820 45724
rect 8988 45668 9044 46398
rect 9212 45890 9268 47292
rect 9212 45838 9214 45890
rect 9266 45838 9268 45890
rect 9212 45826 9268 45838
rect 8988 45602 9044 45612
rect 8764 45388 9156 45444
rect 8764 45108 8820 45118
rect 8764 45014 8820 45052
rect 8652 44604 8820 44660
rect 8540 44258 8596 44268
rect 8652 44434 8708 44446
rect 8652 44382 8654 44434
rect 8706 44382 8708 44434
rect 7980 43486 7982 43538
rect 8034 43486 8036 43538
rect 7980 42868 8036 43486
rect 7980 42802 8036 42812
rect 8092 43820 8484 43876
rect 8092 43426 8148 43820
rect 8316 43652 8372 43662
rect 8092 43374 8094 43426
rect 8146 43374 8148 43426
rect 8092 42532 8148 43374
rect 8092 42466 8148 42476
rect 8204 43650 8372 43652
rect 8204 43598 8318 43650
rect 8370 43598 8372 43650
rect 8204 43596 8372 43598
rect 8204 42308 8260 43596
rect 8316 43586 8372 43596
rect 8316 42868 8372 42878
rect 8652 42868 8708 44382
rect 8764 44100 8820 44604
rect 8764 44044 9044 44100
rect 8876 43652 8932 43662
rect 8316 42754 8372 42812
rect 8316 42702 8318 42754
rect 8370 42702 8372 42754
rect 8316 42690 8372 42702
rect 8540 42866 8708 42868
rect 8540 42814 8654 42866
rect 8706 42814 8708 42866
rect 8540 42812 8708 42814
rect 7868 42030 7870 42082
rect 7922 42030 7924 42082
rect 7868 41636 7924 42030
rect 7980 42252 8260 42308
rect 7980 42082 8036 42252
rect 7980 42030 7982 42082
rect 8034 42030 8036 42082
rect 7980 42018 8036 42030
rect 8092 42084 8148 42094
rect 7868 41570 7924 41580
rect 7700 41244 7812 41300
rect 7644 41234 7700 41244
rect 7532 41188 7588 41198
rect 7532 41094 7588 41132
rect 7756 41076 7812 41086
rect 8092 41076 8148 42028
rect 7756 41074 7924 41076
rect 7756 41022 7758 41074
rect 7810 41022 7924 41074
rect 7756 41020 7924 41022
rect 7756 41010 7812 41020
rect 7644 40964 7700 40974
rect 7532 40516 7588 40526
rect 7532 40422 7588 40460
rect 7420 40350 7422 40402
rect 7474 40350 7476 40402
rect 7420 40338 7476 40350
rect 7308 39732 7364 39742
rect 7308 39506 7364 39676
rect 7308 39454 7310 39506
rect 7362 39454 7364 39506
rect 7308 38946 7364 39454
rect 7308 38894 7310 38946
rect 7362 38894 7364 38946
rect 7308 38724 7364 38894
rect 7532 38836 7588 38846
rect 7644 38836 7700 40908
rect 7756 40628 7812 40638
rect 7756 40534 7812 40572
rect 7868 39844 7924 41020
rect 8092 40516 8148 41020
rect 8204 40964 8260 42252
rect 8316 42308 8372 42318
rect 8316 41970 8372 42252
rect 8316 41918 8318 41970
rect 8370 41918 8372 41970
rect 8316 41188 8372 41918
rect 8540 41412 8596 42812
rect 8652 42802 8708 42812
rect 8764 43596 8876 43652
rect 8652 42420 8708 42430
rect 8764 42420 8820 43596
rect 8876 43558 8932 43596
rect 8988 43540 9044 44044
rect 9100 43652 9156 45388
rect 9324 44548 9380 47406
rect 9436 45332 9492 50540
rect 9548 50482 9604 50764
rect 9996 50708 10052 51772
rect 10108 51762 10164 51772
rect 9548 50430 9550 50482
rect 9602 50430 9604 50482
rect 9548 50418 9604 50430
rect 9884 50594 9940 50606
rect 9884 50542 9886 50594
rect 9938 50542 9940 50594
rect 9660 49924 9716 49934
rect 9548 48130 9604 48142
rect 9548 48078 9550 48130
rect 9602 48078 9604 48130
rect 9548 47348 9604 48078
rect 9548 47282 9604 47292
rect 9660 47236 9716 49868
rect 9884 49140 9940 50542
rect 9996 50428 10052 50652
rect 10220 51602 10276 51884
rect 10220 51550 10222 51602
rect 10274 51550 10276 51602
rect 10220 50820 10276 51550
rect 10108 50596 10164 50634
rect 10108 50530 10164 50540
rect 9996 50372 10164 50428
rect 9884 49074 9940 49084
rect 10108 49138 10164 50372
rect 10220 50034 10276 50764
rect 10220 49982 10222 50034
rect 10274 49982 10276 50034
rect 10220 49970 10276 49982
rect 10332 51938 10500 51940
rect 10332 51886 10446 51938
rect 10498 51886 10500 51938
rect 10332 51884 10500 51886
rect 10108 49086 10110 49138
rect 10162 49086 10164 49138
rect 10108 49074 10164 49086
rect 9660 47170 9716 47180
rect 9772 48130 9828 48142
rect 9772 48078 9774 48130
rect 9826 48078 9828 48130
rect 9660 47012 9716 47022
rect 9548 46676 9604 46686
rect 9548 46582 9604 46620
rect 9660 46676 9716 46956
rect 9772 46900 9828 48078
rect 9884 47796 9940 47806
rect 9940 47740 10052 47796
rect 9884 47730 9940 47740
rect 9772 46834 9828 46844
rect 9884 47124 9940 47134
rect 9772 46676 9828 46686
rect 9660 46674 9828 46676
rect 9660 46622 9774 46674
rect 9826 46622 9828 46674
rect 9660 46620 9828 46622
rect 9660 45892 9716 46620
rect 9772 46610 9828 46620
rect 9772 46116 9828 46126
rect 9884 46116 9940 47068
rect 9772 46114 9940 46116
rect 9772 46062 9774 46114
rect 9826 46062 9940 46114
rect 9772 46060 9940 46062
rect 9996 46114 10052 47740
rect 10332 47684 10388 51884
rect 10444 51874 10500 51884
rect 10668 50596 10724 50606
rect 10444 50372 10500 50382
rect 10444 50278 10500 50316
rect 10444 49140 10500 49150
rect 10444 49046 10500 49084
rect 10668 49026 10724 50540
rect 10668 48974 10670 49026
rect 10722 48974 10724 49026
rect 10668 48692 10724 48974
rect 10108 47628 10388 47684
rect 10444 48636 10724 48692
rect 10108 47012 10164 47628
rect 10332 47460 10388 47470
rect 10444 47460 10500 48636
rect 10668 48356 10724 48366
rect 10668 48354 10836 48356
rect 10668 48302 10670 48354
rect 10722 48302 10836 48354
rect 10668 48300 10836 48302
rect 10668 48290 10724 48300
rect 10556 48244 10612 48254
rect 10556 47796 10612 48188
rect 10556 47740 10724 47796
rect 10332 47458 10500 47460
rect 10332 47406 10334 47458
rect 10386 47406 10500 47458
rect 10332 47404 10500 47406
rect 10556 47572 10612 47582
rect 10556 47458 10612 47516
rect 10556 47406 10558 47458
rect 10610 47406 10612 47458
rect 10332 47394 10388 47404
rect 10556 47394 10612 47406
rect 10108 46946 10164 46956
rect 10332 47236 10388 47246
rect 10220 46900 10276 46910
rect 9996 46062 9998 46114
rect 10050 46062 10052 46114
rect 9772 46050 9828 46060
rect 9996 46050 10052 46062
rect 10108 46450 10164 46462
rect 10108 46398 10110 46450
rect 10162 46398 10164 46450
rect 10108 45892 10164 46398
rect 9660 45836 9828 45892
rect 9660 45668 9716 45678
rect 9660 45574 9716 45612
rect 9772 45556 9828 45836
rect 10108 45826 10164 45836
rect 9772 45490 9828 45500
rect 9436 45276 9940 45332
rect 9548 45108 9604 45118
rect 9548 45014 9604 45052
rect 9324 44482 9380 44492
rect 9100 43586 9156 43596
rect 9660 43652 9716 43662
rect 9660 43558 9716 43596
rect 9884 43652 9940 45276
rect 8988 43446 9044 43484
rect 9548 43540 9604 43550
rect 9548 43446 9604 43484
rect 8876 43316 8932 43326
rect 8876 43222 8932 43260
rect 8708 42364 8820 42420
rect 9884 42644 9940 43596
rect 9996 44994 10052 45006
rect 9996 44942 9998 44994
rect 10050 44942 10052 44994
rect 9996 43540 10052 44942
rect 10220 44436 10276 46844
rect 10332 45444 10388 47180
rect 10668 47236 10724 47740
rect 10444 46788 10500 46798
rect 10668 46788 10724 47180
rect 10444 46694 10500 46732
rect 10556 46786 10724 46788
rect 10556 46734 10670 46786
rect 10722 46734 10724 46786
rect 10556 46732 10724 46734
rect 10556 46564 10612 46732
rect 10668 46722 10724 46732
rect 10780 46786 10836 48300
rect 10892 47572 10948 52780
rect 11228 52834 11284 53452
rect 11228 52782 11230 52834
rect 11282 52782 11284 52834
rect 11228 50932 11284 52782
rect 11564 52834 11620 53676
rect 11564 52782 11566 52834
rect 11618 52782 11620 52834
rect 11564 52770 11620 52782
rect 11340 52724 11396 52734
rect 11676 52724 11732 53790
rect 11900 53620 11956 55022
rect 12348 55076 12404 55086
rect 12348 54982 12404 55020
rect 12684 54740 12740 55132
rect 12572 54738 12740 54740
rect 12572 54686 12686 54738
rect 12738 54686 12740 54738
rect 12572 54684 12740 54686
rect 12460 54514 12516 54526
rect 12460 54462 12462 54514
rect 12514 54462 12516 54514
rect 12124 54404 12180 54414
rect 12124 54310 12180 54348
rect 12236 54292 12292 54302
rect 12236 54198 12292 54236
rect 12460 53956 12516 54462
rect 12460 53890 12516 53900
rect 11900 53554 11956 53564
rect 12348 53620 12404 53630
rect 12348 53526 12404 53564
rect 12572 53618 12628 54684
rect 12684 54674 12740 54684
rect 12572 53566 12574 53618
rect 12626 53566 12628 53618
rect 12572 53554 12628 53566
rect 12796 54516 12852 54526
rect 11340 52722 11508 52724
rect 11340 52670 11342 52722
rect 11394 52670 11508 52722
rect 11340 52668 11508 52670
rect 11340 52658 11396 52668
rect 11228 50866 11284 50876
rect 11228 50482 11284 50494
rect 11228 50430 11230 50482
rect 11282 50430 11284 50482
rect 11228 50428 11284 50430
rect 11228 50372 11396 50428
rect 11004 49252 11060 49262
rect 11004 49158 11060 49196
rect 11340 49138 11396 50372
rect 11340 49086 11342 49138
rect 11394 49086 11396 49138
rect 11340 49074 11396 49086
rect 11340 48916 11396 48926
rect 10892 47506 10948 47516
rect 11228 47684 11284 47694
rect 11228 47458 11284 47628
rect 11228 47406 11230 47458
rect 11282 47406 11284 47458
rect 11228 47394 11284 47406
rect 10780 46734 10782 46786
rect 10834 46734 10836 46786
rect 10780 46722 10836 46734
rect 10892 47234 10948 47246
rect 10892 47182 10894 47234
rect 10946 47182 10948 47234
rect 10892 46788 10948 47182
rect 11116 47234 11172 47246
rect 11116 47182 11118 47234
rect 11170 47182 11172 47234
rect 11116 46900 11172 47182
rect 11116 46834 11172 46844
rect 10892 46722 10948 46732
rect 10444 46508 10612 46564
rect 10444 45890 10500 46508
rect 11004 46452 11060 46462
rect 11228 46452 11284 46462
rect 10444 45838 10446 45890
rect 10498 45838 10500 45890
rect 10444 45826 10500 45838
rect 10668 46450 11060 46452
rect 10668 46398 11006 46450
rect 11058 46398 11060 46450
rect 10668 46396 11060 46398
rect 10556 45778 10612 45790
rect 10556 45726 10558 45778
rect 10610 45726 10612 45778
rect 10556 45444 10612 45726
rect 10332 45388 10612 45444
rect 10220 44370 10276 44380
rect 10332 44548 10388 44558
rect 10332 44434 10388 44492
rect 10332 44382 10334 44434
rect 10386 44382 10388 44434
rect 10332 44370 10388 44382
rect 10220 44100 10276 44110
rect 10220 43762 10276 44044
rect 10220 43710 10222 43762
rect 10274 43710 10276 43762
rect 9996 43474 10052 43484
rect 10108 43650 10164 43662
rect 10108 43598 10110 43650
rect 10162 43598 10164 43650
rect 10108 43428 10164 43598
rect 10108 43362 10164 43372
rect 8652 42354 8708 42364
rect 8652 41972 8708 41982
rect 8652 41878 8708 41916
rect 8876 41860 8932 41870
rect 9772 41860 9828 41870
rect 8932 41804 9044 41860
rect 8876 41794 8932 41804
rect 8764 41746 8820 41758
rect 8764 41694 8766 41746
rect 8818 41694 8820 41746
rect 8764 41636 8820 41694
rect 8764 41570 8820 41580
rect 8652 41412 8708 41422
rect 8540 41410 8708 41412
rect 8540 41358 8654 41410
rect 8706 41358 8708 41410
rect 8540 41356 8708 41358
rect 8652 41346 8708 41356
rect 8316 41094 8372 41132
rect 8988 41188 9044 41804
rect 9772 41766 9828 41804
rect 9660 41746 9716 41758
rect 9660 41694 9662 41746
rect 9714 41694 9716 41746
rect 9324 41188 9380 41198
rect 8988 41186 9380 41188
rect 8988 41134 9326 41186
rect 9378 41134 9380 41186
rect 8988 41132 9380 41134
rect 8204 40908 8372 40964
rect 8092 40450 8148 40460
rect 7868 39778 7924 39788
rect 8316 39842 8372 40908
rect 8316 39790 8318 39842
rect 8370 39790 8372 39842
rect 8316 39778 8372 39790
rect 8540 40402 8596 40414
rect 8540 40350 8542 40402
rect 8594 40350 8596 40402
rect 7532 38834 7700 38836
rect 7532 38782 7534 38834
rect 7586 38782 7700 38834
rect 7532 38780 7700 38782
rect 7756 39730 7812 39742
rect 7756 39678 7758 39730
rect 7810 39678 7812 39730
rect 7532 38770 7588 38780
rect 7308 38658 7364 38668
rect 7756 38052 7812 39678
rect 8540 39732 8596 40350
rect 8988 40402 9044 41132
rect 9324 41122 9380 41132
rect 9548 41076 9604 41086
rect 9548 40982 9604 41020
rect 8988 40350 8990 40402
rect 9042 40350 9044 40402
rect 8988 40338 9044 40350
rect 8540 39666 8596 39676
rect 8876 40292 8932 40302
rect 7868 39620 7924 39630
rect 7868 39526 7924 39564
rect 8876 39618 8932 40236
rect 8876 39566 8878 39618
rect 8930 39566 8932 39618
rect 8876 39554 8932 39566
rect 9660 39618 9716 41694
rect 9884 41412 9940 42588
rect 10108 41748 10164 41758
rect 10220 41748 10276 43710
rect 10332 42644 10388 42654
rect 10332 42550 10388 42588
rect 10164 41692 10276 41748
rect 10108 41682 10164 41692
rect 9884 41186 9940 41356
rect 9884 41134 9886 41186
rect 9938 41134 9940 41186
rect 9884 41122 9940 41134
rect 9772 40964 9828 40974
rect 9772 40870 9828 40908
rect 10332 40628 10388 40638
rect 9884 40404 9940 40414
rect 9884 40290 9940 40348
rect 9884 40238 9886 40290
rect 9938 40238 9940 40290
rect 9884 40226 9940 40238
rect 9772 39844 9828 39854
rect 9828 39788 9940 39844
rect 9772 39778 9828 39788
rect 9660 39566 9662 39618
rect 9714 39566 9716 39618
rect 8540 39508 8596 39518
rect 8540 38836 8596 39452
rect 8652 39508 8708 39518
rect 8652 39506 8820 39508
rect 8652 39454 8654 39506
rect 8706 39454 8820 39506
rect 8652 39452 8820 39454
rect 8652 39442 8708 39452
rect 8428 38834 8596 38836
rect 8428 38782 8542 38834
rect 8594 38782 8596 38834
rect 8428 38780 8596 38782
rect 8316 38722 8372 38734
rect 8316 38670 8318 38722
rect 8370 38670 8372 38722
rect 8316 38668 8372 38670
rect 7868 38612 7924 38622
rect 8092 38612 8372 38668
rect 7868 38610 8036 38612
rect 7868 38558 7870 38610
rect 7922 38558 8036 38610
rect 7868 38556 8036 38558
rect 7868 38546 7924 38556
rect 7756 37996 7924 38052
rect 7756 37826 7812 37838
rect 7756 37774 7758 37826
rect 7810 37774 7812 37826
rect 7196 37436 7364 37492
rect 7196 37266 7252 37278
rect 7196 37214 7198 37266
rect 7250 37214 7252 37266
rect 7196 36708 7252 37214
rect 7084 36652 7196 36708
rect 7084 35812 7140 36652
rect 7196 36642 7252 36652
rect 7308 36484 7364 37436
rect 7084 35698 7140 35756
rect 7084 35646 7086 35698
rect 7138 35646 7140 35698
rect 7084 35634 7140 35646
rect 7196 36428 7364 36484
rect 7420 37380 7476 37390
rect 7756 37380 7812 37774
rect 7868 37716 7924 37996
rect 7868 37650 7924 37660
rect 7420 37378 7812 37380
rect 7420 37326 7422 37378
rect 7474 37326 7812 37378
rect 7420 37324 7812 37326
rect 7980 37380 8036 38556
rect 7196 35924 7252 36428
rect 7084 33908 7140 33918
rect 7084 33814 7140 33852
rect 7196 33572 7252 35868
rect 7308 35810 7364 35822
rect 7308 35758 7310 35810
rect 7362 35758 7364 35810
rect 7308 34916 7364 35758
rect 7420 35700 7476 37324
rect 7980 37314 8036 37324
rect 8092 38050 8148 38612
rect 8428 38500 8484 38780
rect 8540 38770 8596 38780
rect 8652 39172 8708 39182
rect 8652 38668 8708 39116
rect 8764 39060 8820 39452
rect 8876 39060 8932 39070
rect 8764 39058 9604 39060
rect 8764 39006 8878 39058
rect 8930 39006 9604 39058
rect 8764 39004 9604 39006
rect 8876 38994 8932 39004
rect 9548 38834 9604 39004
rect 9548 38782 9550 38834
rect 9602 38782 9604 38834
rect 9548 38770 9604 38782
rect 9660 38668 9716 39566
rect 8652 38612 8820 38668
rect 8316 38444 8484 38500
rect 8316 38052 8372 38444
rect 8092 37998 8094 38050
rect 8146 37998 8148 38050
rect 7980 37042 8036 37054
rect 7980 36990 7982 37042
rect 8034 36990 8036 37042
rect 7868 36260 7924 36270
rect 7420 35634 7476 35644
rect 7644 36258 7924 36260
rect 7644 36206 7870 36258
rect 7922 36206 7924 36258
rect 7644 36204 7924 36206
rect 7644 35364 7700 36204
rect 7868 36194 7924 36204
rect 7756 35812 7812 35822
rect 7756 35698 7812 35756
rect 7980 35812 8036 36990
rect 7980 35718 8036 35756
rect 7756 35646 7758 35698
rect 7810 35646 7812 35698
rect 7756 35634 7812 35646
rect 8092 35476 8148 37998
rect 8204 38050 8372 38052
rect 8204 37998 8318 38050
rect 8370 37998 8372 38050
rect 8204 37996 8372 37998
rect 8204 37268 8260 37996
rect 8316 37986 8372 37996
rect 8652 38052 8708 38062
rect 8652 37958 8708 37996
rect 8316 37716 8372 37726
rect 8316 37490 8372 37660
rect 8316 37438 8318 37490
rect 8370 37438 8372 37490
rect 8316 37426 8372 37438
rect 8652 37492 8708 37502
rect 8652 37398 8708 37436
rect 8204 37212 8372 37268
rect 7644 35298 7700 35308
rect 7756 35420 8148 35476
rect 7308 34850 7364 34860
rect 7420 35252 7476 35262
rect 7196 33516 7364 33572
rect 7084 33460 7140 33470
rect 7084 33366 7140 33404
rect 7196 33348 7252 33358
rect 7196 33254 7252 33292
rect 7308 33124 7364 33516
rect 6636 31154 6692 31164
rect 6748 31948 7028 32004
rect 7196 33068 7364 33124
rect 6636 30100 6692 30110
rect 6524 30098 6692 30100
rect 6524 30046 6638 30098
rect 6690 30046 6692 30098
rect 6524 30044 6692 30046
rect 6636 30034 6692 30044
rect 6300 29250 6356 29260
rect 5964 28590 5966 28642
rect 6018 28590 6020 28642
rect 5964 28578 6020 28590
rect 6188 29204 6244 29214
rect 6188 28642 6244 29148
rect 6188 28590 6190 28642
rect 6242 28590 6244 28642
rect 6188 28578 6244 28590
rect 5740 28530 5908 28532
rect 5740 28478 5742 28530
rect 5794 28478 5908 28530
rect 5740 28476 5908 28478
rect 5740 28466 5796 28476
rect 5404 28252 6132 28308
rect 4508 28196 4564 28206
rect 4564 28140 4676 28196
rect 4508 28130 4564 28140
rect 4172 28082 4340 28084
rect 4172 28030 4286 28082
rect 4338 28030 4340 28082
rect 4172 28028 4340 28030
rect 3500 27918 3502 27970
rect 3554 27918 3556 27970
rect 2940 26572 3108 26628
rect 2940 26402 2996 26414
rect 2940 26350 2942 26402
rect 2994 26350 2996 26402
rect 2940 25732 2996 26350
rect 2940 25666 2996 25676
rect 2940 24500 2996 24510
rect 2828 24444 2940 24500
rect 2940 24434 2996 24444
rect 2716 24220 2996 24276
rect 2604 24108 2884 24164
rect 2380 21810 2548 21812
rect 2380 21758 2382 21810
rect 2434 21758 2548 21810
rect 2380 21756 2548 21758
rect 2604 23940 2660 23950
rect 2604 23266 2660 23884
rect 2604 23214 2606 23266
rect 2658 23214 2660 23266
rect 2604 22596 2660 23214
rect 2828 23156 2884 24108
rect 2380 21746 2436 21756
rect 2492 21588 2548 21598
rect 1932 19180 2100 19236
rect 2156 20132 2324 20188
rect 2380 21532 2492 21588
rect 1484 18386 1540 18396
rect 1596 18676 1652 18686
rect 1372 16706 1428 16716
rect 1260 15474 1316 15484
rect 1596 13186 1652 18620
rect 1932 14980 1988 19180
rect 2044 19010 2100 19022
rect 2044 18958 2046 19010
rect 2098 18958 2100 19010
rect 2044 18564 2100 18958
rect 2044 18498 2100 18508
rect 2044 17780 2100 17790
rect 2044 17686 2100 17724
rect 2156 16996 2212 20132
rect 2268 18338 2324 18350
rect 2268 18286 2270 18338
rect 2322 18286 2324 18338
rect 2268 18228 2324 18286
rect 2268 18162 2324 18172
rect 2044 16940 2212 16996
rect 2044 15540 2100 16940
rect 2156 16770 2212 16782
rect 2156 16718 2158 16770
rect 2210 16718 2212 16770
rect 2156 16658 2212 16718
rect 2156 16606 2158 16658
rect 2210 16606 2212 16658
rect 2156 16594 2212 16606
rect 2268 16772 2324 16782
rect 2268 16210 2324 16716
rect 2268 16158 2270 16210
rect 2322 16158 2324 16210
rect 2268 15988 2324 16158
rect 2268 15922 2324 15932
rect 2380 15540 2436 21532
rect 2492 21522 2548 21532
rect 2604 20804 2660 22540
rect 2604 20738 2660 20748
rect 2716 23154 2884 23156
rect 2716 23102 2830 23154
rect 2882 23102 2884 23154
rect 2716 23100 2884 23102
rect 2716 21028 2772 23100
rect 2828 23090 2884 23100
rect 2716 20802 2772 20972
rect 2716 20750 2718 20802
rect 2770 20750 2772 20802
rect 2716 20738 2772 20750
rect 2604 20580 2660 20590
rect 2604 20486 2660 20524
rect 2492 20356 2548 20366
rect 2492 20130 2548 20300
rect 2940 20188 2996 24220
rect 3052 21588 3108 26572
rect 3500 26404 3556 27918
rect 4060 27972 4116 27982
rect 3724 27860 3780 27870
rect 3724 27766 3780 27804
rect 3948 27860 4004 27870
rect 3500 25508 3556 26348
rect 3500 25442 3556 25452
rect 3724 27074 3780 27086
rect 3724 27022 3726 27074
rect 3778 27022 3780 27074
rect 3724 25284 3780 27022
rect 3948 26908 4004 27804
rect 4060 27076 4116 27916
rect 4172 27188 4228 28028
rect 4284 28018 4340 28028
rect 4508 27972 4564 27982
rect 4508 27878 4564 27916
rect 4620 27970 4676 28140
rect 5516 28084 5572 28094
rect 4620 27918 4622 27970
rect 4674 27918 4676 27970
rect 4620 27906 4676 27918
rect 5404 27970 5460 27982
rect 5404 27918 5406 27970
rect 5458 27918 5460 27970
rect 4956 27858 5012 27870
rect 4956 27806 4958 27858
rect 5010 27806 5012 27858
rect 4620 27748 4676 27758
rect 4620 27746 4900 27748
rect 4620 27694 4622 27746
rect 4674 27694 4900 27746
rect 4620 27692 4900 27694
rect 4620 27682 4676 27692
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4396 27188 4452 27198
rect 4172 27186 4452 27188
rect 4172 27134 4398 27186
rect 4450 27134 4452 27186
rect 4172 27132 4452 27134
rect 4396 27122 4452 27132
rect 4060 27010 4116 27020
rect 4620 27076 4676 27086
rect 4620 26982 4676 27020
rect 3836 26852 4004 26908
rect 4732 26964 4788 26974
rect 4732 26870 4788 26908
rect 3836 25508 3892 26852
rect 4844 26292 4900 27692
rect 4956 26908 5012 27806
rect 5404 26908 5460 27918
rect 5516 27076 5572 28028
rect 5628 27860 5684 27870
rect 5628 27766 5684 27804
rect 5628 27076 5684 27086
rect 5516 27074 5684 27076
rect 5516 27022 5630 27074
rect 5682 27022 5684 27074
rect 5516 27020 5684 27022
rect 5628 27010 5684 27020
rect 4956 26852 5348 26908
rect 5404 26852 5572 26908
rect 4844 26226 4900 26236
rect 5180 26402 5236 26414
rect 5180 26350 5182 26402
rect 5234 26350 5236 26402
rect 4284 26180 4340 26190
rect 3836 25452 4228 25508
rect 4060 25284 4116 25294
rect 3724 25282 3892 25284
rect 3724 25230 3726 25282
rect 3778 25230 3892 25282
rect 3724 25228 3892 25230
rect 3724 25218 3780 25228
rect 3836 25060 3892 25228
rect 3836 24994 3892 25004
rect 3948 25282 4116 25284
rect 3948 25230 4062 25282
rect 4114 25230 4116 25282
rect 3948 25228 4116 25230
rect 3500 24724 3556 24734
rect 3836 24724 3892 24734
rect 3500 24162 3556 24668
rect 3500 24110 3502 24162
rect 3554 24110 3556 24162
rect 3500 24098 3556 24110
rect 3724 24722 3892 24724
rect 3724 24670 3838 24722
rect 3890 24670 3892 24722
rect 3724 24668 3892 24670
rect 3724 23828 3780 24668
rect 3836 24658 3892 24668
rect 3612 23772 3780 23828
rect 3836 24276 3892 24286
rect 3612 23548 3668 23772
rect 3388 23492 3668 23548
rect 3724 23604 3780 23614
rect 3164 23156 3220 23166
rect 3164 23042 3220 23100
rect 3164 22990 3166 23042
rect 3218 22990 3220 23042
rect 3164 22978 3220 22990
rect 3052 21522 3108 21532
rect 3164 22820 3220 22830
rect 3052 20804 3108 20814
rect 3052 20710 3108 20748
rect 2492 20078 2494 20130
rect 2546 20078 2548 20130
rect 2492 20066 2548 20078
rect 2828 20132 2996 20188
rect 2828 18900 2884 20132
rect 2940 19796 2996 19806
rect 2940 19122 2996 19740
rect 2940 19070 2942 19122
rect 2994 19070 2996 19122
rect 2940 19058 2996 19070
rect 2828 18844 2996 18900
rect 2716 18452 2772 18462
rect 2716 18358 2772 18396
rect 2492 17444 2548 17454
rect 2828 17444 2884 17454
rect 2492 17442 2884 17444
rect 2492 17390 2494 17442
rect 2546 17390 2830 17442
rect 2882 17390 2884 17442
rect 2492 17388 2884 17390
rect 2940 17444 2996 18844
rect 3052 18450 3108 18462
rect 3052 18398 3054 18450
rect 3106 18398 3108 18450
rect 3052 17892 3108 18398
rect 3052 17826 3108 17836
rect 2940 17388 3108 17444
rect 2492 17378 2548 17388
rect 2828 17332 2884 17388
rect 2884 17276 2996 17332
rect 2828 17266 2884 17276
rect 2604 17108 2660 17118
rect 2604 17014 2660 17052
rect 2940 17106 2996 17276
rect 2940 17054 2942 17106
rect 2994 17054 2996 17106
rect 2940 17042 2996 17054
rect 3052 16884 3108 17388
rect 2940 16828 3108 16884
rect 2716 15874 2772 15886
rect 2716 15822 2718 15874
rect 2770 15822 2772 15874
rect 2716 15652 2772 15822
rect 2716 15586 2772 15596
rect 2492 15540 2548 15550
rect 2044 15538 2212 15540
rect 2044 15486 2046 15538
rect 2098 15486 2212 15538
rect 2044 15484 2212 15486
rect 2380 15538 2548 15540
rect 2380 15486 2494 15538
rect 2546 15486 2548 15538
rect 2380 15484 2548 15486
rect 2044 15474 2100 15484
rect 2156 15092 2212 15484
rect 2492 15474 2548 15484
rect 2716 15428 2772 15438
rect 2156 15036 2436 15092
rect 1932 14924 2212 14980
rect 1596 13134 1598 13186
rect 1650 13134 1652 13186
rect 1596 13122 1652 13134
rect 1932 14306 1988 14318
rect 1932 14254 1934 14306
rect 1986 14254 1988 14306
rect 1932 13188 1988 14254
rect 2156 13970 2212 14924
rect 2156 13918 2158 13970
rect 2210 13918 2212 13970
rect 2156 13906 2212 13918
rect 2380 13860 2436 15036
rect 2492 14644 2548 14654
rect 2492 14550 2548 14588
rect 2716 13970 2772 15372
rect 2716 13918 2718 13970
rect 2770 13918 2772 13970
rect 2716 13906 2772 13918
rect 2828 15204 2884 15214
rect 2940 15204 2996 16828
rect 3164 16436 3220 22764
rect 3388 21924 3444 23492
rect 3500 23156 3556 23166
rect 3500 23062 3556 23100
rect 3500 22932 3556 22942
rect 3500 22258 3556 22876
rect 3500 22206 3502 22258
rect 3554 22206 3556 22258
rect 3500 22194 3556 22206
rect 3276 21028 3332 21038
rect 3276 20934 3332 20972
rect 2828 15202 2996 15204
rect 2828 15150 2830 15202
rect 2882 15150 2996 15202
rect 2828 15148 2996 15150
rect 3052 16380 3220 16436
rect 3276 19460 3332 19470
rect 3276 16658 3332 19404
rect 3276 16606 3278 16658
rect 3330 16606 3332 16658
rect 2380 13794 2436 13804
rect 1932 13122 1988 13132
rect 2828 13188 2884 15148
rect 2940 14308 2996 14318
rect 2940 14214 2996 14252
rect 3052 13970 3108 16380
rect 3164 16212 3220 16222
rect 3276 16212 3332 16606
rect 3164 16210 3332 16212
rect 3164 16158 3166 16210
rect 3218 16158 3332 16210
rect 3164 16156 3332 16158
rect 3164 16146 3220 16156
rect 3164 15988 3220 15998
rect 3164 14532 3220 15932
rect 3388 15428 3444 21868
rect 3500 21700 3556 21710
rect 3500 21606 3556 21644
rect 3612 20578 3668 20590
rect 3612 20526 3614 20578
rect 3666 20526 3668 20578
rect 3612 18788 3668 20526
rect 3612 18722 3668 18732
rect 3612 18452 3668 18462
rect 3612 18358 3668 18396
rect 3724 17780 3780 23548
rect 3836 23042 3892 24220
rect 3836 22990 3838 23042
rect 3890 22990 3892 23042
rect 3836 22978 3892 22990
rect 3948 21812 4004 25228
rect 4060 25218 4116 25228
rect 4060 24836 4116 24846
rect 4172 24836 4228 25452
rect 4284 25396 4340 26124
rect 4732 26068 4788 26078
rect 4732 26066 4900 26068
rect 4732 26014 4734 26066
rect 4786 26014 4900 26066
rect 4732 26012 4900 26014
rect 4732 26002 4788 26012
rect 4844 25956 4900 26012
rect 5180 25956 5236 26350
rect 4476 25900 4740 25910
rect 4844 25900 5236 25956
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25302 4340 25340
rect 4396 25620 4452 25630
rect 4396 25394 4452 25564
rect 4956 25620 5012 25630
rect 4956 25506 5012 25564
rect 4956 25454 4958 25506
rect 5010 25454 5012 25506
rect 4956 25442 5012 25454
rect 4396 25342 4398 25394
rect 4450 25342 4452 25394
rect 4116 24780 4228 24836
rect 4060 24770 4116 24780
rect 4396 24500 4452 25342
rect 4732 25282 4788 25294
rect 4732 25230 4734 25282
rect 4786 25230 4788 25282
rect 4732 24836 4788 25230
rect 4732 24770 4788 24780
rect 5068 24722 5124 25900
rect 5068 24670 5070 24722
rect 5122 24670 5124 24722
rect 5068 24658 5124 24670
rect 5292 25284 5348 26852
rect 5516 26180 5572 26852
rect 5628 26404 5684 26414
rect 5628 26310 5684 26348
rect 5964 26292 6020 26302
rect 5516 26114 5572 26124
rect 5852 26180 5908 26190
rect 5852 26086 5908 26124
rect 5740 25732 5796 25742
rect 5740 25506 5796 25676
rect 5740 25454 5742 25506
rect 5794 25454 5796 25506
rect 5740 25442 5796 25454
rect 5964 25394 6020 26236
rect 5964 25342 5966 25394
rect 6018 25342 6020 25394
rect 5964 25330 6020 25342
rect 4284 24444 4452 24500
rect 4732 24500 4788 24510
rect 4732 24498 4900 24500
rect 4732 24446 4734 24498
rect 4786 24446 4900 24498
rect 4732 24444 4900 24446
rect 4284 24164 4340 24444
rect 4732 24434 4788 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 24108 4452 24164
rect 4060 23940 4116 23950
rect 4284 23940 4340 23950
rect 4060 23846 4116 23884
rect 4172 23938 4340 23940
rect 4172 23886 4286 23938
rect 4338 23886 4340 23938
rect 4172 23884 4340 23886
rect 3948 21746 4004 21756
rect 4060 23268 4116 23278
rect 3948 20804 4004 20814
rect 4060 20804 4116 23212
rect 4172 21700 4228 23884
rect 4284 23874 4340 23884
rect 4396 23380 4452 24108
rect 4284 23324 4452 23380
rect 4620 23714 4676 23726
rect 4620 23662 4622 23714
rect 4674 23662 4676 23714
rect 4284 21812 4340 23324
rect 4620 23044 4676 23662
rect 4620 22978 4676 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 21746 4340 21756
rect 4620 22482 4676 22494
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 4620 22372 4676 22430
rect 4620 21810 4676 22316
rect 4620 21758 4622 21810
rect 4674 21758 4676 21810
rect 4620 21746 4676 21758
rect 4844 21812 4900 24444
rect 5068 24052 5124 24062
rect 5068 23958 5124 23996
rect 5068 22148 5124 22158
rect 5068 22054 5124 22092
rect 5180 21812 5236 21822
rect 4844 21810 5180 21812
rect 4844 21758 4846 21810
rect 4898 21758 5180 21810
rect 4844 21756 5180 21758
rect 4844 21746 4900 21756
rect 4172 21028 4228 21644
rect 4396 21698 4452 21710
rect 4396 21646 4398 21698
rect 4450 21646 4452 21698
rect 4396 21588 4452 21646
rect 5180 21698 5236 21756
rect 5180 21646 5182 21698
rect 5234 21646 5236 21698
rect 5180 21634 5236 21646
rect 4284 21532 4396 21588
rect 4284 21028 4340 21532
rect 4396 21522 4452 21532
rect 4732 21476 4788 21486
rect 4732 21382 4788 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4508 21028 4564 21038
rect 4284 21026 4564 21028
rect 4284 20974 4510 21026
rect 4562 20974 4564 21026
rect 4284 20972 4564 20974
rect 4172 20934 4228 20972
rect 4508 20962 4564 20972
rect 4844 20804 4900 20814
rect 4060 20748 4228 20804
rect 3948 20710 4004 20748
rect 3948 20580 4004 20590
rect 4004 20524 4116 20580
rect 3948 20514 4004 20524
rect 3724 17714 3780 17724
rect 3836 19796 3892 19806
rect 3836 17554 3892 19740
rect 3948 18564 4004 18574
rect 3948 18338 4004 18508
rect 3948 18286 3950 18338
rect 4002 18286 4004 18338
rect 3948 18228 4004 18286
rect 3948 18162 4004 18172
rect 3836 17502 3838 17554
rect 3890 17502 3892 17554
rect 3836 17490 3892 17502
rect 3948 17108 4004 17118
rect 3948 17014 4004 17052
rect 3388 15362 3444 15372
rect 3500 16770 3556 16782
rect 3500 16718 3502 16770
rect 3554 16718 3556 16770
rect 3388 15204 3444 15242
rect 3388 15138 3444 15148
rect 3276 14532 3332 14542
rect 3164 14530 3332 14532
rect 3164 14478 3278 14530
rect 3330 14478 3332 14530
rect 3164 14476 3332 14478
rect 3276 14466 3332 14476
rect 3500 14532 3556 16718
rect 3612 16212 3668 16222
rect 3612 16118 3668 16156
rect 4060 16212 4116 20524
rect 4172 17892 4228 20748
rect 4844 20802 5124 20804
rect 4844 20750 4846 20802
rect 4898 20750 5124 20802
rect 4844 20748 5124 20750
rect 4844 20738 4900 20748
rect 4956 20578 5012 20590
rect 4956 20526 4958 20578
rect 5010 20526 5012 20578
rect 4620 19906 4676 19918
rect 4620 19854 4622 19906
rect 4674 19854 4676 19906
rect 4620 19796 4676 19854
rect 4956 19796 5012 20526
rect 5068 19908 5124 20748
rect 5180 20580 5236 20590
rect 5180 20486 5236 20524
rect 5292 20356 5348 25228
rect 5628 25282 5684 25294
rect 5628 25230 5630 25282
rect 5682 25230 5684 25282
rect 5628 25060 5684 25230
rect 5852 25284 5908 25322
rect 5852 25218 5908 25228
rect 5964 25172 6020 25182
rect 5852 25060 5908 25070
rect 5628 25004 5796 25060
rect 5628 24836 5684 24846
rect 5628 24742 5684 24780
rect 5740 23380 5796 25004
rect 5852 24724 5908 25004
rect 5852 24630 5908 24668
rect 5852 24052 5908 24062
rect 5964 24052 6020 25116
rect 5852 24050 6020 24052
rect 5852 23998 5854 24050
rect 5906 23998 6020 24050
rect 5852 23996 6020 23998
rect 5852 23604 5908 23996
rect 5852 23538 5908 23548
rect 5740 23324 5908 23380
rect 5628 23044 5684 23054
rect 5628 22370 5684 22988
rect 5628 22318 5630 22370
rect 5682 22318 5684 22370
rect 5628 22306 5684 22318
rect 5404 22148 5460 22158
rect 5404 21588 5460 22092
rect 5404 21586 5684 21588
rect 5404 21534 5406 21586
rect 5458 21534 5684 21586
rect 5404 21532 5684 21534
rect 5404 21522 5460 21532
rect 5628 21026 5684 21532
rect 5628 20974 5630 21026
rect 5682 20974 5684 21026
rect 5628 20962 5684 20974
rect 5740 21028 5796 21038
rect 5516 20916 5572 20926
rect 5292 20300 5460 20356
rect 5180 20132 5236 20142
rect 5180 20038 5236 20076
rect 5292 20130 5348 20142
rect 5292 20078 5294 20130
rect 5346 20078 5348 20130
rect 5292 20020 5348 20078
rect 5292 19954 5348 19964
rect 5068 19852 5236 19908
rect 4676 19740 4900 19796
rect 4620 19730 4676 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4732 19234 4788 19246
rect 4732 19182 4734 19234
rect 4786 19182 4788 19234
rect 4732 19124 4788 19182
rect 4732 19058 4788 19068
rect 4844 18562 4900 19740
rect 4956 19730 5012 19740
rect 4844 18510 4846 18562
rect 4898 18510 4900 18562
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4172 17836 4564 17892
rect 4396 17668 4452 17678
rect 4396 17108 4452 17612
rect 4396 17014 4452 17052
rect 4508 16996 4564 17836
rect 4844 17220 4900 18510
rect 4956 19572 5012 19582
rect 4956 17668 5012 19516
rect 4956 17602 5012 17612
rect 4956 17444 5012 17454
rect 4956 17350 5012 17388
rect 4844 17164 5124 17220
rect 4844 16996 4900 17006
rect 4508 16994 4900 16996
rect 4508 16942 4846 16994
rect 4898 16942 4900 16994
rect 4508 16940 4900 16942
rect 4844 16930 4900 16940
rect 5068 16994 5124 17164
rect 5068 16942 5070 16994
rect 5122 16942 5124 16994
rect 5068 16930 5124 16942
rect 4284 16884 4340 16894
rect 3948 16100 4004 16110
rect 4060 16100 4116 16156
rect 3948 16098 4116 16100
rect 3948 16046 3950 16098
rect 4002 16046 4116 16098
rect 3948 16044 4116 16046
rect 4172 16324 4228 16334
rect 3948 16034 4004 16044
rect 4172 15986 4228 16268
rect 4172 15934 4174 15986
rect 4226 15934 4228 15986
rect 4172 15922 4228 15934
rect 3948 15764 4004 15774
rect 4284 15764 4340 16828
rect 5180 16882 5236 19852
rect 5180 16830 5182 16882
rect 5234 16830 5236 16882
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 5180 16436 5236 16830
rect 5180 16370 5236 16380
rect 4732 16324 4788 16334
rect 4620 16098 4676 16110
rect 4620 16046 4622 16098
rect 4674 16046 4676 16098
rect 4620 15988 4676 16046
rect 4732 16098 4788 16268
rect 5404 16324 5460 20300
rect 5516 20130 5572 20860
rect 5740 20914 5796 20972
rect 5740 20862 5742 20914
rect 5794 20862 5796 20914
rect 5740 20850 5796 20862
rect 5516 20078 5518 20130
rect 5570 20078 5572 20130
rect 5516 20066 5572 20078
rect 5740 20018 5796 20030
rect 5740 19966 5742 20018
rect 5794 19966 5796 20018
rect 5740 19348 5796 19966
rect 5516 19292 5796 19348
rect 5516 18340 5572 19292
rect 5628 19124 5684 19134
rect 5628 19030 5684 19068
rect 5516 18274 5572 18284
rect 5628 17780 5684 17790
rect 5628 17106 5684 17724
rect 5852 17668 5908 23324
rect 5964 23154 6020 23166
rect 5964 23102 5966 23154
rect 6018 23102 6020 23154
rect 5964 20804 6020 23102
rect 6076 22148 6132 28252
rect 6300 28084 6356 28094
rect 6300 27990 6356 28028
rect 6188 27524 6244 27534
rect 6188 27188 6244 27468
rect 6188 27094 6244 27132
rect 6748 27188 6804 31948
rect 7084 31778 7140 31790
rect 7084 31726 7086 31778
rect 7138 31726 7140 31778
rect 6860 31668 6916 31678
rect 6860 31574 6916 31612
rect 6972 31556 7028 31566
rect 6972 31462 7028 31500
rect 6860 31444 6916 31454
rect 6860 31220 6916 31388
rect 6972 31220 7028 31230
rect 6860 31218 7028 31220
rect 6860 31166 6974 31218
rect 7026 31166 7028 31218
rect 6860 31164 7028 31166
rect 6972 31154 7028 31164
rect 6860 30882 6916 30894
rect 6860 30830 6862 30882
rect 6914 30830 6916 30882
rect 6860 29988 6916 30830
rect 7084 30884 7140 31726
rect 7084 30818 7140 30828
rect 6860 29922 6916 29932
rect 7084 30548 7140 30558
rect 6972 29316 7028 29326
rect 6972 29222 7028 29260
rect 6972 28756 7028 28766
rect 7084 28756 7140 30492
rect 7196 29764 7252 33068
rect 7420 32788 7476 35196
rect 7532 35028 7588 35038
rect 7532 34914 7588 34972
rect 7532 34862 7534 34914
rect 7586 34862 7588 34914
rect 7532 34850 7588 34862
rect 7756 34580 7812 35420
rect 7868 34914 7924 34926
rect 7868 34862 7870 34914
rect 7922 34862 7924 34914
rect 7868 34804 7924 34862
rect 7868 34738 7924 34748
rect 7980 34914 8036 34926
rect 7980 34862 7982 34914
rect 8034 34862 8036 34914
rect 7644 34130 7700 34142
rect 7644 34078 7646 34130
rect 7698 34078 7700 34130
rect 7532 34018 7588 34030
rect 7532 33966 7534 34018
rect 7586 33966 7588 34018
rect 7532 33348 7588 33966
rect 7644 33572 7700 34078
rect 7644 33506 7700 33516
rect 7532 33282 7588 33292
rect 7756 33122 7812 34524
rect 7980 33460 8036 34862
rect 8092 34916 8148 34926
rect 8316 34916 8372 37212
rect 8540 35700 8596 35710
rect 8540 35606 8596 35644
rect 8764 35476 8820 38612
rect 8988 38612 9716 38668
rect 9772 39394 9828 39406
rect 9772 39342 9774 39394
rect 9826 39342 9828 39394
rect 9772 38948 9828 39342
rect 9884 39060 9940 39788
rect 9996 39620 10052 39630
rect 9996 39526 10052 39564
rect 10332 39618 10388 40572
rect 10332 39566 10334 39618
rect 10386 39566 10388 39618
rect 10332 39554 10388 39566
rect 10108 39060 10164 39070
rect 9884 39058 10164 39060
rect 9884 39006 10110 39058
rect 10162 39006 10164 39058
rect 9884 39004 10164 39006
rect 10108 38994 10164 39004
rect 8988 38050 9044 38612
rect 8988 37998 8990 38050
rect 9042 37998 9044 38050
rect 8988 37986 9044 37998
rect 9548 38052 9604 38062
rect 9548 37958 9604 37996
rect 9100 37940 9156 37950
rect 9100 37846 9156 37884
rect 9324 37828 9380 37838
rect 9324 37734 9380 37772
rect 8876 37378 8932 37390
rect 8876 37326 8878 37378
rect 8930 37326 8932 37378
rect 8876 36260 8932 37326
rect 8988 37380 9044 37390
rect 8988 37286 9044 37324
rect 8988 36596 9044 36606
rect 9772 36596 9828 38892
rect 9996 38834 10052 38846
rect 9996 38782 9998 38834
rect 10050 38782 10052 38834
rect 9996 38724 10052 38782
rect 9996 38658 10052 38668
rect 10108 38836 10164 38846
rect 10108 37380 10164 38780
rect 10220 38834 10276 38846
rect 10220 38782 10222 38834
rect 10274 38782 10276 38834
rect 10220 38052 10276 38782
rect 10444 38612 10500 45388
rect 10668 45330 10724 46396
rect 11004 46386 11060 46396
rect 11116 46450 11284 46452
rect 11116 46398 11230 46450
rect 11282 46398 11284 46450
rect 11116 46396 11284 46398
rect 11004 46116 11060 46126
rect 10668 45278 10670 45330
rect 10722 45278 10724 45330
rect 10668 45266 10724 45278
rect 10780 45780 10836 45790
rect 10556 45220 10612 45230
rect 10556 45126 10612 45164
rect 10780 45218 10836 45724
rect 10780 45166 10782 45218
rect 10834 45166 10836 45218
rect 10780 45108 10836 45166
rect 10780 45042 10836 45052
rect 10892 44324 10948 44334
rect 11004 44324 11060 46060
rect 11116 44436 11172 46396
rect 11228 46386 11284 46396
rect 11340 46228 11396 48860
rect 11228 46172 11396 46228
rect 11452 46452 11508 52668
rect 11676 52658 11732 52668
rect 11788 53506 11844 53518
rect 11788 53454 11790 53506
rect 11842 53454 11844 53506
rect 11676 52050 11732 52062
rect 11676 51998 11678 52050
rect 11730 51998 11732 52050
rect 11676 51940 11732 51998
rect 11676 51874 11732 51884
rect 11788 51604 11844 53454
rect 12572 52050 12628 52062
rect 12572 51998 12574 52050
rect 12626 51998 12628 52050
rect 12572 51828 12628 51998
rect 12572 51762 12628 51772
rect 11564 51268 11620 51278
rect 11564 50596 11620 51212
rect 11788 50820 11844 51548
rect 12684 51268 12740 51278
rect 12684 51174 12740 51212
rect 12124 51156 12180 51166
rect 12796 51156 12852 54460
rect 12908 53732 12964 58940
rect 13804 58996 13860 59838
rect 14028 59892 14084 59902
rect 14028 59442 14084 59836
rect 14028 59390 14030 59442
rect 14082 59390 14084 59442
rect 14028 59378 14084 59390
rect 14140 59778 14196 59790
rect 14140 59726 14142 59778
rect 14194 59726 14196 59778
rect 14140 59332 14196 59726
rect 14140 59266 14196 59276
rect 14476 59778 14532 59790
rect 14476 59726 14478 59778
rect 14530 59726 14532 59778
rect 13804 58930 13860 58940
rect 13804 58772 13860 58782
rect 13468 58660 13524 58670
rect 13468 58566 13524 58604
rect 13804 58658 13860 58716
rect 13804 58606 13806 58658
rect 13858 58606 13860 58658
rect 13804 58594 13860 58606
rect 14476 58548 14532 59726
rect 14812 59778 14868 59790
rect 14812 59726 14814 59778
rect 14866 59726 14868 59778
rect 14812 59444 14868 59726
rect 14812 59378 14868 59388
rect 14924 59332 14980 59342
rect 14924 59238 14980 59276
rect 14476 58482 14532 58492
rect 15260 58884 15316 59948
rect 15372 59938 15428 59948
rect 16940 60004 16996 60014
rect 16940 60002 17108 60004
rect 16940 59950 16942 60002
rect 16994 59950 17108 60002
rect 16940 59948 17108 59950
rect 16940 59938 16996 59948
rect 14140 58436 14196 58446
rect 14028 58324 14084 58334
rect 13916 58322 14084 58324
rect 13916 58270 14030 58322
rect 14082 58270 14084 58322
rect 13916 58268 14084 58270
rect 13580 57876 13636 57886
rect 13132 57538 13188 57550
rect 13132 57486 13134 57538
rect 13186 57486 13188 57538
rect 13132 56980 13188 57486
rect 13580 57538 13636 57820
rect 13580 57486 13582 57538
rect 13634 57486 13636 57538
rect 13580 57474 13636 57486
rect 13132 56914 13188 56924
rect 13916 56980 13972 58268
rect 14028 58258 14084 58268
rect 14028 57876 14084 57886
rect 14140 57876 14196 58380
rect 14700 58324 14756 58334
rect 14028 57874 14196 57876
rect 14028 57822 14030 57874
rect 14082 57822 14196 57874
rect 14028 57820 14196 57822
rect 14476 58322 14756 58324
rect 14476 58270 14702 58322
rect 14754 58270 14756 58322
rect 14476 58268 14756 58270
rect 14476 57874 14532 58268
rect 14700 58258 14756 58268
rect 14812 58212 14868 58222
rect 14812 57988 14868 58156
rect 14476 57822 14478 57874
rect 14530 57822 14532 57874
rect 14028 57810 14084 57820
rect 14476 57810 14532 57822
rect 14588 57932 14868 57988
rect 14588 57876 14644 57932
rect 14588 57782 14644 57820
rect 14700 57764 14756 57774
rect 14700 57762 14980 57764
rect 14700 57710 14702 57762
rect 14754 57710 14980 57762
rect 14700 57708 14980 57710
rect 14700 57698 14756 57708
rect 14364 57652 14420 57662
rect 14364 57650 14532 57652
rect 14364 57598 14366 57650
rect 14418 57598 14532 57650
rect 14364 57596 14532 57598
rect 14364 57586 14420 57596
rect 13916 56914 13972 56924
rect 14028 57540 14084 57550
rect 14028 57092 14084 57484
rect 14028 56978 14084 57036
rect 14028 56926 14030 56978
rect 14082 56926 14084 56978
rect 14028 56914 14084 56926
rect 13020 56868 13076 56878
rect 13020 56774 13076 56812
rect 13580 56868 13636 56878
rect 13580 56774 13636 56812
rect 14364 56754 14420 56766
rect 14364 56702 14366 56754
rect 14418 56702 14420 56754
rect 14140 56532 14196 56542
rect 13020 55970 13076 55982
rect 13020 55918 13022 55970
rect 13074 55918 13076 55970
rect 13020 55858 13076 55918
rect 13020 55806 13022 55858
rect 13074 55806 13076 55858
rect 13020 55794 13076 55806
rect 13356 55972 13412 55982
rect 13356 55524 13412 55916
rect 13468 55972 13524 55982
rect 13804 55972 13860 55982
rect 13468 55970 13636 55972
rect 13468 55918 13470 55970
rect 13522 55918 13636 55970
rect 13468 55916 13636 55918
rect 13468 55906 13524 55916
rect 13356 55468 13524 55524
rect 13020 55074 13076 55086
rect 13020 55022 13022 55074
rect 13074 55022 13076 55074
rect 13020 54964 13076 55022
rect 13020 54908 13412 54964
rect 13244 54740 13300 54750
rect 13244 54646 13300 54684
rect 12908 53638 12964 53676
rect 13020 54628 13076 54638
rect 12908 52052 12964 52062
rect 13020 52052 13076 54572
rect 13132 54516 13188 54526
rect 13132 54422 13188 54460
rect 13244 54290 13300 54302
rect 13244 54238 13246 54290
rect 13298 54238 13300 54290
rect 13244 53060 13300 54238
rect 13244 52994 13300 53004
rect 12908 52050 13300 52052
rect 12908 51998 12910 52050
rect 12962 51998 13300 52050
rect 12908 51996 13300 51998
rect 12908 51986 12964 51996
rect 12124 51154 12628 51156
rect 12124 51102 12126 51154
rect 12178 51102 12628 51154
rect 12124 51100 12628 51102
rect 12124 51090 12180 51100
rect 11788 50754 11844 50764
rect 12348 50932 12404 50942
rect 11564 50034 11620 50540
rect 11564 49982 11566 50034
rect 11618 49982 11620 50034
rect 11564 49970 11620 49982
rect 12012 50372 12068 50382
rect 11676 49026 11732 49038
rect 11676 48974 11678 49026
rect 11730 48974 11732 49026
rect 11228 45890 11284 46172
rect 11452 46116 11508 46396
rect 11452 46050 11508 46060
rect 11564 48914 11620 48926
rect 11564 48862 11566 48914
rect 11618 48862 11620 48914
rect 11340 46004 11396 46014
rect 11340 45910 11396 45948
rect 11228 45838 11230 45890
rect 11282 45838 11284 45890
rect 11228 45780 11284 45838
rect 11228 45714 11284 45724
rect 11452 45778 11508 45790
rect 11452 45726 11454 45778
rect 11506 45726 11508 45778
rect 11452 45668 11508 45726
rect 11452 45602 11508 45612
rect 11564 45444 11620 48862
rect 11676 47012 11732 48974
rect 11900 48802 11956 48814
rect 11900 48750 11902 48802
rect 11954 48750 11956 48802
rect 11900 48356 11956 48750
rect 11900 48290 11956 48300
rect 11900 47460 11956 47470
rect 11900 47234 11956 47404
rect 12012 47458 12068 50316
rect 12348 50372 12404 50876
rect 12348 50306 12404 50316
rect 12460 50820 12516 50830
rect 12460 50036 12516 50764
rect 12348 49980 12516 50036
rect 12572 50708 12628 51100
rect 12796 51090 12852 51100
rect 12908 51266 12964 51278
rect 12908 51214 12910 51266
rect 12962 51214 12964 51266
rect 12124 49700 12180 49710
rect 12124 49026 12180 49644
rect 12124 48974 12126 49026
rect 12178 48974 12180 49026
rect 12124 48962 12180 48974
rect 12236 49140 12292 49150
rect 12236 47796 12292 49084
rect 12348 48020 12404 49980
rect 12460 49812 12516 49822
rect 12572 49812 12628 50652
rect 12684 50596 12740 50606
rect 12684 49922 12740 50540
rect 12908 50428 12964 51214
rect 13020 50596 13076 50606
rect 13020 50502 13076 50540
rect 12684 49870 12686 49922
rect 12738 49870 12740 49922
rect 12684 49858 12740 49870
rect 12796 50372 12964 50428
rect 12460 49810 12628 49812
rect 12460 49758 12462 49810
rect 12514 49758 12628 49810
rect 12460 49756 12628 49758
rect 12460 48356 12516 49756
rect 12572 48804 12628 48814
rect 12572 48710 12628 48748
rect 12796 48466 12852 50372
rect 13244 49810 13300 51996
rect 13356 51828 13412 54908
rect 13468 52388 13524 55468
rect 13580 54068 13636 55916
rect 13804 55970 14084 55972
rect 13804 55918 13806 55970
rect 13858 55918 14084 55970
rect 13804 55916 14084 55918
rect 13804 55906 13860 55916
rect 13916 55076 13972 55086
rect 13916 54852 13972 55020
rect 13804 54628 13860 54638
rect 13804 54534 13860 54572
rect 13692 54514 13748 54526
rect 13692 54462 13694 54514
rect 13746 54462 13748 54514
rect 13692 54180 13748 54462
rect 13916 54516 13972 54796
rect 13916 54450 13972 54460
rect 13804 54292 13860 54302
rect 13804 54290 13972 54292
rect 13804 54238 13806 54290
rect 13858 54238 13972 54290
rect 13804 54236 13972 54238
rect 13804 54226 13860 54236
rect 13692 54114 13748 54124
rect 13580 54002 13636 54012
rect 13804 54068 13860 54078
rect 13692 53956 13748 53966
rect 13692 53730 13748 53900
rect 13804 53954 13860 54012
rect 13804 53902 13806 53954
rect 13858 53902 13860 53954
rect 13804 53890 13860 53902
rect 13692 53678 13694 53730
rect 13746 53678 13748 53730
rect 13692 53666 13748 53678
rect 13580 53508 13636 53518
rect 13580 53414 13636 53452
rect 13804 53396 13860 53406
rect 13692 52836 13748 52846
rect 13692 52742 13748 52780
rect 13468 52322 13524 52332
rect 13804 52612 13860 53340
rect 13692 52164 13748 52174
rect 13692 52070 13748 52108
rect 13804 52162 13860 52556
rect 13804 52110 13806 52162
rect 13858 52110 13860 52162
rect 13804 52098 13860 52110
rect 13916 52052 13972 54236
rect 13916 51986 13972 51996
rect 14028 53172 14084 55916
rect 14140 55188 14196 56476
rect 14364 56308 14420 56702
rect 14364 56242 14420 56252
rect 14364 55970 14420 55982
rect 14364 55918 14366 55970
rect 14418 55918 14420 55970
rect 14364 55858 14420 55918
rect 14364 55806 14366 55858
rect 14418 55806 14420 55858
rect 14140 55094 14196 55132
rect 14252 55524 14308 55534
rect 14252 54740 14308 55468
rect 14140 54684 14308 54740
rect 14140 53730 14196 54684
rect 14252 54516 14308 54526
rect 14252 54422 14308 54460
rect 14140 53678 14142 53730
rect 14194 53678 14196 53730
rect 14140 53666 14196 53678
rect 14364 53620 14420 55806
rect 14476 53732 14532 57596
rect 14700 56756 14756 56766
rect 14700 56662 14756 56700
rect 14700 55972 14756 55982
rect 14700 55878 14756 55916
rect 14588 55524 14644 55534
rect 14588 54740 14644 55468
rect 14924 54740 14980 57708
rect 15036 57652 15092 57662
rect 15036 57558 15092 57596
rect 15260 57090 15316 58828
rect 15372 59778 15428 59790
rect 15372 59726 15374 59778
rect 15426 59726 15428 59778
rect 15372 58436 15428 59726
rect 15932 59778 15988 59790
rect 16156 59780 16212 59790
rect 15932 59726 15934 59778
rect 15986 59726 15988 59778
rect 15932 58660 15988 59726
rect 15372 58370 15428 58380
rect 15820 58548 15876 58558
rect 15260 57038 15262 57090
rect 15314 57038 15316 57090
rect 15260 57026 15316 57038
rect 15484 58212 15540 58222
rect 15484 57876 15540 58156
rect 15036 56980 15092 56990
rect 15036 56886 15092 56924
rect 15372 56644 15428 56654
rect 15036 56082 15092 56094
rect 15036 56030 15038 56082
rect 15090 56030 15092 56082
rect 15036 55524 15092 56030
rect 15036 55468 15316 55524
rect 15260 55412 15316 55468
rect 15260 55346 15316 55356
rect 15036 54740 15092 54750
rect 14588 54738 14756 54740
rect 14588 54686 14590 54738
rect 14642 54686 14756 54738
rect 14588 54684 14756 54686
rect 14924 54738 15092 54740
rect 14924 54686 15038 54738
rect 15090 54686 15092 54738
rect 14924 54684 15092 54686
rect 14588 54674 14644 54684
rect 14476 53676 14644 53732
rect 14364 53508 14420 53564
rect 14476 53508 14532 53518
rect 14364 53506 14532 53508
rect 14364 53454 14478 53506
rect 14530 53454 14532 53506
rect 14364 53452 14532 53454
rect 13356 51762 13412 51772
rect 13580 51940 13636 51950
rect 13468 51716 13524 51726
rect 13468 51602 13524 51660
rect 13468 51550 13470 51602
rect 13522 51550 13524 51602
rect 13468 51538 13524 51550
rect 13356 51378 13412 51390
rect 13356 51326 13358 51378
rect 13410 51326 13412 51378
rect 13356 51268 13412 51326
rect 13356 50820 13412 51212
rect 13356 50754 13412 50764
rect 13580 50482 13636 51884
rect 14028 51828 14084 53116
rect 14476 53172 14532 53452
rect 14476 53106 14532 53116
rect 13804 51772 14084 51828
rect 14140 52948 14196 52958
rect 14364 52948 14420 52958
rect 14196 52946 14420 52948
rect 14196 52894 14366 52946
rect 14418 52894 14420 52946
rect 14196 52892 14420 52894
rect 13692 51378 13748 51390
rect 13692 51326 13694 51378
rect 13746 51326 13748 51378
rect 13692 50932 13748 51326
rect 13804 50932 13860 51772
rect 14028 51380 14084 51390
rect 14140 51380 14196 52892
rect 14364 52882 14420 52892
rect 14588 52724 14644 53676
rect 14700 53508 14756 54684
rect 15036 54674 15092 54684
rect 15372 54514 15428 56588
rect 15484 56084 15540 57820
rect 15708 57762 15764 57774
rect 15708 57710 15710 57762
rect 15762 57710 15764 57762
rect 15596 57092 15652 57102
rect 15596 56998 15652 57036
rect 15708 56532 15764 57710
rect 15708 56466 15764 56476
rect 15820 56980 15876 58492
rect 15932 57652 15988 58604
rect 16044 59778 16212 59780
rect 16044 59726 16158 59778
rect 16210 59726 16212 59778
rect 16044 59724 16212 59726
rect 16044 58436 16100 59724
rect 16156 59714 16212 59724
rect 16268 59778 16324 59790
rect 16268 59726 16270 59778
rect 16322 59726 16324 59778
rect 16044 58370 16100 58380
rect 16156 59444 16212 59454
rect 16156 57762 16212 59388
rect 16268 59108 16324 59726
rect 16268 59042 16324 59052
rect 16380 59778 16436 59790
rect 16380 59726 16382 59778
rect 16434 59726 16436 59778
rect 16380 57988 16436 59726
rect 16940 59106 16996 59118
rect 16940 59054 16942 59106
rect 16994 59054 16996 59106
rect 16380 57922 16436 57932
rect 16492 58210 16548 58222
rect 16492 58158 16494 58210
rect 16546 58158 16548 58210
rect 16156 57710 16158 57762
rect 16210 57710 16212 57762
rect 16156 57698 16212 57710
rect 15932 57586 15988 57596
rect 16380 57652 16436 57662
rect 16492 57652 16548 58158
rect 16940 58212 16996 59054
rect 16940 57764 16996 58156
rect 16940 57698 16996 57708
rect 16380 57650 16548 57652
rect 16380 57598 16382 57650
rect 16434 57598 16548 57650
rect 16380 57596 16548 57598
rect 16156 57204 16212 57214
rect 15820 56924 16100 56980
rect 15596 56308 15652 56318
rect 15596 56214 15652 56252
rect 15484 56028 15652 56084
rect 15484 55412 15540 55422
rect 15484 55318 15540 55356
rect 15372 54462 15374 54514
rect 15426 54462 15428 54514
rect 15372 54450 15428 54462
rect 15484 55188 15540 55198
rect 14812 54404 14868 54414
rect 14812 53730 14868 54348
rect 15484 53956 15540 55132
rect 15372 53900 15540 53956
rect 14812 53678 14814 53730
rect 14866 53678 14868 53730
rect 14812 53666 14868 53678
rect 15148 53730 15204 53742
rect 15148 53678 15150 53730
rect 15202 53678 15204 53730
rect 14700 53452 14980 53508
rect 14364 52668 14644 52724
rect 14700 53284 14756 53294
rect 14252 52276 14308 52286
rect 14252 51938 14308 52220
rect 14364 52274 14420 52668
rect 14364 52222 14366 52274
rect 14418 52222 14420 52274
rect 14364 52210 14420 52222
rect 14476 52388 14532 52398
rect 14252 51886 14254 51938
rect 14306 51886 14308 51938
rect 14252 51604 14308 51886
rect 14476 52050 14532 52332
rect 14700 52164 14756 53228
rect 14700 52098 14756 52108
rect 14812 52948 14868 52958
rect 14812 52724 14868 52892
rect 14476 51998 14478 52050
rect 14530 51998 14532 52050
rect 14476 51940 14532 51998
rect 14476 51874 14532 51884
rect 14812 51604 14868 52668
rect 14252 51538 14308 51548
rect 14476 51548 14868 51604
rect 14028 51378 14196 51380
rect 14028 51326 14030 51378
rect 14082 51326 14196 51378
rect 14028 51324 14196 51326
rect 14028 51314 14084 51324
rect 13804 50876 13972 50932
rect 13692 50866 13748 50876
rect 13804 50708 13860 50718
rect 13804 50594 13860 50652
rect 13804 50542 13806 50594
rect 13858 50542 13860 50594
rect 13804 50530 13860 50542
rect 13580 50430 13582 50482
rect 13634 50430 13636 50482
rect 13580 50418 13636 50430
rect 13916 50428 13972 50876
rect 14364 50596 14420 50606
rect 14364 50502 14420 50540
rect 13804 50372 13972 50428
rect 13804 49924 13860 50372
rect 14476 50260 14532 51548
rect 14700 51268 14756 51278
rect 14700 51174 14756 51212
rect 14700 50372 14756 50382
rect 13916 50204 14532 50260
rect 14588 50370 14756 50372
rect 14588 50318 14702 50370
rect 14754 50318 14756 50370
rect 14588 50316 14756 50318
rect 13916 50036 13972 50204
rect 13916 49980 14084 50036
rect 13804 49858 13860 49868
rect 13244 49758 13246 49810
rect 13298 49758 13300 49810
rect 13244 49746 13300 49758
rect 13916 49810 13972 49822
rect 13916 49758 13918 49810
rect 13970 49758 13972 49810
rect 13580 49588 13636 49598
rect 13916 49588 13972 49758
rect 13580 49586 13860 49588
rect 13580 49534 13582 49586
rect 13634 49534 13860 49586
rect 13580 49532 13860 49534
rect 13580 49522 13636 49532
rect 13804 49028 13860 49532
rect 13916 49252 13972 49532
rect 13916 49186 13972 49196
rect 13804 48972 13972 49028
rect 12908 48916 12964 48926
rect 12908 48822 12964 48860
rect 13804 48804 13860 48814
rect 12796 48414 12798 48466
rect 12850 48414 12852 48466
rect 12460 48300 12628 48356
rect 12348 47954 12404 47964
rect 12460 48018 12516 48030
rect 12460 47966 12462 48018
rect 12514 47966 12516 48018
rect 12460 47796 12516 47966
rect 12012 47406 12014 47458
rect 12066 47406 12068 47458
rect 12012 47394 12068 47406
rect 12124 47740 12516 47796
rect 11900 47182 11902 47234
rect 11954 47182 11956 47234
rect 11900 47170 11956 47182
rect 12124 47012 12180 47740
rect 11676 46946 11732 46956
rect 11788 46956 12180 47012
rect 11788 46786 11844 46956
rect 11788 46734 11790 46786
rect 11842 46734 11844 46786
rect 11788 46676 11844 46734
rect 11788 46610 11844 46620
rect 12012 46450 12068 46462
rect 12012 46398 12014 46450
rect 12066 46398 12068 46450
rect 11788 46116 11844 46126
rect 11788 46114 11956 46116
rect 11788 46062 11790 46114
rect 11842 46062 11956 46114
rect 11788 46060 11956 46062
rect 11788 46050 11844 46060
rect 11676 46004 11732 46014
rect 11676 45892 11732 45948
rect 11788 45892 11844 45902
rect 11676 45890 11844 45892
rect 11676 45838 11790 45890
rect 11842 45838 11844 45890
rect 11676 45836 11844 45838
rect 11788 45826 11844 45836
rect 11228 45388 11620 45444
rect 11788 45668 11844 45678
rect 11228 45330 11284 45388
rect 11228 45278 11230 45330
rect 11282 45278 11284 45330
rect 11228 45266 11284 45278
rect 11564 45108 11620 45118
rect 11564 44884 11620 45052
rect 11564 44818 11620 44828
rect 11340 44436 11396 44446
rect 11788 44436 11844 45612
rect 11116 44380 11284 44436
rect 11004 44268 11172 44324
rect 10892 44230 10948 44268
rect 11004 43540 11060 43550
rect 11004 43446 11060 43484
rect 10556 42756 10612 42766
rect 10556 42662 10612 42700
rect 10780 42082 10836 42094
rect 10780 42030 10782 42082
rect 10834 42030 10836 42082
rect 10780 41860 10836 42030
rect 10780 41076 10836 41804
rect 11116 41748 11172 44268
rect 11228 43650 11284 44380
rect 11228 43598 11230 43650
rect 11282 43598 11284 43650
rect 11228 43586 11284 43598
rect 11340 43650 11396 44380
rect 11340 43598 11342 43650
rect 11394 43598 11396 43650
rect 11340 43586 11396 43598
rect 11676 44380 11844 44436
rect 11676 43540 11732 44380
rect 11676 43446 11732 43484
rect 11788 44210 11844 44222
rect 11788 44158 11790 44210
rect 11842 44158 11844 44210
rect 11788 43316 11844 44158
rect 11900 43764 11956 46060
rect 12012 45668 12068 46398
rect 12348 46452 12404 46462
rect 12348 46450 12516 46452
rect 12348 46398 12350 46450
rect 12402 46398 12516 46450
rect 12348 46396 12516 46398
rect 12348 46386 12404 46396
rect 12012 45602 12068 45612
rect 12348 45890 12404 45902
rect 12348 45838 12350 45890
rect 12402 45838 12404 45890
rect 12236 45218 12292 45230
rect 12236 45166 12238 45218
rect 12290 45166 12292 45218
rect 12236 44436 12292 45166
rect 12348 45220 12404 45838
rect 12348 45106 12404 45164
rect 12348 45054 12350 45106
rect 12402 45054 12404 45106
rect 12348 45042 12404 45054
rect 12236 44342 12292 44380
rect 12124 44322 12180 44334
rect 12124 44270 12126 44322
rect 12178 44270 12180 44322
rect 12012 43764 12068 43774
rect 11900 43762 12068 43764
rect 11900 43710 12014 43762
rect 12066 43710 12068 43762
rect 11900 43708 12068 43710
rect 12012 43698 12068 43708
rect 12124 43540 12180 44270
rect 12348 44210 12404 44222
rect 12348 44158 12350 44210
rect 12402 44158 12404 44210
rect 12236 43540 12292 43550
rect 12124 43538 12292 43540
rect 12124 43486 12238 43538
rect 12290 43486 12292 43538
rect 12124 43484 12292 43486
rect 12348 43540 12404 44158
rect 12460 43764 12516 46396
rect 12572 46004 12628 48300
rect 12796 48244 12852 48414
rect 13468 48802 13860 48804
rect 13468 48750 13806 48802
rect 13858 48750 13860 48802
rect 13468 48748 13860 48750
rect 13132 48356 13188 48366
rect 12684 47460 12740 47470
rect 12684 47366 12740 47404
rect 12796 47346 12852 48188
rect 12796 47294 12798 47346
rect 12850 47294 12852 47346
rect 12796 47282 12852 47294
rect 12908 48300 13132 48356
rect 12796 46900 12852 46910
rect 12908 46900 12964 48300
rect 13132 48262 13188 48300
rect 13468 47684 13524 48748
rect 13804 48738 13860 48748
rect 13244 47628 13524 47684
rect 13580 48580 13636 48590
rect 13580 48242 13636 48524
rect 13580 48190 13582 48242
rect 13634 48190 13636 48242
rect 13132 47012 13188 47022
rect 12796 46898 12964 46900
rect 12796 46846 12798 46898
rect 12850 46846 12964 46898
rect 12796 46844 12964 46846
rect 13020 46900 13076 46910
rect 12796 46834 12852 46844
rect 13020 46806 13076 46844
rect 13132 46898 13188 46956
rect 13132 46846 13134 46898
rect 13186 46846 13188 46898
rect 13132 46834 13188 46846
rect 13244 46898 13300 47628
rect 13580 47572 13636 48190
rect 13468 47516 13636 47572
rect 13468 47460 13524 47516
rect 13468 47394 13524 47404
rect 13580 47346 13636 47358
rect 13580 47294 13582 47346
rect 13634 47294 13636 47346
rect 13468 47236 13524 47246
rect 13468 47142 13524 47180
rect 13580 47012 13636 47294
rect 13244 46846 13246 46898
rect 13298 46846 13300 46898
rect 13244 46834 13300 46846
rect 13356 46956 13636 47012
rect 13804 47348 13860 47358
rect 12572 45938 12628 45948
rect 13020 46004 13076 46014
rect 13356 46004 13412 46956
rect 13804 46674 13860 47292
rect 13804 46622 13806 46674
rect 13858 46622 13860 46674
rect 13804 46610 13860 46622
rect 13916 46116 13972 48972
rect 14028 47684 14084 49980
rect 14140 49924 14196 49934
rect 14140 49026 14196 49868
rect 14364 49812 14420 49822
rect 14140 48974 14142 49026
rect 14194 48974 14196 49026
rect 14140 47908 14196 48974
rect 14140 47842 14196 47852
rect 14252 49810 14420 49812
rect 14252 49758 14366 49810
rect 14418 49758 14420 49810
rect 14252 49756 14420 49758
rect 14252 48356 14308 49756
rect 14364 49746 14420 49756
rect 14588 49810 14644 50316
rect 14700 50306 14756 50316
rect 14588 49758 14590 49810
rect 14642 49758 14644 49810
rect 14476 49700 14532 49710
rect 14476 49606 14532 49644
rect 14028 47628 14196 47684
rect 14028 47458 14084 47470
rect 14028 47406 14030 47458
rect 14082 47406 14084 47458
rect 14028 46900 14084 47406
rect 14028 46562 14084 46844
rect 14028 46510 14030 46562
rect 14082 46510 14084 46562
rect 14028 46498 14084 46510
rect 14140 46564 14196 47628
rect 14252 47458 14308 48300
rect 14252 47406 14254 47458
rect 14306 47406 14308 47458
rect 14252 47394 14308 47406
rect 14364 49026 14420 49038
rect 14364 48974 14366 49026
rect 14418 48974 14420 49026
rect 14364 48916 14420 48974
rect 14364 47348 14420 48860
rect 14588 48580 14644 49758
rect 14812 49700 14868 49710
rect 14812 48914 14868 49644
rect 14812 48862 14814 48914
rect 14866 48862 14868 48914
rect 14812 48850 14868 48862
rect 14588 48514 14644 48524
rect 14700 48244 14756 48254
rect 14700 48150 14756 48188
rect 14364 47282 14420 47292
rect 14700 47346 14756 47358
rect 14700 47294 14702 47346
rect 14754 47294 14756 47346
rect 14700 47124 14756 47294
rect 14700 47058 14756 47068
rect 14476 46900 14532 46910
rect 14476 46786 14532 46844
rect 14476 46734 14478 46786
rect 14530 46734 14532 46786
rect 14476 46722 14532 46734
rect 14700 46676 14756 46686
rect 14700 46582 14756 46620
rect 14252 46564 14308 46574
rect 14140 46508 14252 46564
rect 14252 46498 14308 46508
rect 13076 45948 13412 46004
rect 13580 46060 13916 46116
rect 13020 45938 13076 45948
rect 13468 45892 13524 45902
rect 13468 45798 13524 45836
rect 12908 45780 12964 45790
rect 12964 45724 13188 45780
rect 12908 45686 12964 45724
rect 12796 45668 12852 45678
rect 12796 45330 12852 45612
rect 12796 45278 12798 45330
rect 12850 45278 12852 45330
rect 12796 45266 12852 45278
rect 13020 45556 13076 45566
rect 13020 45106 13076 45500
rect 13020 45054 13022 45106
rect 13074 45054 13076 45106
rect 12908 44098 12964 44110
rect 12908 44046 12910 44098
rect 12962 44046 12964 44098
rect 12908 43876 12964 44046
rect 12460 43698 12516 43708
rect 12796 43820 12964 43876
rect 12796 43652 12852 43820
rect 12796 43586 12852 43596
rect 12908 43652 12964 43662
rect 13020 43652 13076 45054
rect 12908 43650 13076 43652
rect 12908 43598 12910 43650
rect 12962 43598 13076 43650
rect 12908 43596 13076 43598
rect 12908 43586 12964 43596
rect 12460 43540 12516 43550
rect 13132 43540 13188 45724
rect 13580 45106 13636 46060
rect 13916 46022 13972 46060
rect 14252 46116 14308 46126
rect 14308 46060 14420 46116
rect 14252 46050 14308 46060
rect 14364 45892 14420 46060
rect 14364 45890 14868 45892
rect 14364 45838 14366 45890
rect 14418 45838 14868 45890
rect 14364 45836 14868 45838
rect 14364 45826 14420 45836
rect 14252 45778 14308 45790
rect 14252 45726 14254 45778
rect 14306 45726 14308 45778
rect 14028 45444 14084 45454
rect 13580 45054 13582 45106
rect 13634 45054 13636 45106
rect 13580 45042 13636 45054
rect 13804 45332 13860 45342
rect 13804 44322 13860 45276
rect 13804 44270 13806 44322
rect 13858 44270 13860 44322
rect 13804 44258 13860 44270
rect 12348 43538 12516 43540
rect 12348 43486 12462 43538
rect 12514 43486 12516 43538
rect 12348 43484 12516 43486
rect 12012 43316 12068 43326
rect 11788 43314 12068 43316
rect 11788 43262 12014 43314
rect 12066 43262 12068 43314
rect 11788 43260 12068 43262
rect 12012 42868 12068 43260
rect 12236 43092 12292 43484
rect 12460 43204 12516 43484
rect 13020 43484 13188 43540
rect 13692 43538 13748 43550
rect 13692 43486 13694 43538
rect 13746 43486 13748 43538
rect 12796 43428 12852 43438
rect 13020 43428 13076 43484
rect 12796 43426 13076 43428
rect 12796 43374 12798 43426
rect 12850 43374 13076 43426
rect 12796 43372 13076 43374
rect 13468 43426 13524 43438
rect 13468 43374 13470 43426
rect 13522 43374 13524 43426
rect 12796 43362 12852 43372
rect 12460 43148 13412 43204
rect 12236 43036 12628 43092
rect 12460 42868 12516 42878
rect 12012 42866 12516 42868
rect 12012 42814 12462 42866
rect 12514 42814 12516 42866
rect 12012 42812 12516 42814
rect 12460 42802 12516 42812
rect 12012 42644 12068 42654
rect 12012 42194 12068 42588
rect 12348 42642 12404 42654
rect 12348 42590 12350 42642
rect 12402 42590 12404 42642
rect 12012 42142 12014 42194
rect 12066 42142 12068 42194
rect 12012 42130 12068 42142
rect 12124 42530 12180 42542
rect 12124 42478 12126 42530
rect 12178 42478 12180 42530
rect 12012 41972 12068 41982
rect 11228 41748 11284 41758
rect 11116 41692 11228 41748
rect 11228 41682 11284 41692
rect 11900 41748 11956 41758
rect 11788 41188 11844 41198
rect 10668 41074 10836 41076
rect 10668 41022 10782 41074
rect 10834 41022 10836 41074
rect 10668 41020 10836 41022
rect 10556 38836 10612 38846
rect 10668 38836 10724 41020
rect 10780 41010 10836 41020
rect 11340 41076 11396 41086
rect 11340 40404 11396 41020
rect 11340 40338 11396 40348
rect 11452 40290 11508 40302
rect 11452 40238 11454 40290
rect 11506 40238 11508 40290
rect 11004 40180 11060 40190
rect 10892 40178 11060 40180
rect 10892 40126 11006 40178
rect 11058 40126 11060 40178
rect 10892 40124 11060 40126
rect 10612 38780 10724 38836
rect 10780 39394 10836 39406
rect 10780 39342 10782 39394
rect 10834 39342 10836 39394
rect 10780 38836 10836 39342
rect 10556 38770 10612 38780
rect 10780 38770 10836 38780
rect 10444 38556 10612 38612
rect 10444 38052 10500 38062
rect 10220 38050 10500 38052
rect 10220 37998 10446 38050
rect 10498 37998 10500 38050
rect 10220 37996 10500 37998
rect 10220 37716 10276 37996
rect 10444 37986 10500 37996
rect 10220 37650 10276 37660
rect 10220 37380 10276 37390
rect 10108 37378 10276 37380
rect 10108 37326 10222 37378
rect 10274 37326 10276 37378
rect 10108 37324 10276 37326
rect 8988 36594 9828 36596
rect 8988 36542 8990 36594
rect 9042 36542 9828 36594
rect 8988 36540 9828 36542
rect 9884 37044 9940 37054
rect 8988 36530 9044 36540
rect 9212 36372 9268 36382
rect 9884 36372 9940 36988
rect 9212 36370 9940 36372
rect 9212 36318 9214 36370
rect 9266 36318 9940 36370
rect 9212 36316 9940 36318
rect 10108 36484 10164 36494
rect 9212 36306 9268 36316
rect 8876 36194 8932 36204
rect 8876 35924 8932 35934
rect 8876 35830 8932 35868
rect 10108 35810 10164 36428
rect 10108 35758 10110 35810
rect 10162 35758 10164 35810
rect 10108 35746 10164 35758
rect 9772 35700 9828 35710
rect 9548 35644 9772 35700
rect 8764 35420 8932 35476
rect 8652 34916 8708 34926
rect 8148 34860 8260 34916
rect 8316 34860 8484 34916
rect 8092 34822 8148 34860
rect 8204 33796 8260 34860
rect 8316 34692 8372 34702
rect 8316 34598 8372 34636
rect 8428 34468 8484 34860
rect 8652 34822 8708 34860
rect 8092 33460 8148 33470
rect 7980 33404 8092 33460
rect 8092 33394 8148 33404
rect 8204 33236 8260 33740
rect 7980 33180 8260 33236
rect 8316 34412 8484 34468
rect 8540 34804 8596 34814
rect 7756 33070 7758 33122
rect 7810 33070 7812 33122
rect 7756 33058 7812 33070
rect 7868 33124 7924 33134
rect 7420 32732 7700 32788
rect 7532 32562 7588 32574
rect 7532 32510 7534 32562
rect 7586 32510 7588 32562
rect 7420 31666 7476 31678
rect 7420 31614 7422 31666
rect 7474 31614 7476 31666
rect 7420 31556 7476 31614
rect 7420 31490 7476 31500
rect 7532 30996 7588 32510
rect 7532 30930 7588 30940
rect 7644 31218 7700 32732
rect 7756 31668 7812 31678
rect 7756 31574 7812 31612
rect 7868 31444 7924 33068
rect 7980 31778 8036 33180
rect 8316 32004 8372 34412
rect 8428 34020 8484 34030
rect 8428 32228 8484 33964
rect 8540 33236 8596 34748
rect 8540 32450 8596 33180
rect 8652 34692 8708 34702
rect 8652 32788 8708 34636
rect 8764 34690 8820 34702
rect 8764 34638 8766 34690
rect 8818 34638 8820 34690
rect 8764 33348 8820 34638
rect 8876 34020 8932 35420
rect 9100 34914 9156 34926
rect 9100 34862 9102 34914
rect 9154 34862 9156 34914
rect 9100 34580 9156 34862
rect 9324 34916 9380 34926
rect 9548 34916 9604 35644
rect 9772 35606 9828 35644
rect 9324 34914 9604 34916
rect 9324 34862 9326 34914
rect 9378 34862 9604 34914
rect 9324 34860 9604 34862
rect 9660 34916 9716 34926
rect 9324 34850 9380 34860
rect 9100 34514 9156 34524
rect 8988 34020 9044 34030
rect 8876 34018 9044 34020
rect 8876 33966 8990 34018
rect 9042 33966 9044 34018
rect 8876 33964 9044 33966
rect 8988 33908 9044 33964
rect 8988 33842 9044 33852
rect 8764 33282 8820 33292
rect 9436 33796 9492 34860
rect 9660 34822 9716 34860
rect 9996 34916 10052 34926
rect 9996 34822 10052 34860
rect 10108 34690 10164 34702
rect 10108 34638 10110 34690
rect 10162 34638 10164 34690
rect 9660 33906 9716 33918
rect 9660 33854 9662 33906
rect 9714 33854 9716 33906
rect 9660 33796 9716 33854
rect 9436 33740 9716 33796
rect 9996 33796 10052 33806
rect 8988 32788 9044 32798
rect 9436 32788 9492 33740
rect 8652 32732 8932 32788
rect 8876 32564 8932 32732
rect 8988 32786 9492 32788
rect 8988 32734 8990 32786
rect 9042 32734 9492 32786
rect 8988 32732 9492 32734
rect 9548 33234 9604 33246
rect 9548 33182 9550 33234
rect 9602 33182 9604 33234
rect 9548 32788 9604 33182
rect 9884 32788 9940 32798
rect 9548 32786 9940 32788
rect 9548 32734 9886 32786
rect 9938 32734 9940 32786
rect 9548 32732 9940 32734
rect 8988 32722 9044 32732
rect 9884 32722 9940 32732
rect 9548 32564 9604 32574
rect 8876 32562 9604 32564
rect 8876 32510 9550 32562
rect 9602 32510 9604 32562
rect 8876 32508 9604 32510
rect 9548 32498 9604 32508
rect 9884 32564 9940 32574
rect 9996 32564 10052 33740
rect 10108 32676 10164 34638
rect 10220 34356 10276 37324
rect 10444 35586 10500 35598
rect 10444 35534 10446 35586
rect 10498 35534 10500 35586
rect 10444 34580 10500 35534
rect 10444 34514 10500 34524
rect 10556 35140 10612 38556
rect 10780 35812 10836 35822
rect 10668 35700 10724 35710
rect 10668 35606 10724 35644
rect 10220 34290 10276 34300
rect 10556 34132 10612 35084
rect 10556 34066 10612 34076
rect 10780 34242 10836 35756
rect 10892 35308 10948 40124
rect 11004 40114 11060 40124
rect 11004 39620 11060 39630
rect 11004 39526 11060 39564
rect 11452 39620 11508 40238
rect 11788 39732 11844 41132
rect 11788 39666 11844 39676
rect 11452 39526 11508 39564
rect 11116 38946 11172 38958
rect 11116 38894 11118 38946
rect 11170 38894 11172 38946
rect 11004 38724 11060 38734
rect 11004 38050 11060 38668
rect 11004 37998 11006 38050
rect 11058 37998 11060 38050
rect 11004 37986 11060 37998
rect 11116 37716 11172 38894
rect 11228 38836 11284 38846
rect 11228 38742 11284 38780
rect 11788 38836 11844 38846
rect 11676 38724 11732 38762
rect 11676 38658 11732 38668
rect 11676 38162 11732 38174
rect 11676 38110 11678 38162
rect 11730 38110 11732 38162
rect 11116 37650 11172 37660
rect 11452 37716 11508 37726
rect 11340 37044 11396 37054
rect 11340 36950 11396 36988
rect 11004 36484 11060 36494
rect 11004 36390 11060 36428
rect 11228 36482 11284 36494
rect 11228 36430 11230 36482
rect 11282 36430 11284 36482
rect 11004 35922 11060 35934
rect 11004 35870 11006 35922
rect 11058 35870 11060 35922
rect 11004 35812 11060 35870
rect 11004 35746 11060 35756
rect 11228 35924 11284 36430
rect 11228 35700 11284 35868
rect 11452 35922 11508 37660
rect 11452 35870 11454 35922
rect 11506 35870 11508 35922
rect 11452 35858 11508 35870
rect 11564 36484 11620 36494
rect 11340 35700 11396 35710
rect 11228 35698 11396 35700
rect 11228 35646 11342 35698
rect 11394 35646 11396 35698
rect 11228 35644 11396 35646
rect 10892 35252 11060 35308
rect 10780 34190 10782 34242
rect 10834 34190 10836 34242
rect 10780 33684 10836 34190
rect 10444 33628 10836 33684
rect 11004 35028 11060 35252
rect 10220 33348 10276 33358
rect 10220 33254 10276 33292
rect 10220 33124 10276 33134
rect 10220 33030 10276 33068
rect 10108 32610 10164 32620
rect 10332 33012 10388 33022
rect 9884 32562 10052 32564
rect 9884 32510 9886 32562
rect 9938 32510 10052 32562
rect 9884 32508 10052 32510
rect 10220 32562 10276 32574
rect 10220 32510 10222 32562
rect 10274 32510 10276 32562
rect 9884 32498 9940 32508
rect 8540 32398 8542 32450
rect 8594 32398 8596 32450
rect 8540 32386 8596 32398
rect 8428 32172 8596 32228
rect 8540 32004 8596 32172
rect 8316 31948 8484 32004
rect 7980 31726 7982 31778
rect 8034 31726 8036 31778
rect 7980 31714 8036 31726
rect 8316 31778 8372 31790
rect 8316 31726 8318 31778
rect 8370 31726 8372 31778
rect 8092 31668 8148 31678
rect 8092 31666 8260 31668
rect 8092 31614 8094 31666
rect 8146 31614 8260 31666
rect 8092 31612 8260 31614
rect 8092 31602 8148 31612
rect 7868 31388 8148 31444
rect 7644 31166 7646 31218
rect 7698 31166 7700 31218
rect 7644 30772 7700 31166
rect 7980 31220 8036 31230
rect 7868 30996 7924 31006
rect 7644 30706 7700 30716
rect 7756 30882 7812 30894
rect 7756 30830 7758 30882
rect 7810 30830 7812 30882
rect 7756 30548 7812 30830
rect 7756 30482 7812 30492
rect 7868 30324 7924 30940
rect 7868 30258 7924 30268
rect 7308 30212 7364 30222
rect 7308 30118 7364 30156
rect 7756 30210 7812 30222
rect 7756 30158 7758 30210
rect 7810 30158 7812 30210
rect 7420 30100 7476 30110
rect 7420 30006 7476 30044
rect 7196 29698 7252 29708
rect 7756 29764 7812 30158
rect 7756 29698 7812 29708
rect 7980 29650 8036 31164
rect 8092 30994 8148 31388
rect 8092 30942 8094 30994
rect 8146 30942 8148 30994
rect 8092 30930 8148 30942
rect 8204 30996 8260 31612
rect 8316 31220 8372 31726
rect 8316 31154 8372 31164
rect 8316 30996 8372 31006
rect 8204 30994 8372 30996
rect 8204 30942 8318 30994
rect 8370 30942 8372 30994
rect 8204 30940 8372 30942
rect 8316 30930 8372 30940
rect 7980 29598 7982 29650
rect 8034 29598 8036 29650
rect 7980 29586 8036 29598
rect 8092 30772 8148 30782
rect 7868 29538 7924 29550
rect 7868 29486 7870 29538
rect 7922 29486 7924 29538
rect 6972 28754 7140 28756
rect 6972 28702 6974 28754
rect 7026 28702 7140 28754
rect 6972 28700 7140 28702
rect 7756 29426 7812 29438
rect 7756 29374 7758 29426
rect 7810 29374 7812 29426
rect 6972 28690 7028 28700
rect 7644 28644 7700 28654
rect 7644 28082 7700 28588
rect 7644 28030 7646 28082
rect 7698 28030 7700 28082
rect 7644 28018 7700 28030
rect 7756 27748 7812 29374
rect 6748 27122 6804 27132
rect 7644 27692 7812 27748
rect 6972 27074 7028 27086
rect 6972 27022 6974 27074
rect 7026 27022 7028 27074
rect 6748 26962 6804 26974
rect 6748 26910 6750 26962
rect 6802 26910 6804 26962
rect 6748 26852 6804 26910
rect 6972 26964 7028 27022
rect 7644 27074 7700 27692
rect 7756 27188 7812 27198
rect 7756 27094 7812 27132
rect 7644 27022 7646 27074
rect 7698 27022 7700 27074
rect 6972 26898 7028 26908
rect 7308 26962 7364 26974
rect 7308 26910 7310 26962
rect 7362 26910 7364 26962
rect 6748 26786 6804 26796
rect 6860 26850 6916 26862
rect 6860 26798 6862 26850
rect 6914 26798 6916 26850
rect 6860 26516 6916 26798
rect 6300 26460 6916 26516
rect 6188 26066 6244 26078
rect 6188 26014 6190 26066
rect 6242 26014 6244 26066
rect 6188 23156 6244 26014
rect 6300 23826 6356 26460
rect 6748 26292 6804 26302
rect 6636 26236 6748 26292
rect 6412 26180 6468 26190
rect 6412 25506 6468 26124
rect 6412 25454 6414 25506
rect 6466 25454 6468 25506
rect 6412 25442 6468 25454
rect 6412 24948 6468 24958
rect 6412 24946 6580 24948
rect 6412 24894 6414 24946
rect 6466 24894 6580 24946
rect 6412 24892 6580 24894
rect 6412 24882 6468 24892
rect 6524 24162 6580 24892
rect 6636 24722 6692 26236
rect 6748 26198 6804 26236
rect 6860 26292 6916 26302
rect 7308 26292 7364 26910
rect 7644 26516 7700 27022
rect 7868 27076 7924 29486
rect 8092 27636 8148 30716
rect 8428 29426 8484 31948
rect 8540 31890 8596 31948
rect 9660 32116 9716 32126
rect 8540 31838 8542 31890
rect 8594 31838 8596 31890
rect 8540 31826 8596 31838
rect 9212 31892 9268 31902
rect 9212 31798 9268 31836
rect 8988 31780 9044 31790
rect 8988 31686 9044 31724
rect 9436 31778 9492 31790
rect 9436 31726 9438 31778
rect 9490 31726 9492 31778
rect 9100 31556 9156 31566
rect 9100 31462 9156 31500
rect 9436 31556 9492 31726
rect 9436 31490 9492 31500
rect 8764 31444 8820 31454
rect 8540 31332 8596 31342
rect 8540 31218 8596 31276
rect 8540 31166 8542 31218
rect 8594 31166 8596 31218
rect 8540 31154 8596 31166
rect 8764 31218 8820 31388
rect 9660 31332 9716 32060
rect 9772 32004 9828 32014
rect 9828 31948 9940 32004
rect 9772 31938 9828 31948
rect 9884 31890 9940 31948
rect 10220 32002 10276 32510
rect 10220 31950 10222 32002
rect 10274 31950 10276 32002
rect 10220 31938 10276 31950
rect 9884 31838 9886 31890
rect 9938 31838 9940 31890
rect 9884 31826 9940 31838
rect 9660 31266 9716 31276
rect 9772 31780 9828 31790
rect 10332 31780 10388 32956
rect 8764 31166 8766 31218
rect 8818 31166 8820 31218
rect 8764 31154 8820 31166
rect 9772 31108 9828 31724
rect 10220 31724 10388 31780
rect 10108 31554 10164 31566
rect 10108 31502 10110 31554
rect 10162 31502 10164 31554
rect 10108 31220 10164 31502
rect 10108 31154 10164 31164
rect 9660 31052 9828 31108
rect 8876 30996 8932 31006
rect 8876 30902 8932 30940
rect 8540 30100 8596 30110
rect 8540 30006 8596 30044
rect 8428 29374 8430 29426
rect 8482 29374 8484 29426
rect 8428 28084 8484 29374
rect 8428 28018 8484 28028
rect 8988 29426 9044 29438
rect 9548 29428 9604 29438
rect 8988 29374 8990 29426
rect 9042 29374 9044 29426
rect 8092 27188 8148 27580
rect 8092 27122 8148 27132
rect 7868 26982 7924 27020
rect 8204 26964 8260 27002
rect 8204 26898 8260 26908
rect 8988 26964 9044 29374
rect 9100 29426 9604 29428
rect 9100 29374 9550 29426
rect 9602 29374 9604 29426
rect 9100 29372 9604 29374
rect 9100 28754 9156 29372
rect 9548 29362 9604 29372
rect 9100 28702 9102 28754
rect 9154 28702 9156 28754
rect 9100 28690 9156 28702
rect 9548 29204 9604 29214
rect 9436 28644 9492 28654
rect 9436 28530 9492 28588
rect 9436 28478 9438 28530
rect 9490 28478 9492 28530
rect 9436 28466 9492 28478
rect 9548 28196 9604 29148
rect 9436 28140 9604 28196
rect 9100 27746 9156 27758
rect 9100 27694 9102 27746
rect 9154 27694 9156 27746
rect 9100 27300 9156 27694
rect 9324 27300 9380 27310
rect 9100 27244 9324 27300
rect 9324 27186 9380 27244
rect 9324 27134 9326 27186
rect 9378 27134 9380 27186
rect 9324 27122 9380 27134
rect 8988 26898 9044 26908
rect 8540 26850 8596 26862
rect 8540 26798 8542 26850
rect 8594 26798 8596 26850
rect 8540 26516 8596 26798
rect 7644 26460 8372 26516
rect 6860 26290 7364 26292
rect 6860 26238 6862 26290
rect 6914 26238 7310 26290
rect 7362 26238 7364 26290
rect 6860 26236 7364 26238
rect 6860 26226 6916 26236
rect 7308 26226 7364 26236
rect 7756 26292 7812 26302
rect 7420 26066 7476 26078
rect 7420 26014 7422 26066
rect 7474 26014 7476 26066
rect 6748 25508 6804 25518
rect 6748 25414 6804 25452
rect 6972 25284 7028 25294
rect 6636 24670 6638 24722
rect 6690 24670 6692 24722
rect 6636 24276 6692 24670
rect 6748 24836 6804 24846
rect 6972 24836 7028 25228
rect 6748 24500 6804 24780
rect 6748 24406 6804 24444
rect 6860 24834 7028 24836
rect 6860 24782 6974 24834
rect 7026 24782 7028 24834
rect 6860 24780 7028 24782
rect 6636 24210 6692 24220
rect 6524 24110 6526 24162
rect 6578 24110 6580 24162
rect 6524 24098 6580 24110
rect 6300 23774 6302 23826
rect 6354 23774 6356 23826
rect 6300 23762 6356 23774
rect 6748 23940 6804 23950
rect 6412 23714 6468 23726
rect 6412 23662 6414 23714
rect 6466 23662 6468 23714
rect 6188 23154 6356 23156
rect 6188 23102 6190 23154
rect 6242 23102 6356 23154
rect 6188 23100 6356 23102
rect 6188 23090 6244 23100
rect 6076 22082 6132 22092
rect 6300 21700 6356 23100
rect 6412 22932 6468 23662
rect 6636 23492 6692 23502
rect 6412 22866 6468 22876
rect 6524 23436 6636 23492
rect 6412 22258 6468 22270
rect 6412 22206 6414 22258
rect 6466 22206 6468 22258
rect 6412 22148 6468 22206
rect 6412 22082 6468 22092
rect 6300 21644 6468 21700
rect 6188 21588 6244 21598
rect 6188 21494 6244 21532
rect 5964 20738 6020 20748
rect 6076 21474 6132 21486
rect 6076 21422 6078 21474
rect 6130 21422 6132 21474
rect 6076 20692 6132 21422
rect 6076 20130 6132 20636
rect 6300 21476 6356 21486
rect 6300 20690 6356 21420
rect 6300 20638 6302 20690
rect 6354 20638 6356 20690
rect 6300 20626 6356 20638
rect 6412 20244 6468 21644
rect 6524 21028 6580 23436
rect 6636 23426 6692 23436
rect 6524 20962 6580 20972
rect 6636 23156 6692 23166
rect 6636 21586 6692 23100
rect 6636 21534 6638 21586
rect 6690 21534 6692 21586
rect 6636 20692 6692 21534
rect 6076 20078 6078 20130
rect 6130 20078 6132 20130
rect 6076 20066 6132 20078
rect 6188 20188 6468 20244
rect 6524 20690 6692 20692
rect 6524 20638 6638 20690
rect 6690 20638 6692 20690
rect 6524 20636 6692 20638
rect 5964 20020 6020 20030
rect 5964 19346 6020 19964
rect 6188 19908 6244 20188
rect 5964 19294 5966 19346
rect 6018 19294 6020 19346
rect 5964 19282 6020 19294
rect 6076 19852 6244 19908
rect 6300 20018 6356 20030
rect 6300 19966 6302 20018
rect 6354 19966 6356 20018
rect 5964 18452 6020 18462
rect 5964 17778 6020 18396
rect 5964 17726 5966 17778
rect 6018 17726 6020 17778
rect 5964 17714 6020 17726
rect 5628 17054 5630 17106
rect 5682 17054 5684 17106
rect 5628 17042 5684 17054
rect 5740 17612 5908 17668
rect 5516 16882 5572 16894
rect 5516 16830 5518 16882
rect 5570 16830 5572 16882
rect 5516 16436 5572 16830
rect 5516 16370 5572 16380
rect 5404 16258 5460 16268
rect 4732 16046 4734 16098
rect 4786 16046 4788 16098
rect 4732 16034 4788 16046
rect 5180 16100 5236 16110
rect 5180 16006 5236 16044
rect 4620 15922 4676 15932
rect 4956 15876 5012 15886
rect 4956 15782 5012 15820
rect 3836 15652 3892 15662
rect 3836 15538 3892 15596
rect 3836 15486 3838 15538
rect 3890 15486 3892 15538
rect 3836 15474 3892 15486
rect 3948 15204 4004 15708
rect 3836 15092 4004 15148
rect 4172 15708 4340 15764
rect 3500 14466 3556 14476
rect 3612 14756 3668 14766
rect 3052 13918 3054 13970
rect 3106 13918 3108 13970
rect 3052 13906 3108 13918
rect 3500 14308 3556 14318
rect 2828 13122 2884 13132
rect 2940 13186 2996 13198
rect 2940 13134 2942 13186
rect 2994 13134 2996 13186
rect 2044 13076 2100 13086
rect 2044 12982 2100 13020
rect 2940 13074 2996 13134
rect 2940 13022 2942 13074
rect 2994 13022 2996 13074
rect 2940 13010 2996 13022
rect 3388 13076 3444 13086
rect 2492 12738 2548 12750
rect 2492 12686 2494 12738
rect 2546 12686 2548 12738
rect 2044 12290 2100 12302
rect 2044 12238 2046 12290
rect 2098 12238 2100 12290
rect 1708 12178 1764 12190
rect 1708 12126 1710 12178
rect 1762 12126 1764 12178
rect 1708 11508 1764 12126
rect 1708 11442 1764 11452
rect 2044 10612 2100 12238
rect 2492 12068 2548 12686
rect 3276 12404 3332 12414
rect 3388 12404 3444 13020
rect 3276 12402 3444 12404
rect 3276 12350 3278 12402
rect 3330 12350 3444 12402
rect 3276 12348 3444 12350
rect 3276 12338 3332 12348
rect 2828 12068 2884 12078
rect 2492 12012 2828 12068
rect 2828 11974 2884 12012
rect 3500 12068 3556 14252
rect 3612 13970 3668 14700
rect 3836 14642 3892 15092
rect 3836 14590 3838 14642
rect 3890 14590 3892 14642
rect 3836 14578 3892 14590
rect 4172 14644 4228 15708
rect 4284 15540 4340 15550
rect 4284 15446 4340 15484
rect 5628 15540 5684 15550
rect 5740 15540 5796 17612
rect 5852 17442 5908 17454
rect 5852 17390 5854 17442
rect 5906 17390 5908 17442
rect 5852 17332 5908 17390
rect 5852 17276 6020 17332
rect 5964 17220 6020 17276
rect 5964 17154 6020 17164
rect 5852 17108 5908 17118
rect 5852 17014 5908 17052
rect 6076 16100 6132 19852
rect 6300 19796 6356 19966
rect 6524 20020 6580 20636
rect 6636 20626 6692 20636
rect 6524 19954 6580 19964
rect 6636 20132 6692 20142
rect 6300 17780 6356 19740
rect 6412 19908 6468 19918
rect 6412 19234 6468 19852
rect 6412 19182 6414 19234
rect 6466 19182 6468 19234
rect 6412 19170 6468 19182
rect 6524 19684 6580 19694
rect 6524 18452 6580 19628
rect 6636 19234 6692 20076
rect 6748 19572 6804 23884
rect 6860 23378 6916 24780
rect 6972 24770 7028 24780
rect 7420 24836 7476 26014
rect 7532 25394 7588 25406
rect 7532 25342 7534 25394
rect 7586 25342 7588 25394
rect 7532 24946 7588 25342
rect 7532 24894 7534 24946
rect 7586 24894 7588 24946
rect 7532 24882 7588 24894
rect 7756 25284 7812 26236
rect 7980 26290 8036 26302
rect 8204 26292 8260 26302
rect 7980 26238 7982 26290
rect 8034 26238 8036 26290
rect 7420 24770 7476 24780
rect 7196 24722 7252 24734
rect 7196 24670 7198 24722
rect 7250 24670 7252 24722
rect 7196 24500 7252 24670
rect 7532 24724 7588 24734
rect 7532 24500 7588 24668
rect 7196 24444 7588 24500
rect 7644 24498 7700 24510
rect 7644 24446 7646 24498
rect 7698 24446 7700 24498
rect 7196 24276 7252 24286
rect 6972 24164 7028 24174
rect 6972 24050 7028 24108
rect 6972 23998 6974 24050
rect 7026 23998 7028 24050
rect 6972 23986 7028 23998
rect 7084 23940 7140 23950
rect 7196 23940 7252 24220
rect 7308 23940 7364 23950
rect 7196 23938 7364 23940
rect 7196 23886 7310 23938
rect 7362 23886 7364 23938
rect 7196 23884 7364 23886
rect 7084 23846 7140 23884
rect 7308 23874 7364 23884
rect 7420 23828 7476 24444
rect 7644 24164 7700 24446
rect 7756 24500 7812 25228
rect 7868 26178 7924 26190
rect 7868 26126 7870 26178
rect 7922 26126 7924 26178
rect 7868 24722 7924 26126
rect 7868 24670 7870 24722
rect 7922 24670 7924 24722
rect 7868 24658 7924 24670
rect 7980 24724 8036 26238
rect 7980 24658 8036 24668
rect 8092 26290 8260 26292
rect 8092 26238 8206 26290
rect 8258 26238 8260 26290
rect 8092 26236 8260 26238
rect 7756 24444 8036 24500
rect 7644 24098 7700 24108
rect 7756 23828 7812 23838
rect 7420 23826 7812 23828
rect 7420 23774 7758 23826
rect 7810 23774 7812 23826
rect 7420 23772 7812 23774
rect 6860 23326 6862 23378
rect 6914 23326 6916 23378
rect 6860 23314 6916 23326
rect 7420 23380 7476 23390
rect 7532 23380 7588 23772
rect 7756 23762 7812 23772
rect 7980 23826 8036 24444
rect 8092 24388 8148 26236
rect 8204 26226 8260 26236
rect 8204 24722 8260 24734
rect 8204 24670 8206 24722
rect 8258 24670 8260 24722
rect 8204 24612 8260 24670
rect 8204 24546 8260 24556
rect 8092 24332 8260 24388
rect 8092 24164 8148 24174
rect 8092 24070 8148 24108
rect 7980 23774 7982 23826
rect 8034 23774 8036 23826
rect 7980 23762 8036 23774
rect 8204 23604 8260 24332
rect 7476 23324 7588 23380
rect 7644 23548 8260 23604
rect 7420 23314 7476 23324
rect 7084 23156 7140 23166
rect 7532 23156 7588 23166
rect 6972 23154 7140 23156
rect 6972 23102 7086 23154
rect 7138 23102 7140 23154
rect 6972 23100 7140 23102
rect 6972 22372 7028 23100
rect 7084 23090 7140 23100
rect 7420 23154 7588 23156
rect 7420 23102 7534 23154
rect 7586 23102 7588 23154
rect 7420 23100 7588 23102
rect 6972 22278 7028 22316
rect 6972 20802 7028 20814
rect 6972 20750 6974 20802
rect 7026 20750 7028 20802
rect 6972 20244 7028 20750
rect 6972 20178 7028 20188
rect 7308 20578 7364 20590
rect 7308 20526 7310 20578
rect 7362 20526 7364 20578
rect 7196 20020 7252 20030
rect 7196 19926 7252 19964
rect 6748 19516 7140 19572
rect 6636 19182 6638 19234
rect 6690 19182 6692 19234
rect 6636 19124 6692 19182
rect 6972 19236 7028 19246
rect 6972 19142 7028 19180
rect 6636 19058 6692 19068
rect 6748 19012 6804 19022
rect 6748 18918 6804 18956
rect 6524 18358 6580 18396
rect 6748 18452 6804 18462
rect 6300 17724 6468 17780
rect 6300 17444 6356 17454
rect 6188 17388 6300 17444
rect 6188 16882 6244 17388
rect 6300 17350 6356 17388
rect 6412 16994 6468 17724
rect 6412 16942 6414 16994
rect 6466 16942 6468 16994
rect 6412 16930 6468 16942
rect 6748 16996 6804 18396
rect 6860 17780 6916 17790
rect 6860 17686 6916 17724
rect 6748 16930 6804 16940
rect 6972 16996 7028 17006
rect 6972 16902 7028 16940
rect 6188 16830 6190 16882
rect 6242 16830 6244 16882
rect 6188 16818 6244 16830
rect 6860 16884 6916 16894
rect 6860 16790 6916 16828
rect 6300 16324 6356 16334
rect 6076 16006 6132 16044
rect 6188 16212 6244 16222
rect 6188 15986 6244 16156
rect 6188 15934 6190 15986
rect 6242 15934 6244 15986
rect 6188 15922 6244 15934
rect 5628 15538 5796 15540
rect 5628 15486 5630 15538
rect 5682 15486 5796 15538
rect 5628 15484 5796 15486
rect 5852 15876 5908 15886
rect 5628 15474 5684 15484
rect 4508 15428 4564 15438
rect 4732 15428 4788 15438
rect 4508 15426 4732 15428
rect 4508 15374 4510 15426
rect 4562 15374 4732 15426
rect 4508 15372 4732 15374
rect 4508 15362 4564 15372
rect 4732 15148 4788 15372
rect 5292 15426 5348 15438
rect 5292 15374 5294 15426
rect 5346 15374 5348 15426
rect 4844 15316 4900 15326
rect 4844 15222 4900 15260
rect 5292 15316 5348 15374
rect 5516 15428 5572 15438
rect 5516 15334 5572 15372
rect 5292 15148 5348 15260
rect 4172 14578 4228 14588
rect 4284 15092 4340 15102
rect 4732 15092 4900 15148
rect 4284 14642 4340 15036
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4844 14756 4900 15092
rect 4284 14590 4286 14642
rect 4338 14590 4340 14642
rect 4284 14578 4340 14590
rect 4620 14700 4900 14756
rect 4956 15092 5348 15148
rect 5740 15314 5796 15326
rect 5740 15262 5742 15314
rect 5794 15262 5796 15314
rect 5740 15204 5796 15262
rect 4620 14418 4676 14700
rect 4956 14642 5012 15092
rect 4956 14590 4958 14642
rect 5010 14590 5012 14642
rect 4956 14578 5012 14590
rect 4620 14366 4622 14418
rect 4674 14366 4676 14418
rect 4620 14354 4676 14366
rect 4732 14308 4788 14318
rect 3612 13918 3614 13970
rect 3666 13918 3668 13970
rect 3612 13906 3668 13918
rect 4620 13972 4676 13982
rect 4060 13860 4116 13870
rect 3948 13634 4004 13646
rect 3948 13582 3950 13634
rect 4002 13582 4004 13634
rect 3836 12964 3892 12974
rect 3836 12850 3892 12908
rect 3836 12798 3838 12850
rect 3890 12798 3892 12850
rect 3836 12292 3892 12798
rect 3948 12740 4004 13582
rect 4060 13076 4116 13804
rect 4172 13636 4228 13646
rect 4172 13634 4340 13636
rect 4172 13582 4174 13634
rect 4226 13582 4340 13634
rect 4172 13580 4340 13582
rect 4172 13570 4228 13580
rect 4284 13188 4340 13580
rect 4620 13634 4676 13916
rect 4620 13582 4622 13634
rect 4674 13582 4676 13634
rect 4620 13570 4676 13582
rect 4732 13524 4788 14252
rect 4844 14308 4900 14318
rect 5068 14308 5124 14318
rect 4844 14306 5012 14308
rect 4844 14254 4846 14306
rect 4898 14254 5012 14306
rect 4844 14252 5012 14254
rect 4844 14242 4900 14252
rect 4844 13860 4900 13870
rect 4844 13746 4900 13804
rect 4844 13694 4846 13746
rect 4898 13694 4900 13746
rect 4844 13682 4900 13694
rect 4732 13458 4788 13468
rect 4956 13412 5012 14252
rect 5068 14214 5124 14252
rect 5404 14196 5460 14206
rect 5180 13636 5236 13646
rect 4476 13356 4740 13366
rect 4956 13356 5124 13412
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4956 13188 5012 13198
rect 4284 13186 5012 13188
rect 4284 13134 4958 13186
rect 5010 13134 5012 13186
rect 4284 13132 5012 13134
rect 4060 13010 4116 13020
rect 4060 12740 4116 12750
rect 3948 12684 4060 12740
rect 4060 12674 4116 12684
rect 4508 12402 4564 13132
rect 4956 13122 5012 13132
rect 5068 13076 5124 13356
rect 5068 13010 5124 13020
rect 4508 12350 4510 12402
rect 4562 12350 4564 12402
rect 4508 12338 4564 12350
rect 4060 12292 4116 12302
rect 3500 12002 3556 12012
rect 3612 12290 4116 12292
rect 3612 12238 4062 12290
rect 4114 12238 4116 12290
rect 3612 12236 4116 12238
rect 2492 11508 2548 11518
rect 2492 11414 2548 11452
rect 3612 11282 3668 12236
rect 4060 12226 4116 12236
rect 3724 12068 3780 12078
rect 3724 11974 3780 12012
rect 4956 12066 5012 12078
rect 4956 12014 4958 12066
rect 5010 12014 5012 12066
rect 4172 11956 4228 11966
rect 4172 11862 4228 11900
rect 4956 11844 5012 12014
rect 4476 11788 4740 11798
rect 4956 11788 5124 11844
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 3612 11230 3614 11282
rect 3666 11230 3668 11282
rect 3612 11218 3668 11230
rect 4956 11284 5012 11294
rect 4956 11190 5012 11228
rect 5068 11172 5124 11788
rect 5068 11106 5124 11116
rect 4844 10836 4900 10846
rect 5180 10836 5236 13580
rect 4844 10834 5236 10836
rect 4844 10782 4846 10834
rect 4898 10782 5182 10834
rect 5234 10782 5236 10834
rect 4844 10780 5236 10782
rect 4844 10770 4900 10780
rect 5180 10770 5236 10780
rect 2044 10546 2100 10556
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 5404 9828 5460 14140
rect 5516 14084 5572 14094
rect 5516 13748 5572 14028
rect 5516 10836 5572 13692
rect 5628 13858 5684 13870
rect 5628 13806 5630 13858
rect 5682 13806 5684 13858
rect 5628 13636 5684 13806
rect 5628 13570 5684 13580
rect 5740 12964 5796 15148
rect 5852 15148 5908 15820
rect 6076 15316 6132 15326
rect 6076 15222 6132 15260
rect 6300 15314 6356 16268
rect 6636 16212 6692 16222
rect 6524 16210 6692 16212
rect 6524 16158 6638 16210
rect 6690 16158 6692 16210
rect 6524 16156 6692 16158
rect 6300 15262 6302 15314
rect 6354 15262 6356 15314
rect 6300 15250 6356 15262
rect 6412 15316 6468 15326
rect 5852 15092 6132 15148
rect 5852 14868 5908 14878
rect 5852 14420 5908 14812
rect 5852 13972 5908 14364
rect 5964 14530 6020 14542
rect 5964 14478 5966 14530
rect 6018 14478 6020 14530
rect 5964 14196 6020 14478
rect 5964 14130 6020 14140
rect 5852 13746 5908 13916
rect 5852 13694 5854 13746
rect 5906 13694 5908 13746
rect 5852 13682 5908 13694
rect 6076 13748 6132 15092
rect 6300 14644 6356 14654
rect 6300 14550 6356 14588
rect 6188 14530 6244 14542
rect 6188 14478 6190 14530
rect 6242 14478 6244 14530
rect 6188 13972 6244 14478
rect 6412 14420 6468 15260
rect 6524 15148 6580 16156
rect 6636 16146 6692 16156
rect 7084 15426 7140 19516
rect 7308 19234 7364 20526
rect 7420 20468 7476 23100
rect 7532 23090 7588 23100
rect 7532 22258 7588 22270
rect 7532 22206 7534 22258
rect 7586 22206 7588 22258
rect 7532 21812 7588 22206
rect 7532 21746 7588 21756
rect 7644 21810 7700 23548
rect 8316 23268 8372 26460
rect 8540 26450 8596 26460
rect 8876 26850 8932 26862
rect 8876 26798 8878 26850
rect 8930 26798 8932 26850
rect 8540 26292 8596 26302
rect 8540 26198 8596 26236
rect 8764 26290 8820 26302
rect 8764 26238 8766 26290
rect 8818 26238 8820 26290
rect 8428 26180 8484 26190
rect 8428 26086 8484 26124
rect 8428 25284 8484 25294
rect 8428 24834 8484 25228
rect 8428 24782 8430 24834
rect 8482 24782 8484 24834
rect 8428 24770 8484 24782
rect 8764 24164 8820 26238
rect 8876 25060 8932 26798
rect 9436 25172 9492 28140
rect 9436 25106 9492 25116
rect 9548 27524 9604 27534
rect 8876 24994 8932 25004
rect 8988 24948 9044 24958
rect 9548 24948 9604 27468
rect 9660 27188 9716 31052
rect 9884 29652 9940 29662
rect 9772 29596 9884 29652
rect 9772 28642 9828 29596
rect 9884 29558 9940 29596
rect 9772 28590 9774 28642
rect 9826 28590 9828 28642
rect 9772 28578 9828 28590
rect 10108 29428 10164 29438
rect 9996 27748 10052 27758
rect 9884 27188 9940 27198
rect 9660 27186 9940 27188
rect 9660 27134 9886 27186
rect 9938 27134 9940 27186
rect 9660 27132 9940 27134
rect 9884 27122 9940 27132
rect 9996 26908 10052 27692
rect 9884 26852 10052 26908
rect 9660 25620 9716 25630
rect 9660 25526 9716 25564
rect 8988 24946 9604 24948
rect 8988 24894 8990 24946
rect 9042 24894 9604 24946
rect 8988 24892 9604 24894
rect 8988 24882 9044 24892
rect 9548 24722 9604 24892
rect 9548 24670 9550 24722
rect 9602 24670 9604 24722
rect 9548 24658 9604 24670
rect 9548 24500 9604 24510
rect 8764 24098 8820 24108
rect 8876 24388 8932 24398
rect 7644 21758 7646 21810
rect 7698 21758 7700 21810
rect 7644 21746 7700 21758
rect 7868 23212 8372 23268
rect 8764 23716 8820 23726
rect 8876 23716 8932 24332
rect 8764 23714 8932 23716
rect 8764 23662 8766 23714
rect 8818 23662 8932 23714
rect 8764 23660 8932 23662
rect 9212 23716 9268 23726
rect 9436 23716 9492 23726
rect 8764 23268 8820 23660
rect 9212 23622 9268 23660
rect 9324 23714 9492 23716
rect 9324 23662 9438 23714
rect 9490 23662 9492 23714
rect 9324 23660 9492 23662
rect 9324 23268 9380 23660
rect 9436 23650 9492 23660
rect 7868 21140 7924 23212
rect 8764 23202 8820 23212
rect 8876 23212 9380 23268
rect 8428 23156 8484 23166
rect 8428 23062 8484 23100
rect 8092 23044 8148 23054
rect 8092 22148 8148 22988
rect 8876 22708 8932 23212
rect 8988 23042 9044 23054
rect 8988 22990 8990 23042
rect 9042 22990 9044 23042
rect 8988 22820 9044 22990
rect 8988 22764 9492 22820
rect 8764 22652 8932 22708
rect 8652 22372 8708 22382
rect 8652 22278 8708 22316
rect 8092 22092 8484 22148
rect 8316 21698 8372 21710
rect 8316 21646 8318 21698
rect 8370 21646 8372 21698
rect 7644 21084 7924 21140
rect 7980 21362 8036 21374
rect 7980 21310 7982 21362
rect 8034 21310 8036 21362
rect 7532 20468 7588 20478
rect 7420 20412 7532 20468
rect 7532 20130 7588 20412
rect 7532 20078 7534 20130
rect 7586 20078 7588 20130
rect 7532 20066 7588 20078
rect 7308 19182 7310 19234
rect 7362 19182 7364 19234
rect 7308 17666 7364 19182
rect 7644 19124 7700 21084
rect 7756 20916 7812 20926
rect 7756 20822 7812 20860
rect 7868 20802 7924 20814
rect 7868 20750 7870 20802
rect 7922 20750 7924 20802
rect 7756 20244 7812 20254
rect 7756 20130 7812 20188
rect 7756 20078 7758 20130
rect 7810 20078 7812 20130
rect 7756 20066 7812 20078
rect 7868 20020 7924 20750
rect 7980 20356 8036 21310
rect 8092 20802 8148 20814
rect 8092 20750 8094 20802
rect 8146 20750 8148 20802
rect 8092 20692 8148 20750
rect 8092 20626 8148 20636
rect 8316 20804 8372 21646
rect 8316 20690 8372 20748
rect 8316 20638 8318 20690
rect 8370 20638 8372 20690
rect 8316 20626 8372 20638
rect 8316 20356 8372 20366
rect 7980 20300 8148 20356
rect 7924 19964 8036 20020
rect 7868 19954 7924 19964
rect 7756 19796 7812 19806
rect 7756 19236 7812 19740
rect 7756 19234 7924 19236
rect 7756 19182 7758 19234
rect 7810 19182 7924 19234
rect 7756 19180 7924 19182
rect 7756 19170 7812 19180
rect 7308 17614 7310 17666
rect 7362 17614 7364 17666
rect 7308 17602 7364 17614
rect 7420 19068 7700 19124
rect 7420 17668 7476 19068
rect 7756 18900 7812 18910
rect 7532 18844 7756 18900
rect 7532 18450 7588 18844
rect 7756 18834 7812 18844
rect 7532 18398 7534 18450
rect 7586 18398 7588 18450
rect 7532 18386 7588 18398
rect 7868 18450 7924 19180
rect 7868 18398 7870 18450
rect 7922 18398 7924 18450
rect 7868 18386 7924 18398
rect 7420 16882 7476 17612
rect 7980 17780 8036 19964
rect 8092 19236 8148 20300
rect 8092 19170 8148 19180
rect 8316 18900 8372 20300
rect 8428 20130 8484 22092
rect 8764 21698 8820 22652
rect 9100 22484 9156 22494
rect 9100 22482 9268 22484
rect 9100 22430 9102 22482
rect 9154 22430 9268 22482
rect 9100 22428 9268 22430
rect 9100 22418 9156 22428
rect 8764 21646 8766 21698
rect 8818 21646 8820 21698
rect 8764 21634 8820 21646
rect 8876 22260 8932 22270
rect 8540 20578 8596 20590
rect 8540 20526 8542 20578
rect 8594 20526 8596 20578
rect 8540 20244 8596 20526
rect 8540 20178 8596 20188
rect 8428 20078 8430 20130
rect 8482 20078 8484 20130
rect 8428 20066 8484 20078
rect 8764 20132 8820 20142
rect 8876 20132 8932 22204
rect 9100 21588 9156 21598
rect 8988 20802 9044 20814
rect 8988 20750 8990 20802
rect 9042 20750 9044 20802
rect 8988 20468 9044 20750
rect 8988 20402 9044 20412
rect 8764 20130 8932 20132
rect 8764 20078 8766 20130
rect 8818 20078 8932 20130
rect 8764 20076 8932 20078
rect 8988 20132 9044 20142
rect 8764 20066 8820 20076
rect 8988 20038 9044 20076
rect 8540 20020 8596 20030
rect 8540 20018 8708 20020
rect 8540 19966 8542 20018
rect 8594 19966 8708 20018
rect 8540 19964 8708 19966
rect 8540 19954 8596 19964
rect 8652 19908 8708 19964
rect 8652 19842 8708 19852
rect 9100 19684 9156 21532
rect 9212 20914 9268 22428
rect 9436 22260 9492 22764
rect 9548 22482 9604 24444
rect 9884 23940 9940 26852
rect 9996 26404 10052 26414
rect 9996 26310 10052 26348
rect 10108 24052 10164 29372
rect 10220 28420 10276 31724
rect 10332 28644 10388 28654
rect 10444 28644 10500 33628
rect 10556 33460 10612 33470
rect 10556 33366 10612 33404
rect 11004 33346 11060 34972
rect 11116 34916 11172 34926
rect 11340 34916 11396 35644
rect 11564 35700 11620 36428
rect 11676 36260 11732 38110
rect 11788 36596 11844 38780
rect 11900 36820 11956 41692
rect 12012 41410 12068 41916
rect 12012 41358 12014 41410
rect 12066 41358 12068 41410
rect 12012 40628 12068 41358
rect 12124 41188 12180 42478
rect 12348 41972 12404 42590
rect 12572 42308 12628 43036
rect 12796 42754 12852 42766
rect 12796 42702 12798 42754
rect 12850 42702 12852 42754
rect 12684 42642 12740 42654
rect 12684 42590 12686 42642
rect 12738 42590 12740 42642
rect 12684 42420 12740 42590
rect 12796 42644 12852 42702
rect 12796 42578 12852 42588
rect 12684 42364 12964 42420
rect 12572 42252 12740 42308
rect 12684 42084 12740 42252
rect 12684 41990 12740 42028
rect 12796 42194 12852 42206
rect 12796 42142 12798 42194
rect 12850 42142 12852 42194
rect 12572 41972 12628 41982
rect 12348 41970 12628 41972
rect 12348 41918 12574 41970
rect 12626 41918 12628 41970
rect 12348 41916 12628 41918
rect 12572 41300 12628 41916
rect 12572 41234 12628 41244
rect 12124 41122 12180 41132
rect 12460 41076 12516 41086
rect 12460 40982 12516 41020
rect 12348 40964 12404 40974
rect 12012 40562 12068 40572
rect 12124 40962 12404 40964
rect 12124 40910 12350 40962
rect 12402 40910 12404 40962
rect 12124 40908 12404 40910
rect 12124 40402 12180 40908
rect 12348 40898 12404 40908
rect 12684 40964 12740 40974
rect 12684 40870 12740 40908
rect 12124 40350 12126 40402
rect 12178 40350 12180 40402
rect 12124 40338 12180 40350
rect 12796 40402 12852 42142
rect 12908 42084 12964 42364
rect 13244 42084 13300 42094
rect 12908 42082 13300 42084
rect 12908 42030 13246 42082
rect 13298 42030 13300 42082
rect 12908 42028 13300 42030
rect 13244 41860 13300 42028
rect 12796 40350 12798 40402
rect 12850 40350 12852 40402
rect 12796 40338 12852 40350
rect 12908 41300 12964 41310
rect 12908 41074 12964 41244
rect 12908 41022 12910 41074
rect 12962 41022 12964 41074
rect 12348 39844 12404 39854
rect 12012 39842 12404 39844
rect 12012 39790 12350 39842
rect 12402 39790 12404 39842
rect 12012 39788 12404 39790
rect 12012 39058 12068 39788
rect 12348 39778 12404 39788
rect 12012 39006 12014 39058
rect 12066 39006 12068 39058
rect 12012 37266 12068 39006
rect 12460 39730 12516 39742
rect 12460 39678 12462 39730
rect 12514 39678 12516 39730
rect 12012 37214 12014 37266
rect 12066 37214 12068 37266
rect 12012 37202 12068 37214
rect 12236 37826 12292 37838
rect 12236 37774 12238 37826
rect 12290 37774 12292 37826
rect 12236 37044 12292 37774
rect 12460 37268 12516 39678
rect 12796 39508 12852 39518
rect 12684 39506 12852 39508
rect 12684 39454 12798 39506
rect 12850 39454 12852 39506
rect 12684 39452 12852 39454
rect 12684 38948 12740 39452
rect 12796 39442 12852 39452
rect 12908 39284 12964 41022
rect 13244 40964 13300 41804
rect 13244 40898 13300 40908
rect 12684 38882 12740 38892
rect 12796 39228 12964 39284
rect 13132 40292 13188 40302
rect 12796 38668 12852 39228
rect 13020 38948 13076 38958
rect 12684 38612 12852 38668
rect 12908 38946 13076 38948
rect 12908 38894 13022 38946
rect 13074 38894 13076 38946
rect 12908 38892 13076 38894
rect 12684 38610 12740 38612
rect 12684 38558 12686 38610
rect 12738 38558 12740 38610
rect 12684 38546 12740 38558
rect 12684 38162 12740 38174
rect 12684 38110 12686 38162
rect 12738 38110 12740 38162
rect 12684 37940 12740 38110
rect 12460 37202 12516 37212
rect 12572 37884 12684 37940
rect 12572 37266 12628 37884
rect 12684 37874 12740 37884
rect 12572 37214 12574 37266
rect 12626 37214 12628 37266
rect 12236 36978 12292 36988
rect 11900 36754 11956 36764
rect 11788 36540 12516 36596
rect 11788 36482 11844 36540
rect 11788 36430 11790 36482
rect 11842 36430 11844 36482
rect 11788 36418 11844 36430
rect 12012 36370 12068 36382
rect 12012 36318 12014 36370
rect 12066 36318 12068 36370
rect 11676 36204 11956 36260
rect 11564 35698 11844 35700
rect 11564 35646 11566 35698
rect 11618 35646 11844 35698
rect 11564 35644 11844 35646
rect 11564 35634 11620 35644
rect 11116 34914 11396 34916
rect 11116 34862 11118 34914
rect 11170 34862 11396 34914
rect 11116 34860 11396 34862
rect 11788 34914 11844 35644
rect 11788 34862 11790 34914
rect 11842 34862 11844 34914
rect 11116 34850 11172 34860
rect 11788 34850 11844 34862
rect 11788 34356 11844 34366
rect 11788 34262 11844 34300
rect 11900 33572 11956 36204
rect 12012 35812 12068 36318
rect 12012 35698 12068 35756
rect 12012 35646 12014 35698
rect 12066 35646 12068 35698
rect 12012 35634 12068 35646
rect 12124 36260 12180 36270
rect 12124 34242 12180 36204
rect 12348 36036 12404 36046
rect 12124 34190 12126 34242
rect 12178 34190 12180 34242
rect 12124 34178 12180 34190
rect 12236 35980 12348 36036
rect 11900 33516 12180 33572
rect 11004 33294 11006 33346
rect 11058 33294 11060 33346
rect 11004 33282 11060 33294
rect 12012 33346 12068 33358
rect 12012 33294 12014 33346
rect 12066 33294 12068 33346
rect 10780 33236 10836 33246
rect 10780 33142 10836 33180
rect 11340 33234 11396 33246
rect 11340 33182 11342 33234
rect 11394 33182 11396 33234
rect 11228 32788 11284 32798
rect 11340 32788 11396 33182
rect 11228 32786 11396 32788
rect 11228 32734 11230 32786
rect 11282 32734 11396 32786
rect 11228 32732 11396 32734
rect 11452 33122 11508 33134
rect 11452 33070 11454 33122
rect 11506 33070 11508 33122
rect 10892 32228 10948 32238
rect 10780 32172 10892 32228
rect 10668 32116 10724 32126
rect 10556 31220 10612 31230
rect 10668 31220 10724 32060
rect 10556 31218 10724 31220
rect 10556 31166 10558 31218
rect 10610 31166 10724 31218
rect 10556 31164 10724 31166
rect 10556 31154 10612 31164
rect 10668 30324 10724 31164
rect 10780 30436 10836 32172
rect 10892 32162 10948 32172
rect 11228 32116 11284 32732
rect 11228 32050 11284 32060
rect 11452 31892 11508 33070
rect 12012 32788 12068 33294
rect 11788 32732 12012 32788
rect 10892 31836 11508 31892
rect 11564 32340 11620 32350
rect 10892 30884 10948 31836
rect 11564 31778 11620 32284
rect 11564 31726 11566 31778
rect 11618 31726 11620 31778
rect 11564 31714 11620 31726
rect 11116 31668 11172 31678
rect 11116 31666 11396 31668
rect 11116 31614 11118 31666
rect 11170 31614 11396 31666
rect 11116 31612 11396 31614
rect 11116 31602 11172 31612
rect 11004 31556 11060 31566
rect 11004 31108 11060 31500
rect 11340 31332 11396 31612
rect 11788 31666 11844 32732
rect 12012 32722 12068 32732
rect 12124 31780 12180 33516
rect 12236 32228 12292 35980
rect 12348 35970 12404 35980
rect 12460 35588 12516 36540
rect 12572 35810 12628 37214
rect 12572 35758 12574 35810
rect 12626 35758 12628 35810
rect 12572 35746 12628 35758
rect 12796 36708 12852 36718
rect 12908 36708 12964 38892
rect 13020 38882 13076 38892
rect 13132 38668 13188 40236
rect 13356 40180 13412 43148
rect 13356 40114 13412 40124
rect 13356 38948 13412 38958
rect 13356 38834 13412 38892
rect 13356 38782 13358 38834
rect 13410 38782 13412 38834
rect 13356 38770 13412 38782
rect 12796 36706 12964 36708
rect 12796 36654 12798 36706
rect 12850 36654 12964 36706
rect 12796 36652 12964 36654
rect 13020 38612 13188 38668
rect 13244 38724 13300 38734
rect 12796 35810 12852 36652
rect 13020 35922 13076 38612
rect 13020 35870 13022 35922
rect 13074 35870 13076 35922
rect 13020 35858 13076 35870
rect 13132 35924 13188 35934
rect 13244 35924 13300 38668
rect 13468 38052 13524 43374
rect 13692 42644 13748 43486
rect 13692 42550 13748 42588
rect 13916 41972 13972 41982
rect 13916 41878 13972 41916
rect 14028 41748 14084 45388
rect 14140 45108 14196 45118
rect 14140 43764 14196 45052
rect 14140 43538 14196 43708
rect 14140 43486 14142 43538
rect 14194 43486 14196 43538
rect 14140 43474 14196 43486
rect 14252 42980 14308 45726
rect 14700 45220 14756 45230
rect 14700 45106 14756 45164
rect 14700 45054 14702 45106
rect 14754 45054 14756 45106
rect 14588 44212 14644 44222
rect 14476 44210 14644 44212
rect 14476 44158 14590 44210
rect 14642 44158 14644 44210
rect 14476 44156 14644 44158
rect 14476 43316 14532 44156
rect 14588 44146 14644 44156
rect 14700 43988 14756 45054
rect 14588 43932 14756 43988
rect 14588 43762 14644 43932
rect 14588 43710 14590 43762
rect 14642 43710 14644 43762
rect 14588 43698 14644 43710
rect 14812 43762 14868 45836
rect 14924 45444 14980 53452
rect 15148 53396 15204 53678
rect 15148 53330 15204 53340
rect 15260 53506 15316 53518
rect 15260 53454 15262 53506
rect 15314 53454 15316 53506
rect 15036 53060 15092 53070
rect 15036 52966 15092 53004
rect 15148 52948 15204 52958
rect 15260 52948 15316 53454
rect 15372 53172 15428 53900
rect 15484 53730 15540 53742
rect 15484 53678 15486 53730
rect 15538 53678 15540 53730
rect 15484 53620 15540 53678
rect 15596 53732 15652 56028
rect 15820 54404 15876 56924
rect 16044 56866 16100 56924
rect 16044 56814 16046 56866
rect 16098 56814 16100 56866
rect 16044 56802 16100 56814
rect 16156 56532 16212 57148
rect 16268 56756 16324 56766
rect 16380 56756 16436 57596
rect 16716 57426 16772 57438
rect 16716 57374 16718 57426
rect 16770 57374 16772 57426
rect 16492 56980 16548 56990
rect 16548 56924 16660 56980
rect 16492 56914 16548 56924
rect 16268 56754 16436 56756
rect 16268 56702 16270 56754
rect 16322 56702 16436 56754
rect 16268 56700 16436 56702
rect 16268 56690 16324 56700
rect 16156 56476 16324 56532
rect 16156 56194 16212 56206
rect 16156 56142 16158 56194
rect 16210 56142 16212 56194
rect 15932 56084 15988 56094
rect 15932 55990 15988 56028
rect 16156 55860 16212 56142
rect 15820 54338 15876 54348
rect 15932 54964 15988 54974
rect 15932 54626 15988 54908
rect 15932 54574 15934 54626
rect 15986 54574 15988 54626
rect 15932 54068 15988 54574
rect 16156 54628 16212 55804
rect 16268 55188 16324 56476
rect 16604 56194 16660 56924
rect 16604 56142 16606 56194
rect 16658 56142 16660 56194
rect 16604 56130 16660 56142
rect 16716 56084 16772 57374
rect 16828 56866 16884 56878
rect 16828 56814 16830 56866
rect 16882 56814 16884 56866
rect 16828 56532 16884 56814
rect 17052 56756 17108 59948
rect 23884 59948 24500 60004
rect 19964 59892 20020 59902
rect 19964 59798 20020 59836
rect 20860 59892 20916 59902
rect 20076 59780 20132 59790
rect 20300 59780 20356 59790
rect 20076 59778 20244 59780
rect 20076 59726 20078 59778
rect 20130 59726 20244 59778
rect 20076 59724 20244 59726
rect 20076 59714 20132 59724
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 20188 59444 20244 59724
rect 20300 59686 20356 59724
rect 20076 59388 20244 59444
rect 17948 59332 18004 59342
rect 17948 59238 18004 59276
rect 19404 58996 19460 59006
rect 19404 58994 19572 58996
rect 19404 58942 19406 58994
rect 19458 58942 19572 58994
rect 19404 58940 19572 58942
rect 19404 58930 19460 58940
rect 19516 58884 19572 58940
rect 17948 58434 18004 58446
rect 17948 58382 17950 58434
rect 18002 58382 18004 58434
rect 17164 58212 17220 58222
rect 17164 58210 17332 58212
rect 17164 58158 17166 58210
rect 17218 58158 17332 58210
rect 17164 58156 17332 58158
rect 17164 58146 17220 58156
rect 17164 57988 17220 57998
rect 17164 57090 17220 57932
rect 17164 57038 17166 57090
rect 17218 57038 17220 57090
rect 17164 57026 17220 57038
rect 17052 56690 17108 56700
rect 16828 56466 16884 56476
rect 16716 56018 16772 56028
rect 17276 55636 17332 58156
rect 17836 58210 17892 58222
rect 17836 58158 17838 58210
rect 17890 58158 17892 58210
rect 17612 57428 17668 57438
rect 17500 57426 17668 57428
rect 17500 57374 17614 57426
rect 17666 57374 17668 57426
rect 17500 57372 17668 57374
rect 17500 56082 17556 57372
rect 17612 57362 17668 57372
rect 17836 57204 17892 58158
rect 17948 57764 18004 58382
rect 17948 57698 18004 57708
rect 18508 58434 18564 58446
rect 18508 58382 18510 58434
rect 18562 58382 18564 58434
rect 18172 57538 18228 57550
rect 18172 57486 18174 57538
rect 18226 57486 18228 57538
rect 17836 57138 17892 57148
rect 17948 57426 18004 57438
rect 17948 57374 17950 57426
rect 18002 57374 18004 57426
rect 17948 56868 18004 57374
rect 18172 56980 18228 57486
rect 18508 57092 18564 58382
rect 19180 58434 19236 58446
rect 19180 58382 19182 58434
rect 19234 58382 19236 58434
rect 18844 58100 18900 58110
rect 18844 57876 18900 58044
rect 19180 57988 19236 58382
rect 19180 57922 19236 57932
rect 18844 57650 18900 57820
rect 19404 57764 19460 57774
rect 18844 57598 18846 57650
rect 18898 57598 18900 57650
rect 18844 57586 18900 57598
rect 19180 57650 19236 57662
rect 19180 57598 19182 57650
rect 19234 57598 19236 57650
rect 18508 57026 18564 57036
rect 18228 56924 18452 56980
rect 18172 56914 18228 56924
rect 17836 56812 18004 56868
rect 17500 56030 17502 56082
rect 17554 56030 17556 56082
rect 17500 56018 17556 56030
rect 17612 56754 17668 56766
rect 17612 56702 17614 56754
rect 17666 56702 17668 56754
rect 17276 55570 17332 55580
rect 16492 55188 16548 55198
rect 17612 55188 17668 56702
rect 16268 55122 16324 55132
rect 16380 55186 16548 55188
rect 16380 55134 16494 55186
rect 16546 55134 16548 55186
rect 16380 55132 16548 55134
rect 16156 54516 16212 54572
rect 15596 53666 15652 53676
rect 15708 54012 15988 54068
rect 16044 54514 16212 54516
rect 16044 54462 16158 54514
rect 16210 54462 16212 54514
rect 16044 54460 16212 54462
rect 15708 53730 15764 54012
rect 15708 53678 15710 53730
rect 15762 53678 15764 53730
rect 15708 53666 15764 53678
rect 15932 53844 15988 53854
rect 15484 53172 15540 53564
rect 15820 53506 15876 53518
rect 15820 53454 15822 53506
rect 15874 53454 15876 53506
rect 15484 53116 15764 53172
rect 15372 53106 15428 53116
rect 15596 52948 15652 52958
rect 15260 52946 15652 52948
rect 15260 52894 15598 52946
rect 15650 52894 15652 52946
rect 15260 52892 15652 52894
rect 15148 52854 15204 52892
rect 15596 52882 15652 52892
rect 15148 52724 15204 52734
rect 15148 52630 15204 52668
rect 15372 52724 15428 52734
rect 15260 52276 15316 52286
rect 15260 52182 15316 52220
rect 15036 52164 15092 52174
rect 15036 50036 15092 52108
rect 15148 52162 15204 52174
rect 15148 52110 15150 52162
rect 15202 52110 15204 52162
rect 15148 51604 15204 52110
rect 15372 51940 15428 52668
rect 15708 52274 15764 53116
rect 15820 52946 15876 53454
rect 15932 53508 15988 53788
rect 16044 53730 16100 54460
rect 16156 54450 16212 54460
rect 16268 54404 16324 54414
rect 16044 53678 16046 53730
rect 16098 53678 16100 53730
rect 16044 53666 16100 53678
rect 16156 54292 16212 54302
rect 16156 53732 16212 54236
rect 16268 53954 16324 54348
rect 16268 53902 16270 53954
rect 16322 53902 16324 53954
rect 16268 53890 16324 53902
rect 16380 53956 16436 55132
rect 16492 55122 16548 55132
rect 17276 55132 17668 55188
rect 17724 56642 17780 56654
rect 17724 56590 17726 56642
rect 17778 56590 17780 56642
rect 16716 54628 16772 54638
rect 16380 53890 16436 53900
rect 16492 54626 16772 54628
rect 16492 54574 16718 54626
rect 16770 54574 16772 54626
rect 16492 54572 16772 54574
rect 16268 53732 16324 53742
rect 16156 53676 16268 53732
rect 16268 53638 16324 53676
rect 15932 53452 16100 53508
rect 15820 52894 15822 52946
rect 15874 52894 15876 52946
rect 15820 52882 15876 52894
rect 15932 53060 15988 53070
rect 15708 52222 15710 52274
rect 15762 52222 15764 52274
rect 15708 52210 15764 52222
rect 15820 52612 15876 52622
rect 15148 51538 15204 51548
rect 15260 51884 15428 51940
rect 15820 52162 15876 52556
rect 15820 52110 15822 52162
rect 15874 52110 15876 52162
rect 15260 51380 15316 51884
rect 15820 51716 15876 52110
rect 15596 51660 15876 51716
rect 15148 51324 15316 51380
rect 15484 51380 15540 51390
rect 15148 50594 15204 51324
rect 15148 50542 15150 50594
rect 15202 50542 15204 50594
rect 15148 50530 15204 50542
rect 15260 50708 15316 50718
rect 15260 50482 15316 50652
rect 15484 50594 15540 51324
rect 15484 50542 15486 50594
rect 15538 50542 15540 50594
rect 15484 50530 15540 50542
rect 15260 50430 15262 50482
rect 15314 50430 15316 50482
rect 15260 50418 15316 50430
rect 15036 49980 15316 50036
rect 15260 49476 15316 49980
rect 15484 49924 15540 49934
rect 15484 49698 15540 49868
rect 15484 49646 15486 49698
rect 15538 49646 15540 49698
rect 15484 49634 15540 49646
rect 15260 49410 15316 49420
rect 15372 49588 15428 49598
rect 15260 48914 15316 48926
rect 15260 48862 15262 48914
rect 15314 48862 15316 48914
rect 15260 48804 15316 48862
rect 15260 48738 15316 48748
rect 15372 48242 15428 49532
rect 15484 49476 15540 49486
rect 15484 49028 15540 49420
rect 15596 49252 15652 51660
rect 15820 51268 15876 51278
rect 15820 50706 15876 51212
rect 15820 50654 15822 50706
rect 15874 50654 15876 50706
rect 15820 50642 15876 50654
rect 15932 50594 15988 53004
rect 16044 52948 16100 53452
rect 16380 52948 16436 52958
rect 16044 52946 16436 52948
rect 16044 52894 16382 52946
rect 16434 52894 16436 52946
rect 16044 52892 16436 52894
rect 16044 52724 16100 52734
rect 16044 52162 16100 52668
rect 16044 52110 16046 52162
rect 16098 52110 16100 52162
rect 16044 52098 16100 52110
rect 16268 52164 16324 52174
rect 16156 52052 16212 52062
rect 15932 50542 15934 50594
rect 15986 50542 15988 50594
rect 15932 50530 15988 50542
rect 16044 50820 16100 50830
rect 15708 50484 15764 50522
rect 15708 50418 15764 50428
rect 15708 49812 15764 49822
rect 15708 49718 15764 49756
rect 16044 49700 16100 50764
rect 16156 50482 16212 51996
rect 16268 50708 16324 52108
rect 16380 51156 16436 52892
rect 16380 51090 16436 51100
rect 16268 50642 16324 50652
rect 16156 50430 16158 50482
rect 16210 50430 16212 50482
rect 16156 50418 16212 50430
rect 16492 50428 16548 54572
rect 16716 54562 16772 54572
rect 16828 54516 16884 54526
rect 17276 54516 17332 55132
rect 17388 54964 17444 54974
rect 17388 54626 17444 54908
rect 17388 54574 17390 54626
rect 17442 54574 17444 54626
rect 17388 54562 17444 54574
rect 17612 54628 17668 54638
rect 17612 54534 17668 54572
rect 16828 54514 17332 54516
rect 16828 54462 16830 54514
rect 16882 54462 17332 54514
rect 16828 54460 17332 54462
rect 16828 54450 16884 54460
rect 16716 54290 16772 54302
rect 16716 54238 16718 54290
rect 16770 54238 16772 54290
rect 16604 53060 16660 53070
rect 16604 52612 16660 53004
rect 16604 52546 16660 52556
rect 16716 51716 16772 54238
rect 16828 53620 16884 53630
rect 16828 53526 16884 53564
rect 16940 53508 16996 53518
rect 16940 53414 16996 53452
rect 17052 53284 17108 54460
rect 17500 54402 17556 54414
rect 17500 54350 17502 54402
rect 17554 54350 17556 54402
rect 17500 54068 17556 54350
rect 17500 54002 17556 54012
rect 17612 53844 17668 53854
rect 17276 53732 17332 53742
rect 17276 53638 17332 53676
rect 17164 53620 17220 53630
rect 17164 53526 17220 53564
rect 17052 53218 17108 53228
rect 17500 52948 17556 52958
rect 17500 52836 17556 52892
rect 17388 52834 17556 52836
rect 17388 52782 17502 52834
rect 17554 52782 17556 52834
rect 17388 52780 17556 52782
rect 17388 52164 17444 52780
rect 17500 52770 17556 52780
rect 17612 52612 17668 53788
rect 17388 52098 17444 52108
rect 17500 52556 17668 52612
rect 17276 52050 17332 52062
rect 17276 51998 17278 52050
rect 17330 51998 17332 52050
rect 16940 51940 16996 51950
rect 16940 51938 17220 51940
rect 16940 51886 16942 51938
rect 16994 51886 17220 51938
rect 16940 51884 17220 51886
rect 16940 51874 16996 51884
rect 17164 51716 17220 51884
rect 16716 51660 17108 51716
rect 16828 51492 16884 51502
rect 16828 51266 16884 51436
rect 16828 51214 16830 51266
rect 16882 51214 16884 51266
rect 16828 51202 16884 51214
rect 16044 49634 16100 49644
rect 16268 50372 16548 50428
rect 16604 50372 16660 50382
rect 16044 49476 16100 49486
rect 15596 49196 15764 49252
rect 15596 49028 15652 49038
rect 15484 49026 15652 49028
rect 15484 48974 15598 49026
rect 15650 48974 15652 49026
rect 15484 48972 15652 48974
rect 15596 48962 15652 48972
rect 15372 48190 15374 48242
rect 15426 48190 15428 48242
rect 15372 48178 15428 48190
rect 15484 47908 15540 47918
rect 15484 47458 15540 47852
rect 15484 47406 15486 47458
rect 15538 47406 15540 47458
rect 15484 47394 15540 47406
rect 15372 47348 15428 47358
rect 15372 47254 15428 47292
rect 15484 47124 15540 47134
rect 15372 46900 15428 46910
rect 15372 46786 15428 46844
rect 15372 46734 15374 46786
rect 15426 46734 15428 46786
rect 14924 45378 14980 45388
rect 15036 46564 15092 46574
rect 14812 43710 14814 43762
rect 14866 43710 14868 43762
rect 14812 43698 14868 43710
rect 15036 44772 15092 46508
rect 15372 46452 15428 46734
rect 15372 46386 15428 46396
rect 15148 45892 15204 45902
rect 15148 45798 15204 45836
rect 15372 45108 15428 45146
rect 15372 45042 15428 45052
rect 15484 44996 15540 47068
rect 15484 44930 15540 44940
rect 15596 45108 15652 45118
rect 14700 43652 14756 43662
rect 14700 43558 14756 43596
rect 14476 43260 14756 43316
rect 14140 42924 14308 42980
rect 14700 42978 14756 43260
rect 14700 42926 14702 42978
rect 14754 42926 14756 42978
rect 14140 42196 14196 42924
rect 14700 42914 14756 42926
rect 15036 42868 15092 44716
rect 15372 43650 15428 43662
rect 15372 43598 15374 43650
rect 15426 43598 15428 43650
rect 15260 43538 15316 43550
rect 15260 43486 15262 43538
rect 15314 43486 15316 43538
rect 15148 42980 15204 42990
rect 15260 42980 15316 43486
rect 15204 42924 15316 42980
rect 15372 42980 15428 43598
rect 15596 43650 15652 45052
rect 15596 43598 15598 43650
rect 15650 43598 15652 43650
rect 15596 43586 15652 43598
rect 15148 42914 15204 42924
rect 15372 42914 15428 42924
rect 14812 42812 15092 42868
rect 14252 42756 14308 42766
rect 14252 42662 14308 42700
rect 14588 42754 14644 42766
rect 14588 42702 14590 42754
rect 14642 42702 14644 42754
rect 14588 42532 14644 42702
rect 14812 42754 14868 42812
rect 14812 42702 14814 42754
rect 14866 42702 14868 42754
rect 14812 42690 14868 42702
rect 15148 42754 15204 42766
rect 15148 42702 15150 42754
rect 15202 42702 15204 42754
rect 14588 42476 14756 42532
rect 14140 42140 14308 42196
rect 14140 41970 14196 41982
rect 14140 41918 14142 41970
rect 14194 41918 14196 41970
rect 14140 41860 14196 41918
rect 14140 41794 14196 41804
rect 13916 41692 14084 41748
rect 13804 41074 13860 41086
rect 13804 41022 13806 41074
rect 13858 41022 13860 41074
rect 13580 40964 13636 40974
rect 13580 38274 13636 40908
rect 13692 39956 13748 39966
rect 13692 39730 13748 39900
rect 13692 39678 13694 39730
rect 13746 39678 13748 39730
rect 13692 38668 13748 39678
rect 13804 39620 13860 41022
rect 13804 39554 13860 39564
rect 13692 38612 13860 38668
rect 13580 38222 13582 38274
rect 13634 38222 13636 38274
rect 13580 38210 13636 38222
rect 13468 37986 13524 37996
rect 13692 38050 13748 38062
rect 13692 37998 13694 38050
rect 13746 37998 13748 38050
rect 13692 37940 13748 37998
rect 13692 37874 13748 37884
rect 13132 35922 13300 35924
rect 13132 35870 13134 35922
rect 13186 35870 13300 35922
rect 13132 35868 13300 35870
rect 13356 37604 13412 37614
rect 13356 37380 13412 37548
rect 13804 37380 13860 38612
rect 13916 37604 13972 41692
rect 14140 41076 14196 41086
rect 14028 40962 14084 40974
rect 14028 40910 14030 40962
rect 14082 40910 14084 40962
rect 14028 39844 14084 40910
rect 14028 39778 14084 39788
rect 14028 39620 14084 39630
rect 14028 39526 14084 39564
rect 14140 39506 14196 41020
rect 14252 40404 14308 42140
rect 14700 42194 14756 42476
rect 14700 42142 14702 42194
rect 14754 42142 14756 42194
rect 14700 42130 14756 42142
rect 14924 42082 14980 42094
rect 14924 42030 14926 42082
rect 14978 42030 14980 42082
rect 14476 41970 14532 41982
rect 14476 41918 14478 41970
rect 14530 41918 14532 41970
rect 14364 41858 14420 41870
rect 14364 41806 14366 41858
rect 14418 41806 14420 41858
rect 14364 41074 14420 41806
rect 14476 41300 14532 41918
rect 14924 41300 14980 42030
rect 15036 42084 15092 42094
rect 15036 41990 15092 42028
rect 15148 41972 15204 42702
rect 15372 42754 15428 42766
rect 15372 42702 15374 42754
rect 15426 42702 15428 42754
rect 15148 41906 15204 41916
rect 15260 42644 15316 42654
rect 15260 41972 15316 42588
rect 15372 42196 15428 42702
rect 15484 42196 15540 42206
rect 15372 42194 15540 42196
rect 15372 42142 15486 42194
rect 15538 42142 15540 42194
rect 15372 42140 15540 42142
rect 15484 42130 15540 42140
rect 15372 41972 15428 41982
rect 15260 41970 15428 41972
rect 15260 41918 15374 41970
rect 15426 41918 15428 41970
rect 15260 41916 15428 41918
rect 15260 41636 15316 41916
rect 15372 41906 15428 41916
rect 15596 41970 15652 41982
rect 15596 41918 15598 41970
rect 15650 41918 15652 41970
rect 15260 41580 15540 41636
rect 15260 41412 15316 41422
rect 14924 41244 15204 41300
rect 14476 41234 14532 41244
rect 14364 41022 14366 41074
rect 14418 41022 14420 41074
rect 14364 40964 14420 41022
rect 14924 41074 14980 41086
rect 14924 41022 14926 41074
rect 14978 41022 14980 41074
rect 14364 40908 14868 40964
rect 14588 40404 14644 40442
rect 14252 40348 14532 40404
rect 14140 39454 14142 39506
rect 14194 39454 14196 39506
rect 14140 39442 14196 39454
rect 14252 40180 14308 40190
rect 14252 38668 14308 40124
rect 14476 39620 14532 40348
rect 14588 40338 14644 40348
rect 14700 40290 14756 40302
rect 14700 40238 14702 40290
rect 14754 40238 14756 40290
rect 14476 39554 14532 39564
rect 14588 40178 14644 40190
rect 14588 40126 14590 40178
rect 14642 40126 14644 40178
rect 14364 38836 14420 38846
rect 14364 38742 14420 38780
rect 14252 38612 14532 38668
rect 13916 37538 13972 37548
rect 14364 37938 14420 37950
rect 14364 37886 14366 37938
rect 14418 37886 14420 37938
rect 13132 35858 13188 35868
rect 12796 35758 12798 35810
rect 12850 35758 12852 35810
rect 12796 35746 12852 35758
rect 12908 35810 12964 35822
rect 12908 35758 12910 35810
rect 12962 35758 12964 35810
rect 12460 35532 12628 35588
rect 12572 35476 12628 35532
rect 12908 35476 12964 35758
rect 13356 35700 13412 37324
rect 13692 37324 13860 37380
rect 12572 35420 12964 35476
rect 13020 35644 13412 35700
rect 13580 36484 13636 36494
rect 13692 36484 13748 37324
rect 13916 37268 13972 37278
rect 14252 37268 14308 37278
rect 13972 37266 14308 37268
rect 13972 37214 14254 37266
rect 14306 37214 14308 37266
rect 13972 37212 14308 37214
rect 13916 37156 13972 37212
rect 14252 37202 14308 37212
rect 14364 37268 14420 37886
rect 14476 37378 14532 38612
rect 14588 38276 14644 40126
rect 14700 40180 14756 40238
rect 14700 40114 14756 40124
rect 14812 39730 14868 40908
rect 14924 40628 14980 41022
rect 15036 41076 15092 41086
rect 15036 40982 15092 41020
rect 15148 40852 15204 41244
rect 15260 41186 15316 41356
rect 15260 41134 15262 41186
rect 15314 41134 15316 41186
rect 15260 41122 15316 41134
rect 15372 41300 15428 41310
rect 14924 40562 14980 40572
rect 15036 40796 15204 40852
rect 15036 40180 15092 40796
rect 14812 39678 14814 39730
rect 14866 39678 14868 39730
rect 14812 39666 14868 39678
rect 14924 40124 15092 40180
rect 14812 39508 14868 39518
rect 14812 39414 14868 39452
rect 14700 39396 14756 39406
rect 14700 38724 14756 39340
rect 14700 38658 14756 38668
rect 14588 38220 14868 38276
rect 14476 37326 14478 37378
rect 14530 37326 14532 37378
rect 14476 37314 14532 37326
rect 14588 38052 14644 38062
rect 13636 36428 13748 36484
rect 13804 37100 13972 37156
rect 13580 36258 13636 36428
rect 13580 36206 13582 36258
rect 13634 36206 13636 36258
rect 12796 34802 12852 34814
rect 12796 34750 12798 34802
rect 12850 34750 12852 34802
rect 12684 34690 12740 34702
rect 12684 34638 12686 34690
rect 12738 34638 12740 34690
rect 12684 33684 12740 34638
rect 12796 34356 12852 34750
rect 12908 34356 12964 34366
rect 12796 34354 12964 34356
rect 12796 34302 12910 34354
rect 12962 34302 12964 34354
rect 12796 34300 12964 34302
rect 12908 34290 12964 34300
rect 12684 33618 12740 33628
rect 12796 33460 12852 33470
rect 12796 33366 12852 33404
rect 12236 32162 12292 32172
rect 12348 33348 12404 33358
rect 11788 31614 11790 31666
rect 11842 31614 11844 31666
rect 11788 31602 11844 31614
rect 11900 31724 12180 31780
rect 12236 31892 12292 31902
rect 11900 31444 11956 31724
rect 11788 31388 11956 31444
rect 12124 31554 12180 31566
rect 12124 31502 12126 31554
rect 12178 31502 12180 31554
rect 11340 31276 11732 31332
rect 11676 31220 11732 31276
rect 11676 31126 11732 31164
rect 11004 31052 11396 31108
rect 10892 30818 10948 30828
rect 11228 30884 11284 30894
rect 10780 30380 11172 30436
rect 10668 30322 10836 30324
rect 10668 30270 10670 30322
rect 10722 30270 10836 30322
rect 10668 30268 10836 30270
rect 10668 30258 10724 30268
rect 10780 29538 10836 30268
rect 10780 29486 10782 29538
rect 10834 29486 10836 29538
rect 10780 29474 10836 29486
rect 10556 28756 10612 28766
rect 10556 28662 10612 28700
rect 10388 28588 10500 28644
rect 10332 28578 10388 28588
rect 10220 28364 10388 28420
rect 10220 27412 10276 27422
rect 10220 27188 10276 27356
rect 10220 27094 10276 27132
rect 10332 26908 10388 28364
rect 10556 28084 10612 28094
rect 10556 27990 10612 28028
rect 10892 27972 10948 27982
rect 10892 27074 10948 27916
rect 10892 27022 10894 27074
rect 10946 27022 10948 27074
rect 10892 27010 10948 27022
rect 11004 27076 11060 27086
rect 11116 27076 11172 30380
rect 11228 30210 11284 30828
rect 11228 30158 11230 30210
rect 11282 30158 11284 30210
rect 11228 30146 11284 30158
rect 11340 30098 11396 31052
rect 11564 30212 11620 30222
rect 11564 30118 11620 30156
rect 11340 30046 11342 30098
rect 11394 30046 11396 30098
rect 11340 30034 11396 30046
rect 11340 28530 11396 28542
rect 11340 28478 11342 28530
rect 11394 28478 11396 28530
rect 11340 28084 11396 28478
rect 11340 28018 11396 28028
rect 11564 28084 11620 28094
rect 11340 27860 11396 27870
rect 11340 27298 11396 27804
rect 11340 27246 11342 27298
rect 11394 27246 11396 27298
rect 11340 27234 11396 27246
rect 11564 27300 11620 28028
rect 11676 27972 11732 27982
rect 11676 27878 11732 27916
rect 11676 27300 11732 27310
rect 11564 27298 11732 27300
rect 11564 27246 11678 27298
rect 11730 27246 11732 27298
rect 11564 27244 11732 27246
rect 11116 27020 11396 27076
rect 10108 23986 10164 23996
rect 10220 26852 10388 26908
rect 10444 26964 10500 26974
rect 9884 23884 10052 23940
rect 9772 23828 9828 23838
rect 9772 23826 9940 23828
rect 9772 23774 9774 23826
rect 9826 23774 9940 23826
rect 9772 23772 9940 23774
rect 9772 23762 9828 23772
rect 9548 22430 9550 22482
rect 9602 22430 9604 22482
rect 9548 22418 9604 22430
rect 9660 23714 9716 23726
rect 9660 23662 9662 23714
rect 9714 23662 9716 23714
rect 9548 22260 9604 22270
rect 9436 22258 9604 22260
rect 9436 22206 9550 22258
rect 9602 22206 9604 22258
rect 9436 22204 9604 22206
rect 9212 20862 9214 20914
rect 9266 20862 9268 20914
rect 9212 20850 9268 20862
rect 9324 21812 9380 21822
rect 8316 18834 8372 18844
rect 8428 19628 9156 19684
rect 8428 18674 8484 19628
rect 8428 18622 8430 18674
rect 8482 18622 8484 18674
rect 8204 18450 8260 18462
rect 8204 18398 8206 18450
rect 8258 18398 8260 18450
rect 8204 18228 8260 18398
rect 8316 18340 8372 18350
rect 8316 18246 8372 18284
rect 8204 18162 8260 18172
rect 7980 17666 8036 17724
rect 7980 17614 7982 17666
rect 8034 17614 8036 17666
rect 7980 17602 8036 17614
rect 8316 17220 8372 17230
rect 7420 16830 7422 16882
rect 7474 16830 7476 16882
rect 7420 16818 7476 16830
rect 7980 16994 8036 17006
rect 7980 16942 7982 16994
rect 8034 16942 8036 16994
rect 7196 16770 7252 16782
rect 7196 16718 7198 16770
rect 7250 16718 7252 16770
rect 7196 15764 7252 16718
rect 7420 16098 7476 16110
rect 7420 16046 7422 16098
rect 7474 16046 7476 16098
rect 7420 15988 7476 16046
rect 7980 16100 8036 16942
rect 8316 16994 8372 17164
rect 8316 16942 8318 16994
rect 8370 16942 8372 16994
rect 8316 16930 8372 16942
rect 8428 16996 8484 18622
rect 8652 19460 8708 19470
rect 8652 18564 8708 19404
rect 7980 16034 8036 16044
rect 7420 15922 7476 15932
rect 7196 15708 7700 15764
rect 7084 15374 7086 15426
rect 7138 15374 7140 15426
rect 7084 15362 7140 15374
rect 7308 15428 7364 15438
rect 7308 15314 7364 15372
rect 7308 15262 7310 15314
rect 7362 15262 7364 15314
rect 7084 15204 7140 15242
rect 6524 15092 6916 15148
rect 7084 15138 7140 15148
rect 6860 14532 6916 15092
rect 7084 14532 7140 14542
rect 6860 14438 6916 14476
rect 6972 14530 7140 14532
rect 6972 14478 7086 14530
rect 7138 14478 7140 14530
rect 6972 14476 7140 14478
rect 6300 14364 6468 14420
rect 6300 14306 6356 14364
rect 6300 14254 6302 14306
rect 6354 14254 6356 14306
rect 6300 14242 6356 14254
rect 6188 13906 6244 13916
rect 6300 13748 6356 13758
rect 6076 13746 6356 13748
rect 6076 13694 6302 13746
rect 6354 13694 6356 13746
rect 6076 13692 6356 13694
rect 6300 13682 6356 13692
rect 6636 13522 6692 13534
rect 6636 13470 6638 13522
rect 6690 13470 6692 13522
rect 6300 13412 6356 13422
rect 6356 13356 6468 13412
rect 6300 13346 6356 13356
rect 5964 12964 6020 12974
rect 6188 12964 6244 12974
rect 5740 12908 5908 12964
rect 5628 12850 5684 12862
rect 5628 12798 5630 12850
rect 5682 12798 5684 12850
rect 5628 11956 5684 12798
rect 5740 12740 5796 12750
rect 5740 12646 5796 12684
rect 5852 12180 5908 12908
rect 5964 12962 6244 12964
rect 5964 12910 5966 12962
rect 6018 12910 6190 12962
rect 6242 12910 6244 12962
rect 5964 12908 6244 12910
rect 5964 12898 6020 12908
rect 6188 12898 6244 12908
rect 5964 12180 6020 12190
rect 5852 12124 5964 12180
rect 5964 12066 6020 12124
rect 6076 12180 6132 12190
rect 6076 12178 6356 12180
rect 6076 12126 6078 12178
rect 6130 12126 6356 12178
rect 6076 12124 6356 12126
rect 6076 12114 6132 12124
rect 5964 12014 5966 12066
rect 6018 12014 6020 12066
rect 5964 12002 6020 12014
rect 5628 11620 5684 11900
rect 5628 11564 6020 11620
rect 5740 11394 5796 11406
rect 5740 11342 5742 11394
rect 5794 11342 5796 11394
rect 5740 11284 5796 11342
rect 5740 11218 5796 11228
rect 5852 11282 5908 11294
rect 5852 11230 5854 11282
rect 5906 11230 5908 11282
rect 5628 10836 5684 10846
rect 5516 10834 5684 10836
rect 5516 10782 5630 10834
rect 5682 10782 5684 10834
rect 5516 10780 5684 10782
rect 5628 10050 5684 10780
rect 5852 10724 5908 11230
rect 5852 10658 5908 10668
rect 5964 10948 6020 11564
rect 5964 10722 6020 10892
rect 6076 11172 6132 11182
rect 6076 10834 6132 11116
rect 6076 10782 6078 10834
rect 6130 10782 6132 10834
rect 6076 10770 6132 10782
rect 6300 10834 6356 12124
rect 6300 10782 6302 10834
rect 6354 10782 6356 10834
rect 6300 10770 6356 10782
rect 6412 10836 6468 13356
rect 6524 12850 6580 12862
rect 6524 12798 6526 12850
rect 6578 12798 6580 12850
rect 6524 12068 6580 12798
rect 6636 12852 6692 13470
rect 6860 13300 6916 13310
rect 6636 12786 6692 12796
rect 6748 13244 6860 13300
rect 6524 12002 6580 12012
rect 6524 11396 6580 11406
rect 6748 11396 6804 13244
rect 6860 13234 6916 13244
rect 6972 12740 7028 14476
rect 7084 14466 7140 14476
rect 7196 13972 7252 13982
rect 7196 13878 7252 13916
rect 7308 13858 7364 15262
rect 7644 15148 7700 15708
rect 8428 15314 8484 16940
rect 8428 15262 8430 15314
rect 8482 15262 8484 15314
rect 8428 15250 8484 15262
rect 8540 18562 8708 18564
rect 8540 18510 8654 18562
rect 8706 18510 8708 18562
rect 8540 18508 8708 18510
rect 8540 16770 8596 18508
rect 8652 18498 8708 18508
rect 9324 18340 9380 21756
rect 9548 20804 9604 22204
rect 9660 22260 9716 23662
rect 9772 23380 9828 23390
rect 9772 23286 9828 23324
rect 9772 23044 9828 23054
rect 9884 23044 9940 23772
rect 9828 22988 9940 23044
rect 9772 22978 9828 22988
rect 9660 22194 9716 22204
rect 9772 22370 9828 22382
rect 9772 22318 9774 22370
rect 9826 22318 9828 22370
rect 9548 20710 9604 20748
rect 9436 20692 9492 20702
rect 9436 20598 9492 20636
rect 9772 20356 9828 22318
rect 9884 21476 9940 21486
rect 9884 21382 9940 21420
rect 9436 20300 9828 20356
rect 9436 19236 9492 20300
rect 9996 20244 10052 23884
rect 10220 23716 10276 26852
rect 10332 25844 10388 25854
rect 10332 25618 10388 25788
rect 10332 25566 10334 25618
rect 10386 25566 10388 25618
rect 10332 25554 10388 25566
rect 10332 24612 10388 24622
rect 10332 24518 10388 24556
rect 10332 23716 10388 23726
rect 10220 23714 10388 23716
rect 10220 23662 10334 23714
rect 10386 23662 10388 23714
rect 10220 23660 10388 23662
rect 10220 23492 10276 23502
rect 9884 20188 10052 20244
rect 10108 23154 10164 23166
rect 10108 23102 10110 23154
rect 10162 23102 10164 23154
rect 10108 20692 10164 23102
rect 10220 22370 10276 23436
rect 10220 22318 10222 22370
rect 10274 22318 10276 22370
rect 10220 22306 10276 22318
rect 9436 19170 9492 19180
rect 9548 20018 9604 20030
rect 9548 19966 9550 20018
rect 9602 19966 9604 20018
rect 8540 16718 8542 16770
rect 8594 16718 8596 16770
rect 8540 15148 8596 16718
rect 8652 18284 9380 18340
rect 8652 15764 8708 18284
rect 9548 18228 9604 19966
rect 9772 20020 9828 20030
rect 9772 19926 9828 19964
rect 9884 19572 9940 20188
rect 9884 19506 9940 19516
rect 9996 20020 10052 20030
rect 9548 18162 9604 18172
rect 9660 19234 9716 19246
rect 9660 19182 9662 19234
rect 9714 19182 9716 19234
rect 9660 17668 9716 19182
rect 9884 19236 9940 19246
rect 9996 19236 10052 19964
rect 10108 19906 10164 20636
rect 10108 19854 10110 19906
rect 10162 19854 10164 19906
rect 10108 19842 10164 19854
rect 10220 21362 10276 21374
rect 10220 21310 10222 21362
rect 10274 21310 10276 21362
rect 9940 19180 10052 19236
rect 10220 19236 10276 21310
rect 10332 21028 10388 23660
rect 10444 22484 10500 26908
rect 10668 26964 10724 26974
rect 11004 26964 11060 27020
rect 11004 26908 11284 26964
rect 10556 26852 10612 26862
rect 10668 26852 10724 26908
rect 10556 26850 10724 26852
rect 10556 26798 10558 26850
rect 10610 26798 10724 26850
rect 10556 26796 10724 26798
rect 10556 26786 10612 26796
rect 10668 25618 10724 26796
rect 10668 25566 10670 25618
rect 10722 25566 10724 25618
rect 10668 25554 10724 25566
rect 10780 25396 10836 25406
rect 10780 25302 10836 25340
rect 11228 25394 11284 26908
rect 11228 25342 11230 25394
rect 11282 25342 11284 25394
rect 11228 25330 11284 25342
rect 11340 25394 11396 27020
rect 11340 25342 11342 25394
rect 11394 25342 11396 25394
rect 11004 25284 11060 25294
rect 11004 25190 11060 25228
rect 10892 24276 10948 24286
rect 10892 24050 10948 24220
rect 11340 24164 11396 25342
rect 10892 23998 10894 24050
rect 10946 23998 10948 24050
rect 10892 23986 10948 23998
rect 11116 24108 11396 24164
rect 11452 26852 11508 26862
rect 11116 23826 11172 24108
rect 11452 24052 11508 26796
rect 11676 25394 11732 27244
rect 11788 26852 11844 31388
rect 12124 31220 12180 31502
rect 12124 31154 12180 31164
rect 12124 30100 12180 30110
rect 12236 30100 12292 31836
rect 12348 30772 12404 33292
rect 12684 33234 12740 33246
rect 12684 33182 12686 33234
rect 12738 33182 12740 33234
rect 12572 32452 12628 32462
rect 12572 32358 12628 32396
rect 12684 31892 12740 33182
rect 13020 32004 13076 35644
rect 13580 35364 13636 36206
rect 13132 35308 13636 35364
rect 13132 33572 13188 35308
rect 13580 35140 13636 35150
rect 13804 35140 13860 37100
rect 14028 37044 14084 37054
rect 13916 36594 13972 36606
rect 13916 36542 13918 36594
rect 13970 36542 13972 36594
rect 13916 36260 13972 36542
rect 13916 36194 13972 36204
rect 13580 35138 13860 35140
rect 13580 35086 13582 35138
rect 13634 35086 13860 35138
rect 13580 35084 13860 35086
rect 13916 35140 13972 35150
rect 14028 35140 14084 36988
rect 14140 36596 14196 36606
rect 14196 36540 14308 36596
rect 14140 36530 14196 36540
rect 13916 35138 14084 35140
rect 13916 35086 13918 35138
rect 13970 35086 14084 35138
rect 13916 35084 14084 35086
rect 14140 35810 14196 35822
rect 14140 35758 14142 35810
rect 14194 35758 14196 35810
rect 13580 35074 13636 35084
rect 13916 35074 13972 35084
rect 13804 34692 13860 34702
rect 13580 34636 13804 34692
rect 13468 34244 13524 34254
rect 13356 34242 13524 34244
rect 13356 34190 13470 34242
rect 13522 34190 13524 34242
rect 13356 34188 13524 34190
rect 13132 33506 13188 33516
rect 13244 33908 13300 33918
rect 13132 32450 13188 32462
rect 13132 32398 13134 32450
rect 13186 32398 13188 32450
rect 13132 32340 13188 32398
rect 13132 32274 13188 32284
rect 13020 31938 13076 31948
rect 12684 31826 12740 31836
rect 12684 31666 12740 31678
rect 12684 31614 12686 31666
rect 12738 31614 12740 31666
rect 12684 31444 12740 31614
rect 12572 31220 12628 31230
rect 12684 31220 12740 31388
rect 12572 31218 12740 31220
rect 12572 31166 12574 31218
rect 12626 31166 12740 31218
rect 12572 31164 12740 31166
rect 12796 31220 12852 31230
rect 12572 31154 12628 31164
rect 12796 31126 12852 31164
rect 13244 31108 13300 33852
rect 13356 32562 13412 34188
rect 13468 34178 13524 34188
rect 13356 32510 13358 32562
rect 13410 32510 13412 32562
rect 13356 32452 13412 32510
rect 13356 32386 13412 32396
rect 13468 31778 13524 31790
rect 13468 31726 13470 31778
rect 13522 31726 13524 31778
rect 13468 31220 13524 31726
rect 13468 31154 13524 31164
rect 13356 31108 13412 31118
rect 13244 31106 13412 31108
rect 13244 31054 13358 31106
rect 13410 31054 13412 31106
rect 13244 31052 13412 31054
rect 13356 31042 13412 31052
rect 12460 30996 12516 31006
rect 12460 30902 12516 30940
rect 12908 30994 12964 31006
rect 12908 30942 12910 30994
rect 12962 30942 12964 30994
rect 12348 30716 12628 30772
rect 12572 30212 12628 30716
rect 12796 30212 12852 30222
rect 12572 30210 12852 30212
rect 12572 30158 12798 30210
rect 12850 30158 12852 30210
rect 12572 30156 12852 30158
rect 12796 30146 12852 30156
rect 12908 30212 12964 30942
rect 12908 30146 12964 30156
rect 13132 30996 13188 31006
rect 12124 30098 12292 30100
rect 12124 30046 12126 30098
rect 12178 30046 12292 30098
rect 12124 30044 12292 30046
rect 12348 30098 12404 30110
rect 12348 30046 12350 30098
rect 12402 30046 12404 30098
rect 12124 30034 12180 30044
rect 12348 29650 12404 30046
rect 12348 29598 12350 29650
rect 12402 29598 12404 29650
rect 12236 27972 12292 27982
rect 12236 27858 12292 27916
rect 12236 27806 12238 27858
rect 12290 27806 12292 27858
rect 12236 27794 12292 27806
rect 12348 27860 12404 29598
rect 13020 30098 13076 30110
rect 13020 30046 13022 30098
rect 13074 30046 13076 30098
rect 13020 29092 13076 30046
rect 13020 29026 13076 29036
rect 13132 28756 13188 30940
rect 13356 29316 13412 29326
rect 13132 28690 13188 28700
rect 13244 29314 13412 29316
rect 13244 29262 13358 29314
rect 13410 29262 13412 29314
rect 13244 29260 13412 29262
rect 12796 28644 12852 28654
rect 12796 28550 12852 28588
rect 12460 28084 12516 28094
rect 12460 27970 12516 28028
rect 12460 27918 12462 27970
rect 12514 27918 12516 27970
rect 12460 27906 12516 27918
rect 12348 27794 12404 27804
rect 13020 27636 13076 27646
rect 12460 27634 13076 27636
rect 12460 27582 13022 27634
rect 13074 27582 13076 27634
rect 12460 27580 13076 27582
rect 11900 26964 11956 26974
rect 11900 26870 11956 26908
rect 12460 26962 12516 27580
rect 13020 27570 13076 27580
rect 12460 26910 12462 26962
rect 12514 26910 12516 26962
rect 11788 26786 11844 26796
rect 11788 26628 11844 26638
rect 11788 26514 11844 26572
rect 12460 26628 12516 26910
rect 12460 26562 12516 26572
rect 12572 26852 12628 26862
rect 11788 26462 11790 26514
rect 11842 26462 11844 26514
rect 11788 26450 11844 26462
rect 12236 26516 12292 26526
rect 12236 26422 12292 26460
rect 12572 26290 12628 26796
rect 13244 26852 13300 29260
rect 13356 29250 13412 29260
rect 13468 28644 13524 28654
rect 13356 27972 13412 27982
rect 13356 27878 13412 27916
rect 13244 26786 13300 26796
rect 12908 26740 12964 26750
rect 12572 26238 12574 26290
rect 12626 26238 12628 26290
rect 12572 26226 12628 26238
rect 12684 26292 12740 26302
rect 12012 25732 12068 25742
rect 12012 25508 12068 25676
rect 12572 25508 12628 25518
rect 12012 25506 12292 25508
rect 12012 25454 12014 25506
rect 12066 25454 12292 25506
rect 12012 25452 12292 25454
rect 12012 25442 12068 25452
rect 11676 25342 11678 25394
rect 11730 25342 11732 25394
rect 11676 25330 11732 25342
rect 12012 25284 12068 25294
rect 11788 24612 11844 24622
rect 11788 24162 11844 24556
rect 11788 24110 11790 24162
rect 11842 24110 11844 24162
rect 11788 24098 11844 24110
rect 11900 24500 11956 24510
rect 11116 23774 11118 23826
rect 11170 23774 11172 23826
rect 10556 23044 10612 23054
rect 11004 23044 11060 23054
rect 10556 23042 10948 23044
rect 10556 22990 10558 23042
rect 10610 22990 10948 23042
rect 10556 22988 10948 22990
rect 10556 22978 10612 22988
rect 10780 22596 10836 22606
rect 10668 22484 10724 22494
rect 10444 22482 10724 22484
rect 10444 22430 10670 22482
rect 10722 22430 10724 22482
rect 10444 22428 10724 22430
rect 10668 22418 10724 22428
rect 10780 21700 10836 22540
rect 10892 22260 10948 22988
rect 10892 22166 10948 22204
rect 11004 22370 11060 22988
rect 11004 22318 11006 22370
rect 11058 22318 11060 22370
rect 11004 21924 11060 22318
rect 11004 21858 11060 21868
rect 11116 21812 11172 23774
rect 11340 23996 11508 24052
rect 11228 23714 11284 23726
rect 11228 23662 11230 23714
rect 11282 23662 11284 23714
rect 11228 22484 11284 23662
rect 11228 22418 11284 22428
rect 11340 22036 11396 23996
rect 11900 23938 11956 24444
rect 11900 23886 11902 23938
rect 11954 23886 11956 23938
rect 11452 23828 11508 23838
rect 11676 23828 11732 23838
rect 11452 23826 11732 23828
rect 11452 23774 11454 23826
rect 11506 23774 11678 23826
rect 11730 23774 11732 23826
rect 11452 23772 11732 23774
rect 11452 23762 11508 23772
rect 11676 23762 11732 23772
rect 11788 23604 11844 23614
rect 11564 23266 11620 23278
rect 11564 23214 11566 23266
rect 11618 23214 11620 23266
rect 11564 22372 11620 23214
rect 11788 22596 11844 23548
rect 11900 23492 11956 23886
rect 11900 23426 11956 23436
rect 11788 22530 11844 22540
rect 12012 22596 12068 25228
rect 12236 24612 12292 25452
rect 12348 25394 12404 25406
rect 12348 25342 12350 25394
rect 12402 25342 12404 25394
rect 12348 24836 12404 25342
rect 12460 25284 12516 25294
rect 12460 25190 12516 25228
rect 12348 24770 12404 24780
rect 12460 24612 12516 24622
rect 12236 24610 12516 24612
rect 12236 24558 12462 24610
rect 12514 24558 12516 24610
rect 12236 24556 12516 24558
rect 12460 24546 12516 24556
rect 12236 24164 12292 24174
rect 12236 24070 12292 24108
rect 12460 24164 12516 24174
rect 12572 24164 12628 25452
rect 12684 25506 12740 26236
rect 12796 26180 12852 26190
rect 12796 26086 12852 26124
rect 12684 25454 12686 25506
rect 12738 25454 12740 25506
rect 12684 24948 12740 25454
rect 12908 25394 12964 26684
rect 13132 26516 13188 26526
rect 13020 26514 13188 26516
rect 13020 26462 13134 26514
rect 13186 26462 13188 26514
rect 13020 26460 13188 26462
rect 13020 25508 13076 26460
rect 13132 26450 13188 26460
rect 13020 25442 13076 25452
rect 13132 26290 13188 26302
rect 13132 26238 13134 26290
rect 13186 26238 13188 26290
rect 12908 25342 12910 25394
rect 12962 25342 12964 25394
rect 12908 25060 12964 25342
rect 13132 25396 13188 26238
rect 13132 25284 13188 25340
rect 12908 24994 12964 25004
rect 13020 25228 13188 25284
rect 13356 26066 13412 26078
rect 13356 26014 13358 26066
rect 13410 26014 13412 26066
rect 12684 24882 12740 24892
rect 13020 24722 13076 25228
rect 13020 24670 13022 24722
rect 13074 24670 13076 24722
rect 13020 24658 13076 24670
rect 13132 24948 13188 24958
rect 13132 24834 13188 24892
rect 13356 24948 13412 26014
rect 13468 26068 13524 28588
rect 13468 25506 13524 26012
rect 13468 25454 13470 25506
rect 13522 25454 13524 25506
rect 13468 25442 13524 25454
rect 13580 25284 13636 34636
rect 13804 34626 13860 34636
rect 14028 34356 14084 34366
rect 14028 34242 14084 34300
rect 14028 34190 14030 34242
rect 14082 34190 14084 34242
rect 14028 34178 14084 34190
rect 14140 34020 14196 35758
rect 13916 33964 14196 34020
rect 13804 33124 13860 33134
rect 13916 33124 13972 33964
rect 14252 33684 14308 36540
rect 14364 35474 14420 37212
rect 14364 35422 14366 35474
rect 14418 35422 14420 35474
rect 14364 35410 14420 35422
rect 14588 35698 14644 37996
rect 14700 37828 14756 37838
rect 14700 37266 14756 37772
rect 14700 37214 14702 37266
rect 14754 37214 14756 37266
rect 14700 37202 14756 37214
rect 14588 35646 14590 35698
rect 14642 35646 14644 35698
rect 14588 34914 14644 35646
rect 14588 34862 14590 34914
rect 14642 34862 14644 34914
rect 14588 34850 14644 34862
rect 14700 36708 14756 36718
rect 13804 33122 13972 33124
rect 13804 33070 13806 33122
rect 13858 33070 13972 33122
rect 13804 33068 13972 33070
rect 14028 33628 14308 33684
rect 14476 34802 14532 34814
rect 14476 34750 14478 34802
rect 14530 34750 14532 34802
rect 14028 33346 14084 33628
rect 14476 33572 14532 34750
rect 14140 33516 14532 33572
rect 14140 33458 14196 33516
rect 14140 33406 14142 33458
rect 14194 33406 14196 33458
rect 14140 33394 14196 33406
rect 14028 33294 14030 33346
rect 14082 33294 14084 33346
rect 13804 33012 13860 33068
rect 13804 32946 13860 32956
rect 14028 32788 14084 33294
rect 14588 33346 14644 33358
rect 14588 33294 14590 33346
rect 14642 33294 14644 33346
rect 14252 33124 14308 33134
rect 14252 33030 14308 33068
rect 14588 33012 14644 33294
rect 14700 33124 14756 36652
rect 14812 34692 14868 38220
rect 14924 36260 14980 40124
rect 15036 39620 15092 39630
rect 15036 38052 15092 39564
rect 15260 39620 15316 39630
rect 15260 39526 15316 39564
rect 15260 38276 15316 38286
rect 15148 38052 15204 38062
rect 15036 38050 15204 38052
rect 15036 37998 15150 38050
rect 15202 37998 15204 38050
rect 15036 37996 15204 37998
rect 15148 37940 15204 37996
rect 15148 37044 15204 37884
rect 15148 36978 15204 36988
rect 14924 36194 14980 36204
rect 15148 36708 15204 36718
rect 15148 35698 15204 36652
rect 15148 35646 15150 35698
rect 15202 35646 15204 35698
rect 15148 35634 15204 35646
rect 15260 35588 15316 38220
rect 15372 36820 15428 41244
rect 15484 41186 15540 41580
rect 15484 41134 15486 41186
rect 15538 41134 15540 41186
rect 15484 40964 15540 41134
rect 15596 41076 15652 41918
rect 15708 41300 15764 49196
rect 15932 48802 15988 48814
rect 15932 48750 15934 48802
rect 15986 48750 15988 48802
rect 15932 48244 15988 48750
rect 15932 48178 15988 48188
rect 15820 48132 15876 48142
rect 15820 45108 15876 48076
rect 16044 47458 16100 49420
rect 16156 48580 16212 48590
rect 16156 47570 16212 48524
rect 16268 47796 16324 50372
rect 16380 49924 16436 49934
rect 16380 49830 16436 49868
rect 16492 49922 16548 49934
rect 16492 49870 16494 49922
rect 16546 49870 16548 49922
rect 16268 47730 16324 47740
rect 16380 49700 16436 49710
rect 16156 47518 16158 47570
rect 16210 47518 16212 47570
rect 16156 47506 16212 47518
rect 16044 47406 16046 47458
rect 16098 47406 16100 47458
rect 16044 47394 16100 47406
rect 16268 47348 16324 47358
rect 16268 47254 16324 47292
rect 16380 47068 16436 49644
rect 16492 48356 16548 49870
rect 16604 49922 16660 50316
rect 16828 50372 16884 50382
rect 16828 50370 16996 50372
rect 16828 50318 16830 50370
rect 16882 50318 16996 50370
rect 16828 50316 16996 50318
rect 16828 50306 16884 50316
rect 16716 50036 16772 50046
rect 16716 49942 16772 49980
rect 16604 49870 16606 49922
rect 16658 49870 16660 49922
rect 16604 49028 16660 49870
rect 16828 49810 16884 49822
rect 16828 49758 16830 49810
rect 16882 49758 16884 49810
rect 16828 49364 16884 49758
rect 16828 49298 16884 49308
rect 16940 49140 16996 50316
rect 17052 49588 17108 51660
rect 17164 51650 17220 51660
rect 17276 51604 17332 51998
rect 17276 51538 17332 51548
rect 17388 51940 17444 51950
rect 17388 51490 17444 51884
rect 17500 51602 17556 52556
rect 17612 52388 17668 52398
rect 17612 52274 17668 52332
rect 17612 52222 17614 52274
rect 17666 52222 17668 52274
rect 17612 52210 17668 52222
rect 17500 51550 17502 51602
rect 17554 51550 17556 51602
rect 17500 51538 17556 51550
rect 17612 52052 17668 52062
rect 17388 51438 17390 51490
rect 17442 51438 17444 51490
rect 17388 51426 17444 51438
rect 17500 51156 17556 51166
rect 17612 51156 17668 51996
rect 17500 51154 17668 51156
rect 17500 51102 17502 51154
rect 17554 51102 17668 51154
rect 17500 51100 17668 51102
rect 17500 51090 17556 51100
rect 17724 50428 17780 56590
rect 17836 55524 17892 56812
rect 18172 56754 18228 56766
rect 18172 56702 18174 56754
rect 18226 56702 18228 56754
rect 17948 56644 18004 56654
rect 17948 56642 18116 56644
rect 17948 56590 17950 56642
rect 18002 56590 18116 56642
rect 17948 56588 18116 56590
rect 17948 56578 18004 56588
rect 17948 55524 18004 55534
rect 17836 55468 17948 55524
rect 17948 55458 18004 55468
rect 17948 54516 18004 54526
rect 17948 54422 18004 54460
rect 17836 54404 17892 54414
rect 17836 54310 17892 54348
rect 17836 54180 17892 54190
rect 17836 53618 17892 54124
rect 17836 53566 17838 53618
rect 17890 53566 17892 53618
rect 17836 53554 17892 53566
rect 18060 53508 18116 56588
rect 18172 56196 18228 56702
rect 18284 56644 18340 56654
rect 18284 56550 18340 56588
rect 18172 56140 18340 56196
rect 18172 55970 18228 55982
rect 18172 55918 18174 55970
rect 18226 55918 18228 55970
rect 18172 55300 18228 55918
rect 18284 55524 18340 56140
rect 18284 55458 18340 55468
rect 18396 55410 18452 56924
rect 18508 56868 18564 56878
rect 18508 56774 18564 56812
rect 18732 56756 18788 56766
rect 19180 56756 19236 57598
rect 19292 57540 19348 57550
rect 19292 57446 19348 57484
rect 19404 57316 19460 57708
rect 19404 57250 19460 57260
rect 18732 56754 19012 56756
rect 18732 56702 18734 56754
rect 18786 56702 19012 56754
rect 18732 56700 19012 56702
rect 18732 56690 18788 56700
rect 18956 56308 19012 56700
rect 19180 56690 19236 56700
rect 19404 56978 19460 56990
rect 19404 56926 19406 56978
rect 19458 56926 19460 56978
rect 18508 56084 18564 56094
rect 18508 55990 18564 56028
rect 18396 55358 18398 55410
rect 18450 55358 18452 55410
rect 18396 55346 18452 55358
rect 18732 55300 18788 55310
rect 18172 55244 18340 55300
rect 18060 53442 18116 53452
rect 18172 55076 18228 55086
rect 18172 53730 18228 55020
rect 18284 54852 18340 55244
rect 18284 54786 18340 54796
rect 18620 55188 18676 55198
rect 18172 53678 18174 53730
rect 18226 53678 18228 53730
rect 18060 53284 18116 53294
rect 17836 53060 17892 53070
rect 17836 52966 17892 53004
rect 17612 50372 17780 50428
rect 17948 51378 18004 51390
rect 17948 51326 17950 51378
rect 18002 51326 18004 51378
rect 17612 49924 17668 50372
rect 17052 49532 17556 49588
rect 17388 49364 17444 49374
rect 16940 49084 17332 49140
rect 16604 48962 16660 48972
rect 16940 48914 16996 48926
rect 16940 48862 16942 48914
rect 16994 48862 16996 48914
rect 16492 48290 16548 48300
rect 16604 48804 16660 48814
rect 16940 48804 16996 48862
rect 16604 48242 16660 48748
rect 16604 48190 16606 48242
rect 16658 48190 16660 48242
rect 16604 48178 16660 48190
rect 16716 48748 16996 48804
rect 16716 48020 16772 48748
rect 16492 48018 16772 48020
rect 16492 47966 16718 48018
rect 16770 47966 16772 48018
rect 16492 47964 16772 47966
rect 16492 47458 16548 47964
rect 16716 47954 16772 47964
rect 16492 47406 16494 47458
rect 16546 47406 16548 47458
rect 16492 47394 16548 47406
rect 16604 47796 16660 47806
rect 16604 47346 16660 47740
rect 16604 47294 16606 47346
rect 16658 47294 16660 47346
rect 16604 47282 16660 47294
rect 16156 47012 16212 47022
rect 16380 47012 16772 47068
rect 15932 46788 15988 46798
rect 15932 46694 15988 46732
rect 16156 46676 16212 46956
rect 16156 46582 16212 46620
rect 16268 46564 16324 46574
rect 16492 46564 16548 46574
rect 16268 46470 16324 46508
rect 16380 46562 16548 46564
rect 16380 46510 16494 46562
rect 16546 46510 16548 46562
rect 16380 46508 16548 46510
rect 16268 45108 16324 45118
rect 15820 45106 16324 45108
rect 15820 45054 16270 45106
rect 16322 45054 16324 45106
rect 15820 45052 16324 45054
rect 16268 44548 16324 45052
rect 16268 44482 16324 44492
rect 16380 44324 16436 46508
rect 16492 46498 16548 46508
rect 16716 46340 16772 47012
rect 17276 46788 17332 49084
rect 16716 46274 16772 46284
rect 16828 46562 16884 46574
rect 16828 46510 16830 46562
rect 16882 46510 16884 46562
rect 16828 46116 16884 46510
rect 16828 46050 16884 46060
rect 16716 45780 16772 45790
rect 16380 44258 16436 44268
rect 16492 45778 16772 45780
rect 16492 45726 16718 45778
rect 16770 45726 16772 45778
rect 16492 45724 16772 45726
rect 16156 43652 16212 43662
rect 16492 43652 16548 45724
rect 16716 45714 16772 45724
rect 17276 45780 17332 46732
rect 17388 46676 17444 49308
rect 17500 47458 17556 49532
rect 17612 49028 17668 49868
rect 17612 48934 17668 48972
rect 17500 47406 17502 47458
rect 17554 47406 17556 47458
rect 17500 47394 17556 47406
rect 17948 48914 18004 51326
rect 18060 49700 18116 53228
rect 18172 52388 18228 53678
rect 18508 54740 18564 54750
rect 18508 54626 18564 54684
rect 18508 54574 18510 54626
rect 18562 54574 18564 54626
rect 18508 54180 18564 54574
rect 18620 54516 18676 55132
rect 18620 54422 18676 54460
rect 18508 53732 18564 54124
rect 18508 53676 18676 53732
rect 18508 53506 18564 53518
rect 18508 53454 18510 53506
rect 18562 53454 18564 53506
rect 18508 53396 18564 53454
rect 18508 53330 18564 53340
rect 18620 53060 18676 53676
rect 18732 53730 18788 55244
rect 18956 54514 19012 56252
rect 19180 55186 19236 55198
rect 19180 55134 19182 55186
rect 19234 55134 19236 55186
rect 19180 54740 19236 55134
rect 19180 54674 19236 54684
rect 18956 54462 18958 54514
rect 19010 54462 19012 54514
rect 18956 54450 19012 54462
rect 18732 53678 18734 53730
rect 18786 53678 18788 53730
rect 18732 53666 18788 53678
rect 18844 53842 18900 53854
rect 18844 53790 18846 53842
rect 18898 53790 18900 53842
rect 18844 53732 18900 53790
rect 18844 53666 18900 53676
rect 19068 53730 19124 53742
rect 19068 53678 19070 53730
rect 19122 53678 19124 53730
rect 18732 53060 18788 53070
rect 18620 53058 18788 53060
rect 18620 53006 18734 53058
rect 18786 53006 18788 53058
rect 18620 53004 18788 53006
rect 18732 52994 18788 53004
rect 19068 52724 19124 53678
rect 19404 53620 19460 56926
rect 19516 56866 19572 58828
rect 20076 58548 20132 59388
rect 20524 59218 20580 59230
rect 20524 59166 20526 59218
rect 20578 59166 20580 59218
rect 20076 58482 20132 58492
rect 20412 58546 20468 58558
rect 20412 58494 20414 58546
rect 20466 58494 20468 58546
rect 19628 58436 19684 58446
rect 19628 58342 19684 58380
rect 19628 58100 19684 58110
rect 19628 57876 19684 58044
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19964 57876 20020 57886
rect 19628 57820 19796 57876
rect 19740 57764 19796 57820
rect 19740 57698 19796 57708
rect 19628 57650 19684 57662
rect 19628 57598 19630 57650
rect 19682 57598 19684 57650
rect 19628 57540 19684 57598
rect 19964 57650 20020 57820
rect 19964 57598 19966 57650
rect 20018 57598 20020 57650
rect 19964 57586 20020 57598
rect 19628 57474 19684 57484
rect 19516 56814 19518 56866
rect 19570 56814 19572 56866
rect 19516 56802 19572 56814
rect 20188 56868 20244 56878
rect 20244 56812 20356 56868
rect 20188 56802 20244 56812
rect 19740 56756 19796 56766
rect 19740 56662 19796 56700
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 20188 56420 20244 56430
rect 20188 56196 20244 56364
rect 19740 56082 19796 56094
rect 19740 56030 19742 56082
rect 19794 56030 19796 56082
rect 19516 55412 19572 55422
rect 19516 54628 19572 55356
rect 19740 55188 19796 56030
rect 20188 56082 20244 56140
rect 20188 56030 20190 56082
rect 20242 56030 20244 56082
rect 20188 56018 20244 56030
rect 19740 55122 19796 55132
rect 20188 55524 20244 55534
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19516 54514 19572 54572
rect 19516 54462 19518 54514
rect 19570 54462 19572 54514
rect 19516 54450 19572 54462
rect 20188 54514 20244 55468
rect 20188 54462 20190 54514
rect 20242 54462 20244 54514
rect 19852 54404 19908 54414
rect 19852 54310 19908 54348
rect 19404 53554 19460 53564
rect 19516 54292 19572 54302
rect 19068 52658 19124 52668
rect 19180 53508 19236 53518
rect 18172 52322 18228 52332
rect 18844 51828 18900 51838
rect 18396 51716 18452 51726
rect 18060 49634 18116 49644
rect 18284 51490 18340 51502
rect 18284 51438 18286 51490
rect 18338 51438 18340 51490
rect 18284 49364 18340 51438
rect 18284 49298 18340 49308
rect 18396 50484 18452 51660
rect 18844 51492 18900 51772
rect 18844 51378 18900 51436
rect 18844 51326 18846 51378
rect 18898 51326 18900 51378
rect 18844 51314 18900 51326
rect 18956 51602 19012 51614
rect 18956 51550 18958 51602
rect 19010 51550 19012 51602
rect 18732 50484 18788 50494
rect 18396 50482 18788 50484
rect 18396 50430 18734 50482
rect 18786 50430 18788 50482
rect 18396 50428 18788 50430
rect 18396 49922 18452 50428
rect 18732 50418 18788 50428
rect 18396 49870 18398 49922
rect 18450 49870 18452 49922
rect 18396 49140 18452 49870
rect 18956 49924 19012 51550
rect 18956 49858 19012 49868
rect 18396 49074 18452 49084
rect 18508 49588 18564 49598
rect 17948 48862 17950 48914
rect 18002 48862 18004 48914
rect 17948 47572 18004 48862
rect 18284 49028 18340 49038
rect 18060 48244 18116 48254
rect 18116 48188 18228 48244
rect 18060 48150 18116 48188
rect 18060 47572 18116 47582
rect 17948 47516 18060 47572
rect 17948 47012 18004 47516
rect 18060 47506 18116 47516
rect 18172 47460 18228 48188
rect 18284 48242 18340 48972
rect 18508 49026 18564 49532
rect 18508 48974 18510 49026
rect 18562 48974 18564 49026
rect 18508 48804 18564 48974
rect 18508 48738 18564 48748
rect 18284 48190 18286 48242
rect 18338 48190 18340 48242
rect 18284 48178 18340 48190
rect 18508 48356 18564 48366
rect 18172 47394 18228 47404
rect 18284 48020 18340 48030
rect 17948 46946 18004 46956
rect 18060 47346 18116 47358
rect 18060 47294 18062 47346
rect 18114 47294 18116 47346
rect 18060 47236 18116 47294
rect 18284 47236 18340 47964
rect 18060 47180 18340 47236
rect 17724 46788 17780 46798
rect 17724 46694 17780 46732
rect 17948 46786 18004 46798
rect 17948 46734 17950 46786
rect 18002 46734 18004 46786
rect 17388 46610 17444 46620
rect 17724 46564 17780 46574
rect 17612 46004 17668 46014
rect 17276 45714 17332 45724
rect 17500 45948 17612 46004
rect 17388 45556 17444 45566
rect 17388 45330 17444 45500
rect 17388 45278 17390 45330
rect 17442 45278 17444 45330
rect 17388 45266 17444 45278
rect 16716 44884 16772 44894
rect 16716 44790 16772 44828
rect 16716 44436 16772 44446
rect 16212 43596 16548 43652
rect 16604 44434 16772 44436
rect 16604 44382 16718 44434
rect 16770 44382 16772 44434
rect 16604 44380 16772 44382
rect 16156 43558 16212 43596
rect 15932 43538 15988 43550
rect 16604 43540 16660 44380
rect 16716 44370 16772 44380
rect 17388 44324 17444 44334
rect 17500 44324 17556 45948
rect 17612 45938 17668 45948
rect 17724 45892 17780 46508
rect 17612 45780 17668 45790
rect 17612 45330 17668 45724
rect 17612 45278 17614 45330
rect 17666 45278 17668 45330
rect 17612 44772 17668 45278
rect 17724 45218 17780 45836
rect 17724 45166 17726 45218
rect 17778 45166 17780 45218
rect 17724 45154 17780 45166
rect 17724 44996 17780 45006
rect 17724 44994 17892 44996
rect 17724 44942 17726 44994
rect 17778 44942 17892 44994
rect 17724 44940 17892 44942
rect 17724 44930 17780 44940
rect 17612 44716 17780 44772
rect 17500 44268 17668 44324
rect 17164 44210 17220 44222
rect 17164 44158 17166 44210
rect 17218 44158 17220 44210
rect 17052 44100 17108 44110
rect 15932 43486 15934 43538
rect 15986 43486 15988 43538
rect 15932 43428 15988 43486
rect 16268 43538 16660 43540
rect 16268 43486 16606 43538
rect 16658 43486 16660 43538
rect 16268 43484 16660 43486
rect 16268 43428 16324 43484
rect 16604 43474 16660 43484
rect 16716 44098 17108 44100
rect 16716 44046 17054 44098
rect 17106 44046 17108 44098
rect 16716 44044 17108 44046
rect 15932 43372 16324 43428
rect 16716 42868 16772 44044
rect 17052 44034 17108 44044
rect 16828 43652 16884 43662
rect 16828 43650 16996 43652
rect 16828 43598 16830 43650
rect 16882 43598 16996 43650
rect 16828 43596 16996 43598
rect 16828 43586 16884 43596
rect 16156 42812 16772 42868
rect 16156 41970 16212 42812
rect 16268 42644 16324 42654
rect 16268 42642 16660 42644
rect 16268 42590 16270 42642
rect 16322 42590 16660 42642
rect 16268 42588 16660 42590
rect 16268 42578 16324 42588
rect 16156 41918 16158 41970
rect 16210 41918 16212 41970
rect 16156 41906 16212 41918
rect 16268 42196 16324 42206
rect 16044 41860 16100 41870
rect 15708 41234 15764 41244
rect 15932 41746 15988 41758
rect 15932 41694 15934 41746
rect 15986 41694 15988 41746
rect 15820 41186 15876 41198
rect 15820 41134 15822 41186
rect 15874 41134 15876 41186
rect 15820 41076 15876 41134
rect 15596 41020 15876 41076
rect 15484 40898 15540 40908
rect 15596 40516 15652 40526
rect 15484 40514 15652 40516
rect 15484 40462 15598 40514
rect 15650 40462 15652 40514
rect 15484 40460 15652 40462
rect 15484 40292 15540 40460
rect 15596 40450 15652 40460
rect 15484 40226 15540 40236
rect 15708 40402 15764 40414
rect 15708 40350 15710 40402
rect 15762 40350 15764 40402
rect 15596 40178 15652 40190
rect 15596 40126 15598 40178
rect 15650 40126 15652 40178
rect 15596 38276 15652 40126
rect 15708 38668 15764 40350
rect 15820 39620 15876 41020
rect 15820 39554 15876 39564
rect 15932 41186 15988 41694
rect 15932 41134 15934 41186
rect 15986 41134 15988 41186
rect 15932 39508 15988 41134
rect 16044 41186 16100 41804
rect 16268 41748 16324 42140
rect 16604 42194 16660 42588
rect 16604 42142 16606 42194
rect 16658 42142 16660 42194
rect 16604 42130 16660 42142
rect 16044 41134 16046 41186
rect 16098 41134 16100 41186
rect 16044 41122 16100 41134
rect 16156 41692 16324 41748
rect 16492 41748 16548 41758
rect 16492 41746 16660 41748
rect 16492 41694 16494 41746
rect 16546 41694 16660 41746
rect 16492 41692 16660 41694
rect 15932 39442 15988 39452
rect 16044 40964 16100 40974
rect 16044 39506 16100 40908
rect 16044 39454 16046 39506
rect 16098 39454 16100 39506
rect 16044 39442 16100 39454
rect 16156 40292 16212 41692
rect 16492 41682 16548 41692
rect 16268 40964 16324 40974
rect 16268 40870 16324 40908
rect 16604 40964 16660 41692
rect 16716 41186 16772 42812
rect 16716 41134 16718 41186
rect 16770 41134 16772 41186
rect 16716 41122 16772 41134
rect 16828 41970 16884 41982
rect 16828 41918 16830 41970
rect 16882 41918 16884 41970
rect 16828 40964 16884 41918
rect 16940 41748 16996 43596
rect 17164 41860 17220 44158
rect 17388 44100 17444 44268
rect 17500 44100 17556 44110
rect 17388 44098 17556 44100
rect 17388 44046 17502 44098
rect 17554 44046 17556 44098
rect 17388 44044 17556 44046
rect 17500 44034 17556 44044
rect 17164 41794 17220 41804
rect 17276 41970 17332 41982
rect 17276 41918 17278 41970
rect 17330 41918 17332 41970
rect 16940 41682 16996 41692
rect 16940 41188 16996 41198
rect 16940 41094 16996 41132
rect 17164 41076 17220 41086
rect 17276 41076 17332 41918
rect 17500 41972 17556 41982
rect 17500 41878 17556 41916
rect 17612 41970 17668 44268
rect 17724 43538 17780 44716
rect 17724 43486 17726 43538
rect 17778 43486 17780 43538
rect 17724 43474 17780 43486
rect 17612 41918 17614 41970
rect 17666 41918 17668 41970
rect 17612 41188 17668 41918
rect 17612 41122 17668 41132
rect 17052 41074 17332 41076
rect 17052 41022 17166 41074
rect 17218 41022 17332 41074
rect 17052 41020 17332 41022
rect 16940 40964 16996 40974
rect 16828 40962 16996 40964
rect 16828 40910 16942 40962
rect 16994 40910 16996 40962
rect 16828 40908 16996 40910
rect 16604 40898 16660 40908
rect 16940 40898 16996 40908
rect 16828 40404 16884 40414
rect 16828 40402 16996 40404
rect 16828 40350 16830 40402
rect 16882 40350 16996 40402
rect 16828 40348 16996 40350
rect 16828 40338 16884 40348
rect 16268 40292 16324 40302
rect 16156 40290 16324 40292
rect 16156 40238 16270 40290
rect 16322 40238 16324 40290
rect 16156 40236 16324 40238
rect 16156 39060 16212 40236
rect 16268 40226 16324 40236
rect 16492 40178 16548 40190
rect 16492 40126 16494 40178
rect 16546 40126 16548 40178
rect 16492 39172 16548 40126
rect 16828 40180 16884 40190
rect 16828 40068 16884 40124
rect 16716 40012 16884 40068
rect 16716 39620 16772 40012
rect 16828 39844 16884 39854
rect 16828 39750 16884 39788
rect 16940 39620 16996 40348
rect 16716 39564 16884 39620
rect 16604 39508 16660 39518
rect 16604 39414 16660 39452
rect 16156 39004 16324 39060
rect 16268 38946 16324 39004
rect 16268 38894 16270 38946
rect 16322 38894 16324 38946
rect 16268 38882 16324 38894
rect 16156 38836 16212 38846
rect 15708 38612 15876 38668
rect 15596 38210 15652 38220
rect 15596 38052 15652 38062
rect 15596 37958 15652 37996
rect 15708 37940 15764 37950
rect 15708 37490 15764 37884
rect 15708 37438 15710 37490
rect 15762 37438 15764 37490
rect 15708 37426 15764 37438
rect 15820 37490 15876 38612
rect 15820 37438 15822 37490
rect 15874 37438 15876 37490
rect 15820 37426 15876 37438
rect 15932 38052 15988 38062
rect 15932 37490 15988 37996
rect 15932 37438 15934 37490
rect 15986 37438 15988 37490
rect 15932 37426 15988 37438
rect 16044 37378 16100 37390
rect 16044 37326 16046 37378
rect 16098 37326 16100 37378
rect 16044 37268 16100 37326
rect 16156 37378 16212 38780
rect 16492 38834 16548 39116
rect 16828 39058 16884 39564
rect 16940 39554 16996 39564
rect 16828 39006 16830 39058
rect 16882 39006 16884 39058
rect 16828 38994 16884 39006
rect 16492 38782 16494 38834
rect 16546 38782 16548 38834
rect 16492 38770 16548 38782
rect 16156 37326 16158 37378
rect 16210 37326 16212 37378
rect 16156 37314 16212 37326
rect 16268 38276 16324 38286
rect 16044 37202 16100 37212
rect 15372 36764 15540 36820
rect 15372 36596 15428 36606
rect 15372 35698 15428 36540
rect 15372 35646 15374 35698
rect 15426 35646 15428 35698
rect 15372 35634 15428 35646
rect 15260 34914 15316 35532
rect 15260 34862 15262 34914
rect 15314 34862 15316 34914
rect 15260 34850 15316 34862
rect 15372 35252 15428 35262
rect 15372 34802 15428 35196
rect 15372 34750 15374 34802
rect 15426 34750 15428 34802
rect 15372 34738 15428 34750
rect 14812 34626 14868 34636
rect 15372 34468 15428 34478
rect 15036 34242 15092 34254
rect 15036 34190 15038 34242
rect 15090 34190 15092 34242
rect 15036 34132 15092 34190
rect 15372 34242 15428 34412
rect 15484 34354 15540 36764
rect 16044 36372 16100 36382
rect 16044 36278 16100 36316
rect 16268 36260 16324 38220
rect 17052 36596 17108 41020
rect 17164 41010 17220 41020
rect 17724 40516 17780 40526
rect 17388 40514 17780 40516
rect 17388 40462 17726 40514
rect 17778 40462 17780 40514
rect 17388 40460 17780 40462
rect 17164 39394 17220 39406
rect 17164 39342 17166 39394
rect 17218 39342 17220 39394
rect 17164 38948 17220 39342
rect 17164 38882 17220 38892
rect 17276 39172 17332 39182
rect 17276 38274 17332 39116
rect 17388 39060 17444 40460
rect 17724 40450 17780 40460
rect 17612 39508 17668 39518
rect 17612 39414 17668 39452
rect 17612 39284 17668 39294
rect 17500 39060 17556 39070
rect 17388 39058 17556 39060
rect 17388 39006 17502 39058
rect 17554 39006 17556 39058
rect 17388 39004 17556 39006
rect 17500 38994 17556 39004
rect 17612 38946 17668 39228
rect 17612 38894 17614 38946
rect 17666 38894 17668 38946
rect 17276 38222 17278 38274
rect 17330 38222 17332 38274
rect 17276 38210 17332 38222
rect 17388 38834 17444 38846
rect 17388 38782 17390 38834
rect 17442 38782 17444 38834
rect 17164 36596 17220 36606
rect 17052 36540 17164 36596
rect 17164 36530 17220 36540
rect 16268 36194 16324 36204
rect 16828 36482 16884 36494
rect 16828 36430 16830 36482
rect 16882 36430 16884 36482
rect 16828 35924 16884 36430
rect 17388 35924 17444 38782
rect 17500 37268 17556 37278
rect 17500 37174 17556 37212
rect 17500 36596 17556 36606
rect 17500 36502 17556 36540
rect 17612 36482 17668 38894
rect 17724 38948 17780 38958
rect 17724 38854 17780 38892
rect 17836 38946 17892 44940
rect 17948 43428 18004 46734
rect 18060 45668 18116 47180
rect 18508 46900 18564 48300
rect 19180 48244 19236 53452
rect 19292 53506 19348 53518
rect 19292 53454 19294 53506
rect 19346 53454 19348 53506
rect 19292 53172 19348 53454
rect 19292 53106 19348 53116
rect 19516 51268 19572 54236
rect 19852 54180 19908 54190
rect 19852 53730 19908 54124
rect 20188 53732 20244 54462
rect 19852 53678 19854 53730
rect 19906 53678 19908 53730
rect 19852 53666 19908 53678
rect 20076 53676 20244 53732
rect 20300 54626 20356 56812
rect 20300 54574 20302 54626
rect 20354 54574 20356 54626
rect 20076 53620 20132 53676
rect 20076 53554 20132 53564
rect 20188 53506 20244 53518
rect 20188 53454 20190 53506
rect 20242 53454 20244 53506
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19964 53172 20020 53182
rect 20188 53172 20244 53454
rect 20300 53508 20356 54574
rect 20412 53620 20468 58494
rect 20524 57316 20580 59166
rect 20860 59220 20916 59836
rect 22540 59892 22596 59902
rect 20860 59154 20916 59164
rect 20972 59778 21028 59790
rect 21196 59780 21252 59790
rect 20972 59726 20974 59778
rect 21026 59726 21028 59778
rect 20972 58884 21028 59726
rect 20972 58818 21028 58828
rect 21084 59778 21252 59780
rect 21084 59726 21198 59778
rect 21250 59726 21252 59778
rect 21084 59724 21252 59726
rect 21084 58324 21140 59724
rect 21196 59714 21252 59724
rect 22092 59778 22148 59790
rect 22092 59726 22094 59778
rect 22146 59726 22148 59778
rect 22092 59668 22148 59726
rect 22092 59442 22148 59612
rect 22092 59390 22094 59442
rect 22146 59390 22148 59442
rect 22092 59378 22148 59390
rect 21756 59108 21812 59118
rect 20972 58268 21140 58324
rect 21420 58996 21476 59006
rect 20524 56866 20580 57260
rect 20748 57540 20804 57550
rect 20524 56814 20526 56866
rect 20578 56814 20580 56866
rect 20524 56196 20580 56814
rect 20524 56130 20580 56140
rect 20636 57092 20692 57102
rect 20636 56082 20692 57036
rect 20748 56866 20804 57484
rect 20972 57092 21028 58268
rect 21308 58212 21364 58222
rect 20972 57026 21028 57036
rect 21084 58210 21364 58212
rect 21084 58158 21310 58210
rect 21362 58158 21364 58210
rect 21084 58156 21364 58158
rect 20748 56814 20750 56866
rect 20802 56814 20804 56866
rect 20748 56802 20804 56814
rect 21084 56084 21140 58156
rect 21308 58146 21364 58156
rect 21196 57764 21252 57774
rect 21196 57650 21252 57708
rect 21196 57598 21198 57650
rect 21250 57598 21252 57650
rect 21196 57586 21252 57598
rect 21308 56980 21364 56990
rect 21420 56980 21476 58940
rect 21756 58324 21812 59052
rect 21980 58548 22036 58558
rect 21980 58454 22036 58492
rect 22540 58434 22596 59836
rect 23212 59892 23268 59902
rect 23772 59892 23828 59902
rect 23212 59798 23268 59836
rect 23548 59890 23828 59892
rect 23548 59838 23774 59890
rect 23826 59838 23828 59890
rect 23548 59836 23828 59838
rect 23436 58996 23492 59006
rect 23436 58902 23492 58940
rect 22540 58382 22542 58434
rect 22594 58382 22596 58434
rect 22540 58370 22596 58382
rect 22876 58434 22932 58446
rect 22876 58382 22878 58434
rect 22930 58382 22932 58434
rect 21756 58268 22036 58324
rect 21644 58210 21700 58222
rect 21644 58158 21646 58210
rect 21698 58158 21700 58210
rect 21308 56978 21476 56980
rect 21308 56926 21310 56978
rect 21362 56926 21476 56978
rect 21308 56924 21476 56926
rect 21532 58100 21588 58110
rect 21308 56914 21364 56924
rect 21420 56756 21476 56766
rect 21532 56756 21588 58044
rect 21644 56868 21700 58158
rect 21868 57652 21924 57662
rect 21868 57558 21924 57596
rect 21644 56802 21700 56812
rect 21420 56754 21588 56756
rect 21420 56702 21422 56754
rect 21474 56702 21588 56754
rect 21420 56700 21588 56702
rect 21980 56754 22036 58268
rect 22092 57652 22148 57662
rect 22092 57204 22148 57596
rect 22092 56866 22148 57148
rect 22092 56814 22094 56866
rect 22146 56814 22148 56866
rect 22092 56802 22148 56814
rect 22764 56868 22820 56878
rect 22876 56868 22932 58382
rect 23212 57428 23268 57438
rect 23212 57334 23268 57372
rect 22764 56866 22932 56868
rect 22764 56814 22766 56866
rect 22818 56814 22932 56866
rect 22764 56812 22932 56814
rect 23548 56980 23604 59836
rect 23772 59826 23828 59836
rect 23884 59890 23940 59948
rect 23884 59838 23886 59890
rect 23938 59838 23940 59890
rect 23884 59826 23940 59838
rect 24108 59780 24164 59790
rect 24108 59778 24388 59780
rect 24108 59726 24110 59778
rect 24162 59726 24388 59778
rect 24108 59724 24388 59726
rect 24108 59714 24164 59724
rect 24332 59330 24388 59724
rect 24444 59668 24500 59948
rect 25004 59778 25060 59790
rect 25004 59726 25006 59778
rect 25058 59726 25060 59778
rect 24444 59612 24724 59668
rect 24332 59278 24334 59330
rect 24386 59278 24388 59330
rect 24332 59266 24388 59278
rect 23660 59220 23716 59230
rect 23660 57428 23716 59164
rect 24556 59220 24612 59230
rect 24556 59126 24612 59164
rect 23772 59108 23828 59118
rect 23772 59106 24276 59108
rect 23772 59054 23774 59106
rect 23826 59054 24276 59106
rect 23772 59052 24276 59054
rect 23772 59042 23828 59052
rect 23884 58884 23940 58894
rect 23940 58828 24052 58884
rect 23884 58818 23940 58828
rect 23884 58548 23940 58558
rect 23884 57650 23940 58492
rect 23884 57598 23886 57650
rect 23938 57598 23940 57650
rect 23884 57586 23940 57598
rect 23660 57372 23940 57428
rect 21980 56702 21982 56754
rect 22034 56702 22036 56754
rect 21420 56690 21476 56700
rect 21980 56690 22036 56702
rect 22764 56644 22820 56812
rect 22764 56578 22820 56588
rect 23100 56642 23156 56654
rect 23100 56590 23102 56642
rect 23154 56590 23156 56642
rect 21196 56308 21252 56318
rect 21196 56214 21252 56252
rect 20636 56030 20638 56082
rect 20690 56030 20692 56082
rect 20636 56018 20692 56030
rect 20860 56082 21140 56084
rect 20860 56030 21086 56082
rect 21138 56030 21140 56082
rect 20860 56028 21140 56030
rect 20636 55524 20692 55534
rect 20860 55524 20916 56028
rect 21084 56018 21140 56028
rect 21868 56194 21924 56206
rect 21868 56142 21870 56194
rect 21922 56142 21924 56194
rect 20636 55522 20916 55524
rect 20636 55470 20638 55522
rect 20690 55470 20916 55522
rect 20636 55468 20916 55470
rect 20636 54180 20692 55468
rect 21868 55300 21924 56142
rect 22988 56194 23044 56206
rect 22988 56142 22990 56194
rect 23042 56142 23044 56194
rect 21868 55234 21924 55244
rect 22092 56084 22148 56094
rect 22428 56084 22484 56094
rect 22092 56082 22484 56084
rect 22092 56030 22094 56082
rect 22146 56030 22430 56082
rect 22482 56030 22484 56082
rect 22092 56028 22484 56030
rect 20860 55188 20916 55198
rect 20860 54738 20916 55132
rect 21980 55076 22036 55086
rect 21980 54982 22036 55020
rect 22092 54964 22148 56028
rect 22428 56018 22484 56028
rect 22764 56082 22820 56094
rect 22764 56030 22766 56082
rect 22818 56030 22820 56082
rect 22092 54740 22148 54908
rect 22652 55636 22708 55646
rect 20860 54686 20862 54738
rect 20914 54686 20916 54738
rect 20860 54674 20916 54686
rect 21980 54684 22148 54740
rect 22204 54740 22260 54750
rect 20972 54628 21028 54638
rect 20972 54534 21028 54572
rect 21532 54626 21588 54638
rect 21532 54574 21534 54626
rect 21586 54574 21588 54626
rect 20636 54114 20692 54124
rect 20748 54516 20804 54526
rect 20748 53842 20804 54460
rect 21532 54516 21588 54574
rect 21868 54626 21924 54638
rect 21868 54574 21870 54626
rect 21922 54574 21924 54626
rect 21532 54450 21588 54460
rect 21644 54514 21700 54526
rect 21868 54516 21924 54574
rect 21644 54462 21646 54514
rect 21698 54462 21700 54514
rect 20748 53790 20750 53842
rect 20802 53790 20804 53842
rect 20748 53778 20804 53790
rect 21308 54402 21364 54414
rect 21308 54350 21310 54402
rect 21362 54350 21364 54402
rect 21308 53844 21364 54350
rect 21308 53778 21364 53788
rect 21532 53732 21588 53742
rect 21532 53638 21588 53676
rect 20412 53564 20916 53620
rect 20300 53442 20356 53452
rect 19964 53170 20244 53172
rect 19964 53118 19966 53170
rect 20018 53118 20244 53170
rect 19964 53116 20244 53118
rect 19964 53060 20020 53116
rect 19964 52994 20020 53004
rect 20412 52946 20468 52958
rect 20412 52894 20414 52946
rect 20466 52894 20468 52946
rect 19740 52836 19796 52846
rect 19740 52274 19796 52780
rect 19740 52222 19742 52274
rect 19794 52222 19796 52274
rect 19740 52210 19796 52222
rect 20412 52052 20468 52894
rect 20636 52946 20692 52958
rect 20636 52894 20638 52946
rect 20690 52894 20692 52946
rect 20524 52836 20580 52846
rect 20524 52742 20580 52780
rect 20636 52612 20692 52894
rect 20636 52546 20692 52556
rect 20524 52276 20580 52286
rect 20524 52162 20580 52220
rect 20524 52110 20526 52162
rect 20578 52110 20580 52162
rect 20524 52098 20580 52110
rect 20412 51986 20468 51996
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 20076 51604 20132 51614
rect 20076 51510 20132 51548
rect 19516 51202 19572 51212
rect 20524 50596 20580 50606
rect 20524 50502 20580 50540
rect 20636 50484 20692 50522
rect 20636 50418 20692 50428
rect 20748 50482 20804 50494
rect 20748 50430 20750 50482
rect 20802 50430 20804 50482
rect 19964 50372 20020 50382
rect 19628 50370 20020 50372
rect 19628 50318 19966 50370
rect 20018 50318 20020 50370
rect 19628 50316 20020 50318
rect 19516 49812 19572 49822
rect 19516 49718 19572 49756
rect 19628 49588 19684 50316
rect 19964 50306 20020 50316
rect 20300 50372 20356 50382
rect 20300 50278 20356 50316
rect 20748 50372 20804 50430
rect 20748 50306 20804 50316
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 20300 50148 20356 50158
rect 20076 49812 20132 49822
rect 19180 48178 19236 48188
rect 19516 49532 19684 49588
rect 19964 49588 20020 49598
rect 19292 47796 19348 47806
rect 18508 46834 18564 46844
rect 18620 47684 18676 47694
rect 18620 46898 18676 47628
rect 18620 46846 18622 46898
rect 18674 46846 18676 46898
rect 18620 46834 18676 46846
rect 19292 46674 19348 47740
rect 19292 46622 19294 46674
rect 19346 46622 19348 46674
rect 19292 46610 19348 46622
rect 18284 46564 18340 46574
rect 18284 46470 18340 46508
rect 18172 46116 18228 46126
rect 18172 46022 18228 46060
rect 18844 46116 18900 46126
rect 18620 45892 18676 45902
rect 18844 45892 18900 46060
rect 18956 46004 19012 46014
rect 18956 45910 19012 45948
rect 18620 45798 18676 45836
rect 18732 45890 18900 45892
rect 18732 45838 18846 45890
rect 18898 45838 18900 45890
rect 18732 45836 18900 45838
rect 18060 45602 18116 45612
rect 17948 43334 18004 43372
rect 18060 45108 18116 45118
rect 18060 44322 18116 45052
rect 18620 44994 18676 45006
rect 18620 44942 18622 44994
rect 18674 44942 18676 44994
rect 18620 44660 18676 44942
rect 18620 44594 18676 44604
rect 18060 44270 18062 44322
rect 18114 44270 18116 44322
rect 17948 42756 18004 42766
rect 18060 42756 18116 44270
rect 18508 43540 18564 43550
rect 18004 42700 18116 42756
rect 18396 43426 18452 43438
rect 18396 43374 18398 43426
rect 18450 43374 18452 43426
rect 18396 43316 18452 43374
rect 17948 42690 18004 42700
rect 17948 42532 18004 42542
rect 18396 42532 18452 43260
rect 18508 43092 18564 43484
rect 18620 43540 18676 43550
rect 18732 43540 18788 45836
rect 18844 45826 18900 45836
rect 18956 44322 19012 44334
rect 18956 44270 18958 44322
rect 19010 44270 19012 44322
rect 18620 43538 18732 43540
rect 18620 43486 18622 43538
rect 18674 43486 18732 43538
rect 18620 43484 18732 43486
rect 18620 43474 18676 43484
rect 18732 43446 18788 43484
rect 18844 44210 18900 44222
rect 18844 44158 18846 44210
rect 18898 44158 18900 44210
rect 18508 43026 18564 43036
rect 17948 42530 18452 42532
rect 17948 42478 17950 42530
rect 18002 42478 18452 42530
rect 17948 42476 18452 42478
rect 17948 42196 18004 42476
rect 17948 42130 18004 42140
rect 18060 42252 18340 42308
rect 17948 41970 18004 41982
rect 17948 41918 17950 41970
rect 18002 41918 18004 41970
rect 17948 41860 18004 41918
rect 17948 41794 18004 41804
rect 17948 40962 18004 40974
rect 17948 40910 17950 40962
rect 18002 40910 18004 40962
rect 17948 40516 18004 40910
rect 17948 40450 18004 40460
rect 18060 40180 18116 42252
rect 18172 42084 18228 42094
rect 18172 41300 18228 42028
rect 18284 42082 18340 42252
rect 18396 42196 18452 42206
rect 18396 42102 18452 42140
rect 18284 42030 18286 42082
rect 18338 42030 18340 42082
rect 18284 42018 18340 42030
rect 18396 41746 18452 41758
rect 18396 41694 18398 41746
rect 18450 41694 18452 41746
rect 18284 41300 18340 41310
rect 18172 41298 18340 41300
rect 18172 41246 18286 41298
rect 18338 41246 18340 41298
rect 18172 41244 18340 41246
rect 18284 41234 18340 41244
rect 18396 41188 18452 41694
rect 18844 41188 18900 44158
rect 18956 43762 19012 44270
rect 19516 44100 19572 49532
rect 19964 49494 20020 49532
rect 19740 49476 19796 49486
rect 19740 49026 19796 49420
rect 19740 48974 19742 49026
rect 19794 48974 19796 49026
rect 19740 48962 19796 48974
rect 20076 49026 20132 49756
rect 20300 49810 20356 50092
rect 20300 49758 20302 49810
rect 20354 49758 20356 49810
rect 20300 49746 20356 49758
rect 20076 48974 20078 49026
rect 20130 48974 20132 49026
rect 20076 48962 20132 48974
rect 20636 48914 20692 48926
rect 20636 48862 20638 48914
rect 20690 48862 20692 48914
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20076 48244 20132 48254
rect 19852 48242 20132 48244
rect 19852 48190 20078 48242
rect 20130 48190 20132 48242
rect 19852 48188 20132 48190
rect 19852 47684 19908 48188
rect 20076 48178 20132 48188
rect 20524 48244 20580 48254
rect 20524 48150 20580 48188
rect 19852 47570 19908 47628
rect 19852 47518 19854 47570
rect 19906 47518 19908 47570
rect 19852 47506 19908 47518
rect 19964 47796 20020 47806
rect 19964 47458 20020 47740
rect 20524 47796 20580 47806
rect 20636 47796 20692 48862
rect 20580 47740 20692 47796
rect 20524 47730 20580 47740
rect 19964 47406 19966 47458
rect 20018 47406 20020 47458
rect 19964 47394 20020 47406
rect 20300 47460 20356 47470
rect 20300 47366 20356 47404
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19740 46900 19796 46910
rect 19740 46786 19796 46844
rect 20188 46900 20244 46910
rect 20244 46844 20356 46900
rect 20188 46834 20244 46844
rect 19740 46734 19742 46786
rect 19794 46734 19796 46786
rect 19740 46722 19796 46734
rect 20076 46004 20132 46014
rect 19740 45890 19796 45902
rect 19740 45838 19742 45890
rect 19794 45838 19796 45890
rect 19740 45780 19796 45838
rect 19740 45714 19796 45724
rect 20076 45668 20132 45948
rect 20076 45602 20132 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20188 45108 20244 45118
rect 20188 45014 20244 45052
rect 20300 44882 20356 46844
rect 20860 45892 20916 53564
rect 21644 53060 21700 54462
rect 21756 54460 21924 54516
rect 21756 53284 21812 54460
rect 21980 54404 22036 54684
rect 22092 54516 22148 54526
rect 22204 54516 22260 54684
rect 22540 54626 22596 54638
rect 22540 54574 22542 54626
rect 22594 54574 22596 54626
rect 22540 54516 22596 54574
rect 22092 54514 22484 54516
rect 22092 54462 22094 54514
rect 22146 54462 22484 54514
rect 22092 54460 22484 54462
rect 22092 54450 22148 54460
rect 21756 53218 21812 53228
rect 21868 54348 22036 54404
rect 21756 53060 21812 53070
rect 21644 53004 21756 53060
rect 21756 52994 21812 53004
rect 21084 52946 21140 52958
rect 21084 52894 21086 52946
rect 21138 52894 21140 52946
rect 21084 52164 21140 52894
rect 21308 52948 21364 52958
rect 21532 52948 21588 52958
rect 21364 52946 21588 52948
rect 21364 52894 21534 52946
rect 21586 52894 21588 52946
rect 21364 52892 21588 52894
rect 21308 52882 21364 52892
rect 21420 52724 21476 52734
rect 21420 52630 21476 52668
rect 21532 52612 21588 52892
rect 21532 52546 21588 52556
rect 21756 52836 21812 52846
rect 21196 52164 21252 52174
rect 21084 52162 21252 52164
rect 21084 52110 21198 52162
rect 21250 52110 21252 52162
rect 21084 52108 21252 52110
rect 21196 52098 21252 52108
rect 21532 52052 21588 52062
rect 21532 52050 21700 52052
rect 21532 51998 21534 52050
rect 21586 51998 21700 52050
rect 21532 51996 21700 51998
rect 21532 51986 21588 51996
rect 21420 51938 21476 51950
rect 21420 51886 21422 51938
rect 21474 51886 21476 51938
rect 21420 51828 21476 51886
rect 21420 51762 21476 51772
rect 21532 51492 21588 51502
rect 21196 51268 21252 51278
rect 21084 48130 21140 48142
rect 21084 48078 21086 48130
rect 21138 48078 21140 48130
rect 21084 47908 21140 48078
rect 21084 47842 21140 47852
rect 20860 45826 20916 45836
rect 21084 46674 21140 46686
rect 21084 46622 21086 46674
rect 21138 46622 21140 46674
rect 20860 45668 20916 45678
rect 20860 45574 20916 45612
rect 20300 44830 20302 44882
rect 20354 44830 20356 44882
rect 20300 44818 20356 44830
rect 20524 45332 20580 45342
rect 20524 44324 20580 45276
rect 20524 44230 20580 44268
rect 20636 45108 20692 45118
rect 20636 44210 20692 45052
rect 21084 45106 21140 46622
rect 21084 45054 21086 45106
rect 21138 45054 21140 45106
rect 21084 44996 21140 45054
rect 20636 44158 20638 44210
rect 20690 44158 20692 44210
rect 19516 44034 19572 44044
rect 20524 44100 20580 44110
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20300 43876 20356 43886
rect 19836 43866 20100 43876
rect 20188 43820 20300 43876
rect 20188 43764 20244 43820
rect 20300 43810 20356 43820
rect 18956 43710 18958 43762
rect 19010 43710 19012 43762
rect 18956 43698 19012 43710
rect 20076 43708 20244 43764
rect 19068 43652 19124 43662
rect 19068 42642 19124 43596
rect 19852 43652 19908 43662
rect 19516 43540 19572 43550
rect 19516 43446 19572 43484
rect 19292 43426 19348 43438
rect 19292 43374 19294 43426
rect 19346 43374 19348 43426
rect 19292 43316 19348 43374
rect 19852 43426 19908 43596
rect 19852 43374 19854 43426
rect 19906 43374 19908 43426
rect 19852 43362 19908 43374
rect 19292 43250 19348 43260
rect 19068 42590 19070 42642
rect 19122 42590 19124 42642
rect 19068 42578 19124 42590
rect 20076 42532 20132 43708
rect 20300 43540 20356 43550
rect 20300 43426 20356 43484
rect 20300 43374 20302 43426
rect 20354 43374 20356 43426
rect 20300 43362 20356 43374
rect 20076 42476 20244 42532
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20188 42196 20244 42476
rect 20076 42140 20244 42196
rect 20300 42530 20356 42542
rect 20300 42478 20302 42530
rect 20354 42478 20356 42530
rect 19180 42082 19236 42094
rect 19180 42030 19182 42082
rect 19234 42030 19236 42082
rect 18396 41132 18564 41188
rect 18844 41132 19012 41188
rect 18172 40962 18228 40974
rect 18172 40910 18174 40962
rect 18226 40910 18228 40962
rect 18172 40404 18228 40910
rect 18396 40964 18452 40974
rect 18396 40870 18452 40908
rect 18172 40338 18228 40348
rect 18060 40114 18116 40124
rect 18396 39620 18452 39630
rect 18508 39620 18564 41132
rect 18844 40964 18900 40974
rect 18844 40870 18900 40908
rect 18508 39564 18676 39620
rect 18396 39526 18452 39564
rect 17948 39508 18004 39518
rect 17948 39172 18004 39452
rect 18508 39396 18564 39406
rect 18508 39302 18564 39340
rect 17948 39106 18004 39116
rect 18508 39060 18564 39070
rect 18620 39060 18676 39564
rect 18508 39058 18676 39060
rect 18508 39006 18510 39058
rect 18562 39006 18676 39058
rect 18508 39004 18676 39006
rect 18508 38994 18564 39004
rect 17836 38894 17838 38946
rect 17890 38894 17892 38946
rect 17836 38882 17892 38894
rect 18732 38834 18788 38846
rect 18732 38782 18734 38834
rect 18786 38782 18788 38834
rect 18620 38722 18676 38734
rect 18620 38670 18622 38722
rect 18674 38670 18676 38722
rect 18508 37940 18564 37950
rect 18508 37846 18564 37884
rect 18620 37378 18676 38670
rect 18620 37326 18622 37378
rect 18674 37326 18676 37378
rect 18620 37314 18676 37326
rect 17948 37268 18004 37278
rect 17948 37174 18004 37212
rect 18620 36820 18676 36830
rect 18732 36820 18788 38782
rect 18676 36764 18788 36820
rect 18284 36596 18340 36606
rect 17612 36430 17614 36482
rect 17666 36430 17668 36482
rect 17612 36418 17668 36430
rect 17836 36594 18340 36596
rect 17836 36542 18286 36594
rect 18338 36542 18340 36594
rect 17836 36540 18340 36542
rect 17612 36148 17668 36158
rect 17500 35924 17556 35934
rect 17388 35922 17556 35924
rect 17388 35870 17502 35922
rect 17554 35870 17556 35922
rect 17388 35868 17556 35870
rect 16828 35858 16884 35868
rect 17500 35858 17556 35868
rect 15596 35700 15652 35710
rect 15596 34914 15652 35644
rect 17388 35698 17444 35710
rect 17388 35646 17390 35698
rect 17442 35646 17444 35698
rect 17052 35476 17108 35486
rect 15596 34862 15598 34914
rect 15650 34862 15652 34914
rect 15596 34850 15652 34862
rect 15820 34916 15876 34926
rect 16044 34916 16100 34926
rect 15820 34914 15988 34916
rect 15820 34862 15822 34914
rect 15874 34862 15988 34914
rect 15820 34860 15988 34862
rect 15820 34850 15876 34860
rect 15484 34302 15486 34354
rect 15538 34302 15540 34354
rect 15484 34290 15540 34302
rect 15372 34190 15374 34242
rect 15426 34190 15428 34242
rect 15092 34076 15204 34132
rect 15036 34038 15092 34076
rect 14700 33058 14756 33068
rect 14588 32946 14644 32956
rect 14924 32900 14980 32910
rect 14028 32732 14308 32788
rect 14028 32450 14084 32462
rect 14028 32398 14030 32450
rect 14082 32398 14084 32450
rect 14028 32116 14084 32398
rect 13804 31220 13860 31230
rect 13692 31108 13748 31118
rect 13692 30994 13748 31052
rect 13692 30942 13694 30994
rect 13746 30942 13748 30994
rect 13692 30436 13748 30942
rect 13692 30370 13748 30380
rect 13804 30210 13860 31164
rect 14028 30996 14084 32060
rect 14028 30930 14084 30940
rect 14028 30660 14084 30670
rect 13804 30158 13806 30210
rect 13858 30158 13860 30210
rect 13804 29428 13860 30158
rect 13804 29362 13860 29372
rect 13916 30604 14028 30660
rect 13692 29314 13748 29326
rect 13692 29262 13694 29314
rect 13746 29262 13748 29314
rect 13692 26908 13748 29262
rect 13804 28756 13860 28766
rect 13916 28756 13972 30604
rect 14028 30594 14084 30604
rect 14140 30436 14196 30446
rect 14252 30436 14308 32732
rect 14812 32564 14868 32574
rect 14924 32564 14980 32844
rect 14812 32562 14924 32564
rect 14812 32510 14814 32562
rect 14866 32510 14924 32562
rect 14812 32508 14924 32510
rect 14812 32498 14868 32508
rect 14924 32470 14980 32508
rect 14476 32340 14532 32350
rect 14476 32338 14644 32340
rect 14476 32286 14478 32338
rect 14530 32286 14644 32338
rect 14476 32284 14644 32286
rect 14476 32274 14532 32284
rect 14364 31780 14420 31790
rect 14364 31686 14420 31724
rect 14476 31778 14532 31790
rect 14476 31726 14478 31778
rect 14530 31726 14532 31778
rect 14476 31108 14532 31726
rect 14476 31042 14532 31052
rect 14588 31780 14644 32284
rect 15148 31892 15204 34076
rect 15260 31892 15316 31902
rect 15148 31836 15260 31892
rect 14588 30770 14644 31724
rect 14588 30718 14590 30770
rect 14642 30718 14644 30770
rect 14588 30706 14644 30718
rect 14700 31668 14756 31678
rect 14700 30660 14756 31612
rect 15148 31668 15204 31678
rect 15036 31444 15092 31454
rect 14812 31108 14868 31118
rect 14812 31014 14868 31052
rect 14700 30604 14868 30660
rect 14252 30380 14644 30436
rect 14140 29650 14196 30380
rect 14140 29598 14142 29650
rect 14194 29598 14196 29650
rect 14140 29586 14196 29598
rect 14252 30210 14308 30222
rect 14252 30158 14254 30210
rect 14306 30158 14308 30210
rect 14252 29428 14308 30158
rect 13804 28754 13972 28756
rect 13804 28702 13806 28754
rect 13858 28702 13972 28754
rect 13804 28700 13972 28702
rect 14140 28980 14196 28990
rect 13804 28690 13860 28700
rect 14140 28642 14196 28924
rect 14140 28590 14142 28642
rect 14194 28590 14196 28642
rect 14140 28578 14196 28590
rect 13804 27860 13860 27870
rect 13804 27766 13860 27804
rect 14252 27746 14308 29372
rect 14476 29204 14532 29214
rect 14476 29110 14532 29148
rect 14364 29092 14420 29102
rect 14364 28644 14420 29036
rect 14588 28644 14644 30380
rect 14700 28756 14756 28766
rect 14700 28662 14756 28700
rect 14364 28550 14420 28588
rect 14476 28588 14644 28644
rect 14252 27694 14254 27746
rect 14306 27694 14308 27746
rect 14252 27682 14308 27694
rect 14028 27076 14084 27086
rect 14028 26962 14084 27020
rect 14028 26910 14030 26962
rect 14082 26910 14084 26962
rect 13692 26852 13860 26908
rect 14028 26898 14084 26910
rect 14476 26908 14532 28588
rect 14812 28532 14868 30604
rect 15036 30210 15092 31388
rect 15148 31218 15204 31612
rect 15148 31166 15150 31218
rect 15202 31166 15204 31218
rect 15148 31154 15204 31166
rect 15148 30436 15204 30446
rect 15260 30436 15316 31836
rect 15372 31220 15428 34190
rect 15820 34132 15876 34142
rect 15708 34076 15820 34132
rect 15708 33348 15764 34076
rect 15820 34038 15876 34076
rect 15708 33282 15764 33292
rect 15932 33124 15988 34860
rect 16044 33908 16100 34860
rect 16380 34692 16436 34702
rect 16716 34692 16772 34702
rect 16380 34690 16772 34692
rect 16380 34638 16382 34690
rect 16434 34638 16718 34690
rect 16770 34638 16772 34690
rect 16380 34636 16772 34638
rect 16380 34626 16436 34636
rect 16716 34626 16772 34636
rect 16828 34692 16884 34702
rect 16828 34598 16884 34636
rect 16940 34690 16996 34702
rect 16940 34638 16942 34690
rect 16994 34638 16996 34690
rect 16044 33842 16100 33852
rect 16268 34130 16324 34142
rect 16268 34078 16270 34130
rect 16322 34078 16324 34130
rect 16044 33348 16100 33358
rect 16044 33254 16100 33292
rect 15932 33058 15988 33068
rect 16268 33012 16324 34078
rect 16828 34018 16884 34030
rect 16828 33966 16830 34018
rect 16882 33966 16884 34018
rect 16828 33796 16884 33966
rect 16828 33730 16884 33740
rect 16940 33460 16996 34638
rect 16940 33394 16996 33404
rect 16044 32956 16324 33012
rect 16380 33348 16436 33358
rect 16044 32788 16100 32956
rect 15932 32732 16100 32788
rect 15596 32674 15652 32686
rect 15596 32622 15598 32674
rect 15650 32622 15652 32674
rect 15484 32562 15540 32574
rect 15484 32510 15486 32562
rect 15538 32510 15540 32562
rect 15484 32452 15540 32510
rect 15484 32386 15540 32396
rect 15596 31892 15652 32622
rect 15596 31826 15652 31836
rect 15932 31668 15988 32732
rect 16268 32674 16324 32686
rect 16268 32622 16270 32674
rect 16322 32622 16324 32674
rect 16044 32564 16100 32574
rect 16044 32470 16100 32508
rect 16268 32564 16324 32622
rect 16268 32498 16324 32508
rect 16156 32450 16212 32462
rect 16156 32398 16158 32450
rect 16210 32398 16212 32450
rect 15932 31612 16100 31668
rect 15372 31162 15428 31164
rect 15372 31110 15374 31162
rect 15426 31110 15428 31162
rect 15372 31098 15428 31110
rect 15484 31106 15540 31118
rect 15484 31054 15486 31106
rect 15538 31054 15540 31106
rect 15484 30996 15540 31054
rect 15708 31108 15764 31118
rect 15708 31014 15764 31052
rect 15148 30434 15316 30436
rect 15148 30382 15150 30434
rect 15202 30382 15316 30434
rect 15148 30380 15316 30382
rect 15372 30940 15540 30996
rect 16044 30996 16100 31612
rect 15148 30370 15204 30380
rect 15036 30158 15038 30210
rect 15090 30158 15092 30210
rect 15036 30146 15092 30158
rect 15372 30100 15428 30940
rect 16044 30930 16100 30940
rect 15932 30884 15988 30894
rect 15708 30882 15988 30884
rect 15708 30830 15934 30882
rect 15986 30830 15988 30882
rect 15708 30828 15988 30830
rect 15596 30100 15652 30110
rect 15372 30098 15652 30100
rect 15372 30046 15598 30098
rect 15650 30046 15652 30098
rect 15372 30044 15652 30046
rect 14700 28530 14868 28532
rect 14700 28478 14814 28530
rect 14866 28478 14868 28530
rect 14700 28476 14868 28478
rect 14588 28418 14644 28430
rect 14588 28366 14590 28418
rect 14642 28366 14644 28418
rect 14588 27860 14644 28366
rect 14588 27794 14644 27804
rect 14700 27970 14756 28476
rect 14812 28466 14868 28476
rect 15036 29538 15092 29550
rect 15036 29486 15038 29538
rect 15090 29486 15092 29538
rect 15036 28196 15092 29486
rect 15260 29428 15316 29438
rect 15260 29334 15316 29372
rect 14700 27918 14702 27970
rect 14754 27918 14756 27970
rect 14700 27748 14756 27918
rect 14700 27682 14756 27692
rect 14812 28140 15092 28196
rect 15260 28980 15316 28990
rect 14476 26852 14756 26908
rect 13692 26290 13748 26302
rect 13692 26238 13694 26290
rect 13746 26238 13748 26290
rect 13692 25284 13748 26238
rect 13804 26292 13860 26852
rect 14588 26516 14644 26526
rect 14588 26422 14644 26460
rect 13804 26226 13860 26236
rect 13916 26292 13972 26302
rect 13916 26290 14084 26292
rect 13916 26238 13918 26290
rect 13970 26238 14084 26290
rect 13916 26236 14084 26238
rect 13916 26226 13972 26236
rect 13804 25284 13860 25294
rect 13692 25282 13860 25284
rect 13692 25230 13806 25282
rect 13858 25230 13860 25282
rect 13692 25228 13860 25230
rect 13580 25218 13636 25228
rect 13356 24882 13412 24892
rect 13580 25060 13636 25070
rect 13132 24782 13134 24834
rect 13186 24782 13188 24834
rect 12460 24162 12628 24164
rect 12460 24110 12462 24162
rect 12514 24110 12628 24162
rect 12460 24108 12628 24110
rect 12460 24098 12516 24108
rect 13132 22596 13188 24782
rect 13468 24836 13524 24846
rect 13356 24724 13412 24734
rect 13356 24630 13412 24668
rect 13468 24722 13524 24780
rect 13468 24670 13470 24722
rect 13522 24670 13524 24722
rect 13468 23156 13524 24670
rect 13580 23938 13636 25004
rect 13692 24948 13748 24958
rect 13692 24164 13748 24892
rect 13804 24724 13860 25228
rect 14028 24836 14084 26236
rect 14700 25620 14756 26852
rect 14812 26516 14868 28140
rect 14924 27860 14980 27870
rect 14924 27766 14980 27804
rect 15148 27300 15204 27310
rect 15036 26964 15092 26974
rect 14924 26516 14980 26526
rect 14812 26514 14980 26516
rect 14812 26462 14926 26514
rect 14978 26462 14980 26514
rect 14812 26460 14980 26462
rect 14924 26450 14980 26460
rect 15036 26514 15092 26908
rect 15036 26462 15038 26514
rect 15090 26462 15092 26514
rect 15036 26450 15092 26462
rect 14812 26292 14868 26302
rect 14812 26198 14868 26236
rect 14700 25564 14980 25620
rect 14700 25394 14756 25406
rect 14700 25342 14702 25394
rect 14754 25342 14756 25394
rect 14476 25284 14532 25294
rect 14252 24836 14308 24846
rect 14028 24834 14252 24836
rect 14028 24782 14030 24834
rect 14082 24782 14252 24834
rect 14028 24780 14252 24782
rect 14028 24770 14084 24780
rect 13916 24724 13972 24734
rect 13804 24722 13972 24724
rect 13804 24670 13918 24722
rect 13970 24670 13972 24722
rect 13804 24668 13972 24670
rect 13692 24070 13748 24108
rect 13580 23886 13582 23938
rect 13634 23886 13636 23938
rect 13580 23874 13636 23886
rect 13916 23828 13972 24668
rect 14252 23938 14308 24780
rect 14252 23886 14254 23938
rect 14306 23886 14308 23938
rect 14252 23874 14308 23886
rect 14028 23828 14084 23838
rect 13916 23826 14084 23828
rect 13916 23774 14030 23826
rect 14082 23774 14084 23826
rect 13916 23772 14084 23774
rect 13356 23100 13524 23156
rect 13580 23492 13636 23502
rect 13916 23492 13972 23502
rect 13356 22708 13412 23100
rect 13468 22932 13524 22942
rect 13468 22838 13524 22876
rect 13580 22708 13636 23436
rect 13356 22652 13524 22708
rect 12012 22530 12068 22540
rect 12908 22540 13188 22596
rect 12460 22484 12516 22494
rect 12460 22482 12740 22484
rect 12460 22430 12462 22482
rect 12514 22430 12740 22482
rect 12460 22428 12740 22430
rect 12460 22418 12516 22428
rect 11564 22306 11620 22316
rect 11788 22372 11844 22382
rect 11788 22370 11956 22372
rect 11788 22318 11790 22370
rect 11842 22318 11956 22370
rect 11788 22316 11956 22318
rect 11788 22306 11844 22316
rect 11676 22260 11732 22270
rect 11676 22148 11732 22204
rect 11676 22092 11844 22148
rect 11116 21746 11172 21756
rect 11228 21980 11396 22036
rect 10668 21644 10836 21700
rect 10556 21364 10612 21374
rect 10556 21270 10612 21308
rect 10332 20972 10500 21028
rect 9884 19142 9940 19180
rect 10220 19170 10276 19180
rect 10332 20580 10388 20590
rect 10332 19234 10388 20524
rect 10332 19182 10334 19234
rect 10386 19182 10388 19234
rect 10332 19170 10388 19182
rect 10444 19012 10500 20972
rect 10668 20804 10724 21644
rect 11116 21588 11172 21598
rect 11116 21494 11172 21532
rect 10780 21476 10836 21486
rect 10780 21382 10836 21420
rect 10556 20748 10724 20804
rect 10556 20244 10612 20748
rect 10668 20580 10724 20590
rect 10668 20578 11172 20580
rect 10668 20526 10670 20578
rect 10722 20526 11172 20578
rect 10668 20524 11172 20526
rect 10668 20514 10724 20524
rect 10556 20188 10836 20244
rect 10668 20018 10724 20030
rect 10668 19966 10670 20018
rect 10722 19966 10724 20018
rect 10220 18956 10500 19012
rect 10556 19124 10612 19134
rect 9996 18450 10052 18462
rect 9996 18398 9998 18450
rect 10050 18398 10052 18450
rect 9772 18340 9828 18350
rect 9772 18246 9828 18284
rect 8876 17666 9716 17668
rect 8876 17614 9662 17666
rect 9714 17614 9716 17666
rect 8876 17612 9716 17614
rect 8876 17106 8932 17612
rect 9660 17602 9716 17612
rect 9884 17668 9940 17678
rect 9884 17574 9940 17612
rect 9436 17444 9492 17454
rect 8876 17054 8878 17106
rect 8930 17054 8932 17106
rect 8876 17042 8932 17054
rect 8988 17220 9044 17230
rect 8988 16884 9044 17164
rect 8876 16828 9044 16884
rect 8652 15698 8708 15708
rect 8764 16100 8820 16110
rect 7644 15092 8148 15148
rect 7308 13806 7310 13858
rect 7362 13806 7364 13858
rect 7308 13794 7364 13806
rect 7532 14532 7588 14542
rect 7084 13746 7140 13758
rect 7084 13694 7086 13746
rect 7138 13694 7140 13746
rect 7084 13636 7140 13694
rect 7532 13746 7588 14476
rect 7532 13694 7534 13746
rect 7586 13694 7588 13746
rect 7532 13682 7588 13694
rect 7868 13748 7924 13758
rect 7868 13746 8036 13748
rect 7868 13694 7870 13746
rect 7922 13694 8036 13746
rect 7868 13692 8036 13694
rect 7868 13682 7924 13692
rect 7084 13570 7140 13580
rect 7980 13522 8036 13692
rect 7980 13470 7982 13522
rect 8034 13470 8036 13522
rect 7980 13458 8036 13470
rect 7532 13186 7588 13198
rect 7532 13134 7534 13186
rect 7586 13134 7588 13186
rect 7532 12852 7588 13134
rect 7644 13076 7700 13086
rect 7644 13074 7812 13076
rect 7644 13022 7646 13074
rect 7698 13022 7812 13074
rect 7644 13020 7812 13022
rect 7644 13010 7700 13020
rect 7644 12852 7700 12862
rect 7532 12796 7644 12852
rect 7644 12786 7700 12796
rect 7084 12740 7140 12750
rect 6972 12684 7084 12740
rect 7084 12674 7140 12684
rect 7756 12068 7812 13020
rect 7980 12850 8036 12862
rect 7980 12798 7982 12850
rect 8034 12798 8036 12850
rect 7980 12740 8036 12798
rect 7868 12068 7924 12078
rect 6860 12066 7924 12068
rect 6860 12014 7870 12066
rect 7922 12014 7924 12066
rect 6860 12012 7924 12014
rect 6860 11618 6916 12012
rect 7868 12002 7924 12012
rect 6860 11566 6862 11618
rect 6914 11566 6916 11618
rect 6860 11554 6916 11566
rect 7308 11844 7364 11854
rect 6748 11340 7028 11396
rect 6524 11302 6580 11340
rect 6412 10770 6468 10780
rect 6636 11284 6692 11294
rect 5964 10670 5966 10722
rect 6018 10670 6020 10722
rect 5964 10658 6020 10670
rect 6636 10610 6692 11228
rect 6636 10558 6638 10610
rect 6690 10558 6692 10610
rect 6636 10500 6692 10558
rect 6860 10612 6916 10622
rect 6860 10518 6916 10556
rect 6636 10434 6692 10444
rect 5628 9998 5630 10050
rect 5682 9998 5684 10050
rect 5628 9986 5684 9998
rect 6300 10050 6356 10062
rect 6300 9998 6302 10050
rect 6354 9998 6356 10050
rect 6300 9938 6356 9998
rect 6300 9886 6302 9938
rect 6354 9886 6356 9938
rect 6300 9874 6356 9886
rect 5964 9828 6020 9838
rect 5404 9826 6020 9828
rect 5404 9774 5966 9826
rect 6018 9774 6020 9826
rect 5404 9772 6020 9774
rect 5964 9762 6020 9772
rect 6860 9604 6916 9614
rect 6972 9604 7028 11340
rect 7084 10500 7140 10510
rect 7308 10500 7364 11788
rect 7756 11844 7812 11854
rect 7420 11394 7476 11406
rect 7420 11342 7422 11394
rect 7474 11342 7476 11394
rect 7420 10724 7476 11342
rect 7756 11394 7812 11788
rect 7756 11342 7758 11394
rect 7810 11342 7812 11394
rect 7756 11172 7812 11342
rect 7756 11106 7812 11116
rect 7756 10836 7812 10846
rect 7756 10742 7812 10780
rect 7420 10722 7700 10724
rect 7420 10670 7422 10722
rect 7474 10670 7700 10722
rect 7420 10668 7700 10670
rect 7420 10658 7476 10668
rect 7308 10444 7588 10500
rect 7084 9826 7140 10444
rect 7084 9774 7086 9826
rect 7138 9774 7140 9826
rect 7084 9762 7140 9774
rect 7308 10164 7364 10174
rect 6860 9602 7028 9604
rect 6860 9550 6862 9602
rect 6914 9550 7028 9602
rect 6860 9548 7028 9550
rect 6860 9538 6916 9548
rect 6748 9268 6804 9278
rect 6748 9174 6804 9212
rect 7308 9042 7364 10108
rect 7532 9940 7588 10444
rect 7644 10388 7700 10668
rect 7980 10610 8036 12684
rect 7980 10558 7982 10610
rect 8034 10558 8036 10610
rect 7980 10546 8036 10558
rect 7980 10388 8036 10398
rect 7644 10386 8036 10388
rect 7644 10334 7982 10386
rect 8034 10334 8036 10386
rect 7644 10332 8036 10334
rect 7980 10322 8036 10332
rect 7532 9938 7700 9940
rect 7532 9886 7534 9938
rect 7586 9886 7700 9938
rect 7532 9884 7700 9886
rect 7532 9874 7588 9884
rect 7308 8990 7310 9042
rect 7362 8990 7364 9042
rect 7308 8978 7364 8990
rect 7084 8932 7140 8942
rect 7084 8838 7140 8876
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 7644 8260 7700 9884
rect 8092 9042 8148 15092
rect 8428 15092 8596 15148
rect 8204 13522 8260 13534
rect 8204 13470 8206 13522
rect 8258 13470 8260 13522
rect 8204 12178 8260 13470
rect 8428 13300 8484 15092
rect 8764 13972 8820 16044
rect 8876 15314 8932 16828
rect 8988 16100 9044 16110
rect 8988 16098 9156 16100
rect 8988 16046 8990 16098
rect 9042 16046 9156 16098
rect 8988 16044 9156 16046
rect 8988 16034 9044 16044
rect 8876 15262 8878 15314
rect 8930 15262 8932 15314
rect 8876 15250 8932 15262
rect 9100 14420 9156 16044
rect 9100 14354 9156 14364
rect 9324 15540 9380 15550
rect 9212 14308 9268 14318
rect 8876 13972 8932 13982
rect 8764 13970 8932 13972
rect 8764 13918 8878 13970
rect 8930 13918 8932 13970
rect 8764 13916 8932 13918
rect 8876 13906 8932 13916
rect 8540 13858 8596 13870
rect 8540 13806 8542 13858
rect 8594 13806 8596 13858
rect 8540 13412 8596 13806
rect 8764 13746 8820 13758
rect 8764 13694 8766 13746
rect 8818 13694 8820 13746
rect 8764 13524 8820 13694
rect 8988 13748 9044 13758
rect 8988 13654 9044 13692
rect 8764 13458 8820 13468
rect 8540 13346 8596 13356
rect 8428 13234 8484 13244
rect 8652 13076 8708 13086
rect 9212 13076 9268 14252
rect 8652 12962 8708 13020
rect 9100 13074 9268 13076
rect 9100 13022 9214 13074
rect 9266 13022 9268 13074
rect 9100 13020 9268 13022
rect 8652 12910 8654 12962
rect 8706 12910 8708 12962
rect 8652 12898 8708 12910
rect 8988 12962 9044 12974
rect 8988 12910 8990 12962
rect 9042 12910 9044 12962
rect 8204 12126 8206 12178
rect 8258 12126 8260 12178
rect 8204 11844 8260 12126
rect 8540 12852 8596 12862
rect 8540 12178 8596 12796
rect 8540 12126 8542 12178
rect 8594 12126 8596 12178
rect 8540 12114 8596 12126
rect 8988 12292 9044 12910
rect 8988 11956 9044 12236
rect 8988 11890 9044 11900
rect 8204 11778 8260 11788
rect 8428 11732 8484 11742
rect 8092 8990 8094 9042
rect 8146 8990 8148 9042
rect 8092 8978 8148 8990
rect 8204 11508 8260 11518
rect 7756 8820 7812 8830
rect 7756 8818 7924 8820
rect 7756 8766 7758 8818
rect 7810 8766 7924 8818
rect 7756 8764 7924 8766
rect 7756 8754 7812 8764
rect 7756 8260 7812 8270
rect 7644 8258 7812 8260
rect 7644 8206 7758 8258
rect 7810 8206 7812 8258
rect 7644 8204 7812 8206
rect 7756 8194 7812 8204
rect 7868 7812 7924 8764
rect 7980 8596 8036 8606
rect 7980 7924 8036 8540
rect 8204 8258 8260 11452
rect 8316 10836 8372 10846
rect 8316 10722 8372 10780
rect 8316 10670 8318 10722
rect 8370 10670 8372 10722
rect 8316 10658 8372 10670
rect 8316 9828 8372 9838
rect 8428 9828 8484 11676
rect 8876 11396 8932 11406
rect 8876 10834 8932 11340
rect 8876 10782 8878 10834
rect 8930 10782 8932 10834
rect 8876 10770 8932 10782
rect 8540 10724 8596 10734
rect 8540 10630 8596 10668
rect 8988 10612 9044 10622
rect 8988 10518 9044 10556
rect 9100 10052 9156 13020
rect 9212 13010 9268 13020
rect 9324 11732 9380 15484
rect 9436 15316 9492 17388
rect 9884 17220 9940 17230
rect 9548 16996 9604 17006
rect 9548 15764 9604 16940
rect 9884 16098 9940 17164
rect 9884 16046 9886 16098
rect 9938 16046 9940 16098
rect 9884 16034 9940 16046
rect 9996 16100 10052 18398
rect 10220 18452 10276 18956
rect 10332 18676 10388 18686
rect 10332 18582 10388 18620
rect 10556 18562 10612 19068
rect 10556 18510 10558 18562
rect 10610 18510 10612 18562
rect 10556 18498 10612 18510
rect 10220 18396 10388 18452
rect 10220 18228 10276 18238
rect 10108 17666 10164 17678
rect 10108 17614 10110 17666
rect 10162 17614 10164 17666
rect 10108 17108 10164 17614
rect 10108 17042 10164 17052
rect 10108 16882 10164 16894
rect 10108 16830 10110 16882
rect 10162 16830 10164 16882
rect 10108 16772 10164 16830
rect 10108 16706 10164 16716
rect 10220 16322 10276 18172
rect 10332 16772 10388 18396
rect 10332 16706 10388 16716
rect 10444 18338 10500 18350
rect 10444 18286 10446 18338
rect 10498 18286 10500 18338
rect 10220 16270 10222 16322
rect 10274 16270 10276 16322
rect 10220 16258 10276 16270
rect 10444 16324 10500 18286
rect 10668 17220 10724 19966
rect 10668 17154 10724 17164
rect 10780 17332 10836 20188
rect 11116 19124 11172 20524
rect 11228 20130 11284 21980
rect 11228 20078 11230 20130
rect 11282 20078 11284 20130
rect 11228 19460 11284 20078
rect 11228 19394 11284 19404
rect 11340 21810 11396 21822
rect 11340 21758 11342 21810
rect 11394 21758 11396 21810
rect 10780 16436 10836 17276
rect 11004 19122 11172 19124
rect 11004 19070 11118 19122
rect 11170 19070 11172 19122
rect 11004 19068 11172 19070
rect 11004 17892 11060 19068
rect 11116 19058 11172 19068
rect 11340 18788 11396 21758
rect 11788 21698 11844 22092
rect 11788 21646 11790 21698
rect 11842 21646 11844 21698
rect 11788 21634 11844 21646
rect 11900 20916 11956 22316
rect 12348 22260 12404 22298
rect 12348 22194 12404 22204
rect 12012 22148 12068 22158
rect 12012 22054 12068 22092
rect 12572 22148 12628 22158
rect 12572 22054 12628 22092
rect 12012 21812 12068 21822
rect 12012 21586 12068 21756
rect 12684 21700 12740 22428
rect 12684 21634 12740 21644
rect 12012 21534 12014 21586
rect 12066 21534 12068 21586
rect 12012 21522 12068 21534
rect 12572 21476 12628 21486
rect 12572 21382 12628 21420
rect 12012 21364 12068 21374
rect 12012 21026 12068 21308
rect 12012 20974 12014 21026
rect 12066 20974 12068 21026
rect 12012 20962 12068 20974
rect 12460 21364 12516 21374
rect 12460 21252 12516 21308
rect 12796 21362 12852 21374
rect 12796 21310 12798 21362
rect 12850 21310 12852 21362
rect 12796 21252 12852 21310
rect 12460 21196 12852 21252
rect 11900 20850 11956 20860
rect 12460 20914 12516 21196
rect 12460 20862 12462 20914
rect 12514 20862 12516 20914
rect 12460 20850 12516 20862
rect 12572 20916 12628 20926
rect 12572 20578 12628 20860
rect 12572 20526 12574 20578
rect 12626 20526 12628 20578
rect 11900 20244 11956 20254
rect 11788 20132 11844 20142
rect 11788 20038 11844 20076
rect 11788 19236 11844 19246
rect 11788 19142 11844 19180
rect 11452 19124 11508 19134
rect 11452 19122 11620 19124
rect 11452 19070 11454 19122
rect 11506 19070 11620 19122
rect 11452 19068 11620 19070
rect 11452 19058 11508 19068
rect 11004 17106 11060 17836
rect 11004 17054 11006 17106
rect 11058 17054 11060 17106
rect 11004 17042 11060 17054
rect 11116 18732 11396 18788
rect 10444 16258 10500 16268
rect 10556 16380 10836 16436
rect 11004 16884 11060 16894
rect 11116 16884 11172 18732
rect 11340 18562 11396 18574
rect 11340 18510 11342 18562
rect 11394 18510 11396 18562
rect 11340 18452 11396 18510
rect 11340 18386 11396 18396
rect 11340 18004 11396 18014
rect 11340 17778 11396 17948
rect 11340 17726 11342 17778
rect 11394 17726 11396 17778
rect 11340 17714 11396 17726
rect 11060 16828 11172 16884
rect 9996 16034 10052 16044
rect 9660 15988 9716 15998
rect 9660 15986 9828 15988
rect 9660 15934 9662 15986
rect 9714 15934 9828 15986
rect 9660 15932 9828 15934
rect 9660 15922 9716 15932
rect 9548 15708 9716 15764
rect 9660 15426 9716 15708
rect 9660 15374 9662 15426
rect 9714 15374 9716 15426
rect 9660 15362 9716 15374
rect 9548 15316 9604 15326
rect 9436 15314 9604 15316
rect 9436 15262 9550 15314
rect 9602 15262 9604 15314
rect 9436 15260 9604 15262
rect 9548 15250 9604 15260
rect 9772 15148 9828 15932
rect 9548 15092 9828 15148
rect 10108 15202 10164 15214
rect 10108 15150 10110 15202
rect 10162 15150 10164 15202
rect 9324 11666 9380 11676
rect 9436 14530 9492 14542
rect 9436 14478 9438 14530
rect 9490 14478 9492 14530
rect 9436 13636 9492 14478
rect 9436 11508 9492 13580
rect 9548 13412 9604 15092
rect 9884 14420 9940 14430
rect 9884 14326 9940 14364
rect 9660 14308 9716 14318
rect 9660 13746 9716 14252
rect 9660 13694 9662 13746
rect 9714 13694 9716 13746
rect 9660 13682 9716 13694
rect 9996 13746 10052 13758
rect 9996 13694 9998 13746
rect 10050 13694 10052 13746
rect 9548 13346 9604 13356
rect 9884 13074 9940 13086
rect 9884 13022 9886 13074
rect 9938 13022 9940 13074
rect 9884 12852 9940 13022
rect 9884 12786 9940 12796
rect 9996 13076 10052 13694
rect 9660 12740 9716 12750
rect 9660 12738 9828 12740
rect 9660 12686 9662 12738
rect 9714 12686 9828 12738
rect 9660 12684 9828 12686
rect 9660 12674 9716 12684
rect 8316 9826 8484 9828
rect 8316 9774 8318 9826
rect 8370 9774 8484 9826
rect 8316 9772 8484 9774
rect 8764 9996 9156 10052
rect 9324 11452 9492 11508
rect 9548 12178 9604 12190
rect 9548 12126 9550 12178
rect 9602 12126 9604 12178
rect 8316 9762 8372 9772
rect 8316 9604 8372 9614
rect 8652 9604 8708 9614
rect 8316 8370 8372 9548
rect 8540 9602 8708 9604
rect 8540 9550 8654 9602
rect 8706 9550 8708 9602
rect 8540 9548 8708 9550
rect 8540 8596 8596 9548
rect 8652 9538 8708 9548
rect 8764 9268 8820 9996
rect 8540 8530 8596 8540
rect 8652 9212 8820 9268
rect 8988 9826 9044 9838
rect 8988 9774 8990 9826
rect 9042 9774 9044 9826
rect 8316 8318 8318 8370
rect 8370 8318 8372 8370
rect 8316 8306 8372 8318
rect 8652 8260 8708 9212
rect 8876 9156 8932 9166
rect 8876 9062 8932 9100
rect 8764 9044 8820 9054
rect 8764 8950 8820 8988
rect 8988 8372 9044 9774
rect 9324 9716 9380 11452
rect 9324 9650 9380 9660
rect 9436 10836 9492 10846
rect 9436 9380 9492 10780
rect 9548 9604 9604 12126
rect 9660 10612 9716 10622
rect 9660 9714 9716 10556
rect 9772 10612 9828 12684
rect 9996 12404 10052 13020
rect 9884 12348 10052 12404
rect 9884 11508 9940 12348
rect 10108 12292 10164 15150
rect 10556 15148 10612 16380
rect 10332 15092 10612 15148
rect 10668 16210 10724 16222
rect 10668 16158 10670 16210
rect 10722 16158 10724 16210
rect 9996 12236 10164 12292
rect 10220 13972 10276 13982
rect 9996 11844 10052 12236
rect 10220 12178 10276 13916
rect 10332 12290 10388 15092
rect 10668 13748 10724 16158
rect 10780 15314 10836 15326
rect 10780 15262 10782 15314
rect 10834 15262 10836 15314
rect 10780 15148 10836 15262
rect 11004 15314 11060 16828
rect 11116 16100 11172 16110
rect 11116 16098 11284 16100
rect 11116 16046 11118 16098
rect 11170 16046 11284 16098
rect 11116 16044 11284 16046
rect 11116 16034 11172 16044
rect 11004 15262 11006 15314
rect 11058 15262 11060 15314
rect 11004 15250 11060 15262
rect 10780 15092 10948 15148
rect 10332 12238 10334 12290
rect 10386 12238 10388 12290
rect 10332 12226 10388 12238
rect 10444 13524 10500 13534
rect 10220 12126 10222 12178
rect 10274 12126 10276 12178
rect 10108 12068 10164 12078
rect 10108 11974 10164 12012
rect 9996 11788 10164 11844
rect 10108 11620 10164 11788
rect 10108 11554 10164 11564
rect 9884 11414 9940 11452
rect 10220 10836 10276 12126
rect 10444 12068 10500 13468
rect 10220 10770 10276 10780
rect 10332 12012 10500 12068
rect 10556 12292 10612 12302
rect 9772 10610 10052 10612
rect 9772 10558 9774 10610
rect 9826 10558 10052 10610
rect 9772 10556 10052 10558
rect 9772 10546 9828 10556
rect 9772 10388 9828 10398
rect 9772 9826 9828 10332
rect 9996 10164 10052 10556
rect 10220 10610 10276 10622
rect 10220 10558 10222 10610
rect 10274 10558 10276 10610
rect 10220 10388 10276 10558
rect 10220 10322 10276 10332
rect 9996 10108 10164 10164
rect 9772 9774 9774 9826
rect 9826 9774 9828 9826
rect 9772 9762 9828 9774
rect 9996 9940 10052 9950
rect 9660 9662 9662 9714
rect 9714 9662 9716 9714
rect 9660 9650 9716 9662
rect 9884 9716 9940 9726
rect 9548 9538 9604 9548
rect 9436 9324 9828 9380
rect 8988 8316 9716 8372
rect 8204 8206 8206 8258
rect 8258 8206 8260 8258
rect 8204 8194 8260 8206
rect 8428 8204 8708 8260
rect 8428 8146 8484 8204
rect 9100 8148 9156 8158
rect 8428 8094 8430 8146
rect 8482 8094 8484 8146
rect 8428 8082 8484 8094
rect 8540 8146 9156 8148
rect 8540 8094 9102 8146
rect 9154 8094 9156 8146
rect 8540 8092 9156 8094
rect 7980 7868 8372 7924
rect 7868 7756 8260 7812
rect 8204 7586 8260 7756
rect 8316 7698 8372 7868
rect 8316 7646 8318 7698
rect 8370 7646 8372 7698
rect 8316 7634 8372 7646
rect 8540 7698 8596 8092
rect 9100 8082 9156 8092
rect 9548 8148 9604 8158
rect 8540 7646 8542 7698
rect 8594 7646 8596 7698
rect 8540 7634 8596 7646
rect 8204 7534 8206 7586
rect 8258 7534 8260 7586
rect 8204 7522 8260 7534
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 9548 6690 9604 8092
rect 9548 6638 9550 6690
rect 9602 6638 9604 6690
rect 9548 6626 9604 6638
rect 9660 6690 9716 8316
rect 9660 6638 9662 6690
rect 9714 6638 9716 6690
rect 9660 6626 9716 6638
rect 9772 6690 9828 9324
rect 9884 7700 9940 9660
rect 9996 9266 10052 9884
rect 9996 9214 9998 9266
rect 10050 9214 10052 9266
rect 9996 9202 10052 9214
rect 9996 7700 10052 7710
rect 9884 7698 10052 7700
rect 9884 7646 9998 7698
rect 10050 7646 10052 7698
rect 9884 7644 10052 7646
rect 9996 7634 10052 7644
rect 9772 6638 9774 6690
rect 9826 6638 9828 6690
rect 9772 6626 9828 6638
rect 10108 6690 10164 10108
rect 10220 9828 10276 9838
rect 10332 9828 10388 12012
rect 10556 11396 10612 12236
rect 10444 11340 10612 11396
rect 10444 11282 10500 11340
rect 10444 11230 10446 11282
rect 10498 11230 10500 11282
rect 10444 11218 10500 11230
rect 10220 9826 10388 9828
rect 10220 9774 10222 9826
rect 10274 9774 10388 9826
rect 10220 9772 10388 9774
rect 10220 9044 10276 9772
rect 10220 8978 10276 8988
rect 10556 9716 10612 9726
rect 10668 9716 10724 13692
rect 10892 14642 10948 15092
rect 10892 14590 10894 14642
rect 10946 14590 10948 14642
rect 10892 13636 10948 14590
rect 11228 14530 11284 16044
rect 11452 15316 11508 15326
rect 11452 15222 11508 15260
rect 11228 14478 11230 14530
rect 11282 14478 11284 14530
rect 11228 14420 11284 14478
rect 11564 14532 11620 19068
rect 11900 19010 11956 20188
rect 12572 20132 12628 20526
rect 12012 20020 12068 20030
rect 12012 19926 12068 19964
rect 12236 19906 12292 19918
rect 12236 19854 12238 19906
rect 12290 19854 12292 19906
rect 11900 18958 11902 19010
rect 11954 18958 11956 19010
rect 11900 18946 11956 18958
rect 12124 19124 12180 19134
rect 11900 18564 11956 18574
rect 11676 17444 11732 17454
rect 11676 17350 11732 17388
rect 11900 15652 11956 18508
rect 12012 17892 12068 17902
rect 12012 17798 12068 17836
rect 11900 15586 11956 15596
rect 12012 16548 12068 16558
rect 11788 15540 11844 15550
rect 11788 15314 11844 15484
rect 12012 15428 12068 16492
rect 12124 16322 12180 19068
rect 12124 16270 12126 16322
rect 12178 16270 12180 16322
rect 12124 16258 12180 16270
rect 12236 18676 12292 19854
rect 12348 19908 12404 19918
rect 12348 19814 12404 19852
rect 12348 19236 12404 19246
rect 12348 19142 12404 19180
rect 12572 19122 12628 20076
rect 12684 20018 12740 21196
rect 12684 19966 12686 20018
rect 12738 19966 12740 20018
rect 12684 19954 12740 19966
rect 12572 19070 12574 19122
rect 12626 19070 12628 19122
rect 12572 19058 12628 19070
rect 12236 16324 12292 18620
rect 12684 18564 12740 18574
rect 12908 18564 12964 22540
rect 13020 22372 13076 22382
rect 13020 22370 13188 22372
rect 13020 22318 13022 22370
rect 13074 22318 13188 22370
rect 13020 22316 13188 22318
rect 13020 22306 13076 22316
rect 13020 21476 13076 21486
rect 13020 19348 13076 21420
rect 13132 21362 13188 22316
rect 13132 21310 13134 21362
rect 13186 21310 13188 21362
rect 13132 20020 13188 21310
rect 13468 20356 13524 22652
rect 13580 22482 13636 22652
rect 13580 22430 13582 22482
rect 13634 22430 13636 22482
rect 13580 22418 13636 22430
rect 13692 23436 13916 23492
rect 14028 23492 14084 23772
rect 14140 23716 14196 23726
rect 14140 23622 14196 23660
rect 14028 23436 14196 23492
rect 13580 21588 13636 21598
rect 13692 21588 13748 23436
rect 13916 23426 13972 23436
rect 14028 23268 14084 23278
rect 14140 23268 14196 23436
rect 14140 23212 14420 23268
rect 13916 23156 13972 23166
rect 13916 22372 13972 23100
rect 14028 22482 14084 23212
rect 14364 23154 14420 23212
rect 14364 23102 14366 23154
rect 14418 23102 14420 23154
rect 14364 23090 14420 23102
rect 14028 22430 14030 22482
rect 14082 22430 14084 22482
rect 14028 22418 14084 22430
rect 14140 22932 14196 22942
rect 13580 21586 13748 21588
rect 13580 21534 13582 21586
rect 13634 21534 13748 21586
rect 13580 21532 13748 21534
rect 13580 21522 13636 21532
rect 13692 20804 13748 21532
rect 13692 20738 13748 20748
rect 13804 22370 13972 22372
rect 13804 22318 13918 22370
rect 13970 22318 13972 22370
rect 13804 22316 13972 22318
rect 13804 21586 13860 22316
rect 13916 22306 13972 22316
rect 14140 22370 14196 22876
rect 14476 22596 14532 25228
rect 14700 24948 14756 25342
rect 14700 24882 14756 24892
rect 14700 24500 14756 24510
rect 14588 24498 14756 24500
rect 14588 24446 14702 24498
rect 14754 24446 14756 24498
rect 14588 24444 14756 24446
rect 14588 23268 14644 24444
rect 14700 24434 14756 24444
rect 14700 24164 14756 24174
rect 14700 23268 14756 24108
rect 14812 23714 14868 23726
rect 14812 23662 14814 23714
rect 14866 23662 14868 23714
rect 14812 23492 14868 23662
rect 14812 23426 14868 23436
rect 14812 23268 14868 23278
rect 14700 23266 14868 23268
rect 14700 23214 14814 23266
rect 14866 23214 14868 23266
rect 14700 23212 14868 23214
rect 14588 23202 14644 23212
rect 14812 23202 14868 23212
rect 14700 23044 14756 23054
rect 14476 22530 14532 22540
rect 14588 23042 14756 23044
rect 14588 22990 14702 23042
rect 14754 22990 14756 23042
rect 14588 22988 14756 22990
rect 14588 22484 14644 22988
rect 14700 22978 14756 22988
rect 14924 22820 14980 25564
rect 15148 25508 15204 27244
rect 15148 25442 15204 25452
rect 15260 26180 15316 28924
rect 15596 28866 15652 30044
rect 15708 29538 15764 30828
rect 15932 30818 15988 30828
rect 15820 29652 15876 29662
rect 16156 29652 16212 32398
rect 16380 32452 16436 33292
rect 16828 33346 16884 33358
rect 16828 33294 16830 33346
rect 16882 33294 16884 33346
rect 16492 32676 16548 32686
rect 16492 32562 16548 32620
rect 16492 32510 16494 32562
rect 16546 32510 16548 32562
rect 16492 32498 16548 32510
rect 16604 32674 16660 32686
rect 16604 32622 16606 32674
rect 16658 32622 16660 32674
rect 16380 32386 16436 32396
rect 16268 31892 16324 31902
rect 16324 31836 16436 31892
rect 16268 31826 16324 31836
rect 16268 31220 16324 31230
rect 16268 31126 16324 31164
rect 16380 31218 16436 31836
rect 16492 31780 16548 31790
rect 16604 31780 16660 32622
rect 16828 31948 16884 33294
rect 16492 31778 16660 31780
rect 16492 31726 16494 31778
rect 16546 31726 16660 31778
rect 16492 31724 16660 31726
rect 16716 31892 16884 31948
rect 16492 31444 16548 31724
rect 16492 31378 16548 31388
rect 16604 31556 16660 31566
rect 16380 31166 16382 31218
rect 16434 31166 16436 31218
rect 16380 31154 16436 31166
rect 16492 30996 16548 31006
rect 16492 30902 16548 30940
rect 16604 30884 16660 31500
rect 16716 31108 16772 31892
rect 16828 31780 16884 31790
rect 16828 31686 16884 31724
rect 16716 31042 16772 31052
rect 16940 31444 16996 31454
rect 16940 30994 16996 31388
rect 16940 30942 16942 30994
rect 16994 30942 16996 30994
rect 16940 30930 16996 30942
rect 16604 30828 16772 30884
rect 16716 30322 16772 30828
rect 16716 30270 16718 30322
rect 16770 30270 16772 30322
rect 16604 30210 16660 30222
rect 16604 30158 16606 30210
rect 16658 30158 16660 30210
rect 15820 29650 16212 29652
rect 15820 29598 15822 29650
rect 15874 29598 16212 29650
rect 15820 29596 16212 29598
rect 16380 30100 16436 30110
rect 16380 29650 16436 30044
rect 16380 29598 16382 29650
rect 16434 29598 16436 29650
rect 15820 29586 15876 29596
rect 16380 29586 16436 29598
rect 15708 29486 15710 29538
rect 15762 29486 15764 29538
rect 15708 29474 15764 29486
rect 16492 29540 16548 29550
rect 16492 29446 16548 29484
rect 16044 29428 16100 29438
rect 16268 29428 16324 29438
rect 16044 29426 16324 29428
rect 16044 29374 16046 29426
rect 16098 29374 16270 29426
rect 16322 29374 16324 29426
rect 16044 29372 16324 29374
rect 16044 29362 16100 29372
rect 16268 29362 16324 29372
rect 16604 29428 16660 30158
rect 16604 29204 16660 29372
rect 16380 29148 16660 29204
rect 16716 29204 16772 30270
rect 16940 29652 16996 29662
rect 16940 29426 16996 29596
rect 16940 29374 16942 29426
rect 16994 29374 16996 29426
rect 16940 29362 16996 29374
rect 15596 28814 15598 28866
rect 15650 28814 15652 28866
rect 15596 28802 15652 28814
rect 16156 29092 16212 29102
rect 15820 28530 15876 28542
rect 15820 28478 15822 28530
rect 15874 28478 15876 28530
rect 15484 26962 15540 26974
rect 15484 26910 15486 26962
rect 15538 26910 15540 26962
rect 15484 26852 15540 26910
rect 15484 26786 15540 26796
rect 15484 26628 15540 26638
rect 15372 26180 15428 26190
rect 15260 26178 15428 26180
rect 15260 26126 15374 26178
rect 15426 26126 15428 26178
rect 15260 26124 15428 26126
rect 15036 25060 15092 25070
rect 15036 24946 15092 25004
rect 15036 24894 15038 24946
rect 15090 24894 15092 24946
rect 15036 24882 15092 24894
rect 14924 22754 14980 22764
rect 15036 23938 15092 23950
rect 15036 23886 15038 23938
rect 15090 23886 15092 23938
rect 15036 22596 15092 23886
rect 15148 23156 15204 23166
rect 15148 23062 15204 23100
rect 15036 22530 15092 22540
rect 14924 22484 14980 22494
rect 14588 22482 14980 22484
rect 14588 22430 14926 22482
rect 14978 22430 14980 22482
rect 14588 22428 14980 22430
rect 14140 22318 14142 22370
rect 14194 22318 14196 22370
rect 14140 22306 14196 22318
rect 14476 22372 14532 22382
rect 14588 22372 14644 22428
rect 14924 22418 14980 22428
rect 14476 22370 14644 22372
rect 14476 22318 14478 22370
rect 14530 22318 14644 22370
rect 14476 22316 14644 22318
rect 15036 22370 15092 22382
rect 15036 22318 15038 22370
rect 15090 22318 15092 22370
rect 14476 22306 14532 22316
rect 14812 22258 14868 22270
rect 14812 22206 14814 22258
rect 14866 22206 14868 22258
rect 13804 21534 13806 21586
rect 13858 21534 13860 21586
rect 13468 20300 13748 20356
rect 13132 19954 13188 19964
rect 13468 20018 13524 20030
rect 13468 19966 13470 20018
rect 13522 19966 13524 20018
rect 13468 19796 13524 19966
rect 13468 19730 13524 19740
rect 13692 19572 13748 20300
rect 13692 19506 13748 19516
rect 13804 19460 13860 21534
rect 13804 19394 13860 19404
rect 13916 22148 13972 22158
rect 13020 19292 13300 19348
rect 13020 19012 13076 19022
rect 13020 18676 13076 18956
rect 13020 18610 13076 18620
rect 12740 18508 12964 18564
rect 12684 18498 12740 18508
rect 13132 18226 13188 18238
rect 13132 18174 13134 18226
rect 13186 18174 13188 18226
rect 13132 17780 13188 18174
rect 12684 17666 12740 17678
rect 12684 17614 12686 17666
rect 12738 17614 12740 17666
rect 12684 16884 12740 17614
rect 12796 17556 12852 17566
rect 13132 17556 13188 17724
rect 12796 17554 13188 17556
rect 12796 17502 12798 17554
rect 12850 17502 13188 17554
rect 12796 17500 13188 17502
rect 12796 17490 12852 17500
rect 13132 17108 13188 17118
rect 13020 17052 13132 17108
rect 12908 16884 12964 16894
rect 12684 16828 12908 16884
rect 12908 16790 12964 16828
rect 12908 16660 12964 16670
rect 12348 16324 12404 16334
rect 12908 16324 12964 16604
rect 12236 16322 12404 16324
rect 12236 16270 12350 16322
rect 12402 16270 12404 16322
rect 12236 16268 12404 16270
rect 12348 16258 12404 16268
rect 12796 16322 12964 16324
rect 12796 16270 12910 16322
rect 12962 16270 12964 16322
rect 12796 16268 12964 16270
rect 12684 16100 12740 16110
rect 12684 16006 12740 16044
rect 12572 15986 12628 15998
rect 12572 15934 12574 15986
rect 12626 15934 12628 15986
rect 12012 15426 12180 15428
rect 12012 15374 12014 15426
rect 12066 15374 12180 15426
rect 12012 15372 12180 15374
rect 12012 15362 12068 15372
rect 11788 15262 11790 15314
rect 11842 15262 11844 15314
rect 11788 15250 11844 15262
rect 11900 15202 11956 15214
rect 11900 15150 11902 15202
rect 11954 15150 11956 15202
rect 11564 14466 11620 14476
rect 11788 14530 11844 14542
rect 11788 14478 11790 14530
rect 11842 14478 11844 14530
rect 11228 14354 11284 14364
rect 11564 14084 11620 14094
rect 11004 13860 11060 13870
rect 11004 13746 11060 13804
rect 11004 13694 11006 13746
rect 11058 13694 11060 13746
rect 11004 13636 11060 13694
rect 11564 13746 11620 14028
rect 11564 13694 11566 13746
rect 11618 13694 11620 13746
rect 11564 13682 11620 13694
rect 11676 13748 11732 13758
rect 11116 13636 11172 13646
rect 11004 13580 11116 13636
rect 10892 13570 10948 13580
rect 11116 13570 11172 13580
rect 10780 13524 10836 13534
rect 10780 13430 10836 13468
rect 11228 13412 11284 13422
rect 11228 12402 11284 13356
rect 11228 12350 11230 12402
rect 11282 12350 11284 12402
rect 11228 12338 11284 12350
rect 10892 12068 10948 12078
rect 10780 11394 10836 11406
rect 10780 11342 10782 11394
rect 10834 11342 10836 11394
rect 10780 10724 10836 11342
rect 10780 10658 10836 10668
rect 10556 9714 10724 9716
rect 10556 9662 10558 9714
rect 10610 9662 10724 9714
rect 10556 9660 10724 9662
rect 10892 10610 10948 12012
rect 11564 11956 11620 11966
rect 11676 11956 11732 13692
rect 11788 12292 11844 14478
rect 11900 13076 11956 15150
rect 12012 13076 12068 13086
rect 11900 13074 12068 13076
rect 11900 13022 12014 13074
rect 12066 13022 12068 13074
rect 11900 13020 12068 13022
rect 12012 13010 12068 13020
rect 11788 12226 11844 12236
rect 11900 12180 11956 12190
rect 11564 11954 11732 11956
rect 11564 11902 11566 11954
rect 11618 11902 11732 11954
rect 11564 11900 11732 11902
rect 11788 12066 11844 12078
rect 11788 12014 11790 12066
rect 11842 12014 11844 12066
rect 11004 10836 11060 10846
rect 11004 10722 11060 10780
rect 11004 10670 11006 10722
rect 11058 10670 11060 10722
rect 11004 10658 11060 10670
rect 10892 10558 10894 10610
rect 10946 10558 10948 10610
rect 10444 8932 10500 8942
rect 10444 8838 10500 8876
rect 10556 6914 10612 9660
rect 10892 8148 10948 10558
rect 11228 10500 11284 10510
rect 11228 10406 11284 10444
rect 11564 10052 11620 11900
rect 11788 11732 11844 12014
rect 11676 11676 11844 11732
rect 11676 11284 11732 11676
rect 11788 11508 11844 11518
rect 11900 11508 11956 12124
rect 12124 11788 12180 15372
rect 12572 15314 12628 15934
rect 12572 15262 12574 15314
rect 12626 15262 12628 15314
rect 12572 15250 12628 15262
rect 12236 14530 12292 14542
rect 12236 14478 12238 14530
rect 12290 14478 12292 14530
rect 12236 13972 12292 14478
rect 12572 14420 12628 14430
rect 12572 14326 12628 14364
rect 12684 14418 12740 14430
rect 12684 14366 12686 14418
rect 12738 14366 12740 14418
rect 12236 13906 12292 13916
rect 12572 14084 12628 14094
rect 12460 13860 12516 13870
rect 12348 13804 12460 13860
rect 12348 13746 12404 13804
rect 12460 13794 12516 13804
rect 12348 13694 12350 13746
rect 12402 13694 12404 13746
rect 12348 13682 12404 13694
rect 12572 12964 12628 14028
rect 12684 13748 12740 14366
rect 12684 13682 12740 13692
rect 12684 12964 12740 12974
rect 12572 12962 12740 12964
rect 12572 12910 12686 12962
rect 12738 12910 12740 12962
rect 12572 12908 12740 12910
rect 12460 12180 12516 12190
rect 12348 12124 12460 12180
rect 12348 11844 12404 12124
rect 12460 12086 12516 12124
rect 12348 11788 12516 11844
rect 11788 11506 11956 11508
rect 11788 11454 11790 11506
rect 11842 11454 11956 11506
rect 11788 11452 11956 11454
rect 12012 11732 12180 11788
rect 11788 11442 11844 11452
rect 11676 11228 11844 11284
rect 11676 11060 11732 11070
rect 11676 10612 11732 11004
rect 11676 10518 11732 10556
rect 11788 10164 11844 11228
rect 11900 10610 11956 10622
rect 11900 10558 11902 10610
rect 11954 10558 11956 10610
rect 11900 10388 11956 10558
rect 11900 10322 11956 10332
rect 11788 10098 11844 10108
rect 12012 10052 12068 11732
rect 12124 11620 12180 11630
rect 12348 11620 12404 11630
rect 12124 10276 12180 11564
rect 12236 11564 12348 11620
rect 12236 10500 12292 11564
rect 12348 11554 12404 11564
rect 12348 11396 12404 11406
rect 12348 11302 12404 11340
rect 12460 11284 12516 11788
rect 12572 11508 12628 12908
rect 12684 12898 12740 12908
rect 12684 11954 12740 11966
rect 12684 11902 12686 11954
rect 12738 11902 12740 11954
rect 12684 11620 12740 11902
rect 12796 11788 12852 16268
rect 12908 16258 12964 16268
rect 13020 16100 13076 17052
rect 13132 17042 13188 17052
rect 12908 16044 13076 16100
rect 13132 16436 13188 16446
rect 12908 15314 12964 16044
rect 13020 15540 13076 15550
rect 13132 15540 13188 16380
rect 13244 16212 13300 19292
rect 13916 19236 13972 22092
rect 14476 21588 14532 21598
rect 14364 21586 14532 21588
rect 14364 21534 14478 21586
rect 14530 21534 14532 21586
rect 14364 21532 14532 21534
rect 14140 21476 14196 21486
rect 14364 21476 14420 21532
rect 14476 21522 14532 21532
rect 14700 21586 14756 21598
rect 14700 21534 14702 21586
rect 14754 21534 14756 21586
rect 14140 21474 14420 21476
rect 14140 21422 14142 21474
rect 14194 21422 14420 21474
rect 14140 21420 14420 21422
rect 14588 21474 14644 21486
rect 14588 21422 14590 21474
rect 14642 21422 14644 21474
rect 14140 21410 14196 21420
rect 14028 21364 14084 21374
rect 14028 20916 14084 21308
rect 14588 21252 14644 21422
rect 14700 21364 14756 21534
rect 14700 21298 14756 21308
rect 14364 21196 14644 21252
rect 14028 20914 14196 20916
rect 14028 20862 14030 20914
rect 14082 20862 14196 20914
rect 14028 20860 14196 20862
rect 14028 20850 14084 20860
rect 14140 19346 14196 20860
rect 14140 19294 14142 19346
rect 14194 19294 14196 19346
rect 14140 19282 14196 19294
rect 13580 19234 13972 19236
rect 13580 19182 13918 19234
rect 13970 19182 13972 19234
rect 13580 19180 13972 19182
rect 13356 18676 13412 18714
rect 13356 18610 13412 18620
rect 13580 18674 13636 19180
rect 13916 19170 13972 19180
rect 14252 19124 14308 19134
rect 14252 19030 14308 19068
rect 13580 18622 13582 18674
rect 13634 18622 13636 18674
rect 13580 18610 13636 18622
rect 13916 18562 13972 18574
rect 13916 18510 13918 18562
rect 13970 18510 13972 18562
rect 13468 18452 13524 18462
rect 13468 18358 13524 18396
rect 13804 18452 13860 18462
rect 13804 18358 13860 18396
rect 13580 17892 13636 17902
rect 13580 17554 13636 17836
rect 13580 17502 13582 17554
rect 13634 17502 13636 17554
rect 13580 17490 13636 17502
rect 13916 17106 13972 18510
rect 14364 18452 14420 21196
rect 14812 21028 14868 22206
rect 14924 22148 14980 22158
rect 14924 21810 14980 22092
rect 14924 21758 14926 21810
rect 14978 21758 14980 21810
rect 14924 21746 14980 21758
rect 15036 21028 15092 22318
rect 15260 22260 15316 26124
rect 15372 26114 15428 26124
rect 15484 25844 15540 26572
rect 15820 26516 15876 28478
rect 15820 26450 15876 26460
rect 15932 27858 15988 27870
rect 15932 27806 15934 27858
rect 15986 27806 15988 27858
rect 15932 26852 15988 27806
rect 15820 26292 15876 26302
rect 15820 26198 15876 26236
rect 15484 25778 15540 25788
rect 15596 26180 15652 26190
rect 15596 24610 15652 26124
rect 15820 24724 15876 24734
rect 15932 24724 15988 26796
rect 16044 27746 16100 27758
rect 16044 27694 16046 27746
rect 16098 27694 16100 27746
rect 16044 25620 16100 27694
rect 16156 27748 16212 29036
rect 16268 28644 16324 28654
rect 16268 27970 16324 28588
rect 16380 28642 16436 29148
rect 16716 29138 16772 29148
rect 17052 28868 17108 35420
rect 17052 28802 17108 28812
rect 17164 35364 17220 35374
rect 16380 28590 16382 28642
rect 16434 28590 16436 28642
rect 16380 28578 16436 28590
rect 16940 28642 16996 28654
rect 16940 28590 16942 28642
rect 16994 28590 16996 28642
rect 16268 27918 16270 27970
rect 16322 27918 16324 27970
rect 16268 27906 16324 27918
rect 16604 28420 16660 28430
rect 16156 27692 16324 27748
rect 16044 25554 16100 25564
rect 16156 27074 16212 27086
rect 16156 27022 16158 27074
rect 16210 27022 16212 27074
rect 16156 24946 16212 27022
rect 16268 26292 16324 27692
rect 16268 26290 16436 26292
rect 16268 26238 16270 26290
rect 16322 26238 16436 26290
rect 16268 26236 16436 26238
rect 16268 26226 16324 26236
rect 16380 25732 16436 26236
rect 16492 26068 16548 26078
rect 16492 25974 16548 26012
rect 16492 25732 16548 25742
rect 16380 25730 16548 25732
rect 16380 25678 16494 25730
rect 16546 25678 16548 25730
rect 16380 25676 16548 25678
rect 16492 25666 16548 25676
rect 16604 25172 16660 28364
rect 16716 27748 16772 27758
rect 16716 27654 16772 27692
rect 16828 27634 16884 27646
rect 16828 27582 16830 27634
rect 16882 27582 16884 27634
rect 16828 26740 16884 27582
rect 16940 27074 16996 28590
rect 17164 28420 17220 35308
rect 17388 35140 17444 35646
rect 17612 35698 17668 36092
rect 17612 35646 17614 35698
rect 17666 35646 17668 35698
rect 17612 35364 17668 35646
rect 17612 35298 17668 35308
rect 17836 35140 17892 36540
rect 18284 36530 18340 36540
rect 18396 36482 18452 36494
rect 18396 36430 18398 36482
rect 18450 36430 18452 36482
rect 17948 36370 18004 36382
rect 17948 36318 17950 36370
rect 18002 36318 18004 36370
rect 17948 35700 18004 36318
rect 18284 36260 18340 36270
rect 18284 35922 18340 36204
rect 18396 36148 18452 36430
rect 18396 36082 18452 36092
rect 18508 36372 18564 36382
rect 18284 35870 18286 35922
rect 18338 35870 18340 35922
rect 18284 35858 18340 35870
rect 18396 35924 18452 35934
rect 18508 35924 18564 36316
rect 18396 35922 18564 35924
rect 18396 35870 18398 35922
rect 18450 35870 18564 35922
rect 18396 35868 18564 35870
rect 18396 35858 18452 35868
rect 18060 35700 18116 35710
rect 17948 35698 18116 35700
rect 17948 35646 18062 35698
rect 18114 35646 18116 35698
rect 17948 35644 18116 35646
rect 17388 35084 17892 35140
rect 17388 34914 17444 34926
rect 17388 34862 17390 34914
rect 17442 34862 17444 34914
rect 17276 34356 17332 34366
rect 17276 34262 17332 34300
rect 17388 33796 17444 34862
rect 17836 34468 17892 35084
rect 17500 34244 17556 34254
rect 17500 34150 17556 34188
rect 17612 34132 17668 34142
rect 17668 34076 17780 34132
rect 17612 34038 17668 34076
rect 17388 33730 17444 33740
rect 17276 33684 17332 33694
rect 17276 31220 17332 33628
rect 17724 33570 17780 34076
rect 17836 33908 17892 34412
rect 17836 33842 17892 33852
rect 17724 33518 17726 33570
rect 17778 33518 17780 33570
rect 17724 33506 17780 33518
rect 17388 33234 17444 33246
rect 17388 33182 17390 33234
rect 17442 33182 17444 33234
rect 17388 32676 17444 33182
rect 17388 32340 17444 32620
rect 17948 32674 18004 32686
rect 17948 32622 17950 32674
rect 18002 32622 18004 32674
rect 17612 32562 17668 32574
rect 17612 32510 17614 32562
rect 17666 32510 17668 32562
rect 17612 32452 17668 32510
rect 17612 32386 17668 32396
rect 17500 32340 17556 32350
rect 17388 32338 17556 32340
rect 17388 32286 17502 32338
rect 17554 32286 17556 32338
rect 17388 32284 17556 32286
rect 17500 32274 17556 32284
rect 17948 32116 18004 32622
rect 18060 32228 18116 35644
rect 18508 35698 18564 35710
rect 18508 35646 18510 35698
rect 18562 35646 18564 35698
rect 18508 35476 18564 35646
rect 18620 35476 18676 36764
rect 18844 35700 18900 35710
rect 18844 35606 18900 35644
rect 18956 35588 19012 41132
rect 19180 41186 19236 42030
rect 19292 41972 19348 41982
rect 19292 41878 19348 41916
rect 20076 41970 20132 42140
rect 20076 41918 20078 41970
rect 20130 41918 20132 41970
rect 20076 41906 20132 41918
rect 20300 41972 20356 42478
rect 20524 42420 20580 44044
rect 20636 43876 20692 44158
rect 20636 43810 20692 43820
rect 20748 44940 21140 44996
rect 20636 43540 20692 43550
rect 20748 43540 20804 44940
rect 20636 43538 20804 43540
rect 20636 43486 20638 43538
rect 20690 43486 20804 43538
rect 20636 43484 20804 43486
rect 20636 43428 20692 43484
rect 20636 43362 20692 43372
rect 21196 42756 21252 51212
rect 21532 50428 21588 51436
rect 21644 51268 21700 51996
rect 21644 51202 21700 51212
rect 21756 51156 21812 52780
rect 21868 52724 21924 54348
rect 21868 52658 21924 52668
rect 21980 53842 22036 53854
rect 21980 53790 21982 53842
rect 22034 53790 22036 53842
rect 21868 52162 21924 52174
rect 21868 52110 21870 52162
rect 21922 52110 21924 52162
rect 21868 51380 21924 52110
rect 21868 51314 21924 51324
rect 21756 51100 21924 51156
rect 21868 50594 21924 51100
rect 21868 50542 21870 50594
rect 21922 50542 21924 50594
rect 21756 50484 21812 50522
rect 21532 50372 21700 50428
rect 21756 50418 21812 50428
rect 21308 50260 21364 50270
rect 21364 50204 21476 50260
rect 21308 50194 21364 50204
rect 21420 49924 21476 50204
rect 21644 50148 21700 50372
rect 21868 50260 21924 50542
rect 21644 50082 21700 50092
rect 21756 50204 21924 50260
rect 21420 49922 21700 49924
rect 21420 49870 21422 49922
rect 21474 49870 21700 49922
rect 21420 49868 21700 49870
rect 21420 49858 21476 49868
rect 21308 49700 21364 49710
rect 21308 49250 21364 49644
rect 21308 49198 21310 49250
rect 21362 49198 21364 49250
rect 21308 49186 21364 49198
rect 21532 49364 21588 49374
rect 21420 49140 21476 49150
rect 21420 49046 21476 49084
rect 21308 47572 21364 47582
rect 21308 47458 21364 47516
rect 21308 47406 21310 47458
rect 21362 47406 21364 47458
rect 21308 47394 21364 47406
rect 21420 47348 21476 47358
rect 21532 47348 21588 49308
rect 21644 49252 21700 49868
rect 21756 49810 21812 50204
rect 21756 49758 21758 49810
rect 21810 49758 21812 49810
rect 21756 49746 21812 49758
rect 21756 49252 21812 49262
rect 21644 49250 21812 49252
rect 21644 49198 21758 49250
rect 21810 49198 21812 49250
rect 21644 49196 21812 49198
rect 21756 49186 21812 49196
rect 21420 47346 21588 47348
rect 21420 47294 21422 47346
rect 21474 47294 21588 47346
rect 21420 47292 21588 47294
rect 21756 48916 21812 48926
rect 21756 47348 21812 48860
rect 21980 47572 22036 53790
rect 22204 53842 22260 53854
rect 22204 53790 22206 53842
rect 22258 53790 22260 53842
rect 22204 53620 22260 53790
rect 22092 53564 22204 53620
rect 22092 52276 22148 53564
rect 22204 53554 22260 53564
rect 22316 53730 22372 53742
rect 22316 53678 22318 53730
rect 22370 53678 22372 53730
rect 22316 53508 22372 53678
rect 22428 53508 22484 54460
rect 22540 53844 22596 54460
rect 22540 53778 22596 53788
rect 22652 53620 22708 55580
rect 22764 55300 22820 56030
rect 22764 53956 22820 55244
rect 22988 55188 23044 56142
rect 23100 56084 23156 56590
rect 23548 56420 23604 56924
rect 23100 56018 23156 56028
rect 23436 56364 23604 56420
rect 23660 56756 23716 56766
rect 23436 56082 23492 56364
rect 23660 56306 23716 56700
rect 23884 56532 23940 57372
rect 23996 56868 24052 58828
rect 24108 58434 24164 58446
rect 24108 58382 24110 58434
rect 24162 58382 24164 58434
rect 24108 57652 24164 58382
rect 24108 57586 24164 57596
rect 23996 56754 24052 56812
rect 24108 57428 24164 57438
rect 24108 56866 24164 57372
rect 24108 56814 24110 56866
rect 24162 56814 24164 56866
rect 24108 56802 24164 56814
rect 23996 56702 23998 56754
rect 24050 56702 24052 56754
rect 23996 56690 24052 56702
rect 23884 56476 24052 56532
rect 23660 56254 23662 56306
rect 23714 56254 23716 56306
rect 23660 56242 23716 56254
rect 23548 56196 23604 56206
rect 23548 56102 23604 56140
rect 23436 56030 23438 56082
rect 23490 56030 23492 56082
rect 23436 56018 23492 56030
rect 23100 55858 23156 55870
rect 23100 55806 23102 55858
rect 23154 55806 23156 55858
rect 23100 55300 23156 55806
rect 23772 55412 23828 55422
rect 23772 55318 23828 55356
rect 23436 55300 23492 55310
rect 23100 55298 23492 55300
rect 23100 55246 23438 55298
rect 23490 55246 23492 55298
rect 23100 55244 23492 55246
rect 23436 55234 23492 55244
rect 23884 55300 23940 55310
rect 22988 55122 23044 55132
rect 23100 55076 23156 55086
rect 23100 54982 23156 55020
rect 23212 54740 23268 54750
rect 23268 54684 23380 54740
rect 23212 54674 23268 54684
rect 22764 53890 22820 53900
rect 22988 54290 23044 54302
rect 22988 54238 22990 54290
rect 23042 54238 23044 54290
rect 22652 53554 22708 53564
rect 22428 53452 22596 53508
rect 22316 53442 22372 53452
rect 22204 53060 22260 53070
rect 22204 52724 22260 53004
rect 22204 52668 22484 52724
rect 22204 52276 22260 52286
rect 22092 52274 22260 52276
rect 22092 52222 22206 52274
rect 22258 52222 22260 52274
rect 22092 52220 22260 52222
rect 22204 52210 22260 52220
rect 22316 51156 22372 51166
rect 22316 49700 22372 51100
rect 22428 50428 22484 52668
rect 22540 50818 22596 53452
rect 22988 52388 23044 54238
rect 23212 53172 23268 53182
rect 23212 52946 23268 53116
rect 23212 52894 23214 52946
rect 23266 52894 23268 52946
rect 23212 52882 23268 52894
rect 23324 52834 23380 54684
rect 23884 54626 23940 55244
rect 23884 54574 23886 54626
rect 23938 54574 23940 54626
rect 23884 54562 23940 54574
rect 23324 52782 23326 52834
rect 23378 52782 23380 52834
rect 23324 52770 23380 52782
rect 23436 54514 23492 54526
rect 23436 54462 23438 54514
rect 23490 54462 23492 54514
rect 23100 52388 23156 52398
rect 22876 52386 23156 52388
rect 22876 52334 23102 52386
rect 23154 52334 23156 52386
rect 22876 52332 23156 52334
rect 22540 50766 22542 50818
rect 22594 50766 22596 50818
rect 22540 50754 22596 50766
rect 22652 51266 22708 51278
rect 22652 51214 22654 51266
rect 22706 51214 22708 51266
rect 22652 50708 22708 51214
rect 22876 50818 22932 52332
rect 23100 52322 23156 52332
rect 23324 52276 23380 52286
rect 23436 52276 23492 54462
rect 23996 54180 24052 56476
rect 24220 56196 24276 59052
rect 24556 58884 24612 58894
rect 24556 57874 24612 58828
rect 24668 58660 24724 59612
rect 25004 59220 25060 59726
rect 25228 59668 25284 59678
rect 25284 59612 25396 59668
rect 25228 59602 25284 59612
rect 25004 59154 25060 59164
rect 24892 58660 24948 58670
rect 24668 58658 24948 58660
rect 24668 58606 24894 58658
rect 24946 58606 24948 58658
rect 24668 58604 24948 58606
rect 24780 58434 24836 58446
rect 24780 58382 24782 58434
rect 24834 58382 24836 58434
rect 24556 57822 24558 57874
rect 24610 57822 24612 57874
rect 24556 57810 24612 57822
rect 24668 58212 24724 58222
rect 24668 57874 24724 58156
rect 24668 57822 24670 57874
rect 24722 57822 24724 57874
rect 24332 57764 24388 57802
rect 24332 57698 24388 57708
rect 24444 57762 24500 57774
rect 24444 57710 24446 57762
rect 24498 57710 24500 57762
rect 24444 57204 24500 57710
rect 24668 57316 24724 57822
rect 24780 57428 24836 58382
rect 24780 57362 24836 57372
rect 24668 57250 24724 57260
rect 24444 57138 24500 57148
rect 24556 56756 24612 56766
rect 24556 56662 24612 56700
rect 24332 56642 24388 56654
rect 24332 56590 24334 56642
rect 24386 56590 24388 56642
rect 24332 56420 24388 56590
rect 24444 56644 24500 56654
rect 24444 56550 24500 56588
rect 24332 56354 24388 56364
rect 24220 56130 24276 56140
rect 24332 56196 24388 56206
rect 24332 56194 24500 56196
rect 24332 56142 24334 56194
rect 24386 56142 24500 56194
rect 24332 56140 24500 56142
rect 24332 56130 24388 56140
rect 24444 55972 24500 56140
rect 24444 55906 24500 55916
rect 24892 55972 24948 58604
rect 25004 58548 25060 58558
rect 25004 58434 25060 58492
rect 25004 58382 25006 58434
rect 25058 58382 25060 58434
rect 25004 57652 25060 58382
rect 25004 57586 25060 57596
rect 25116 57988 25172 57998
rect 25116 56756 25172 57932
rect 25116 56690 25172 56700
rect 25228 57092 25284 57102
rect 25228 56082 25284 57036
rect 25228 56030 25230 56082
rect 25282 56030 25284 56082
rect 25228 56018 25284 56030
rect 24892 55906 24948 55916
rect 24332 55860 24388 55870
rect 24220 55298 24276 55310
rect 24220 55246 24222 55298
rect 24274 55246 24276 55298
rect 24220 55188 24276 55246
rect 24220 55122 24276 55132
rect 24332 54514 24388 55804
rect 25340 55636 25396 59612
rect 25116 55580 25396 55636
rect 24780 55300 24836 55310
rect 24780 55206 24836 55244
rect 24556 54628 24612 54638
rect 25116 54628 25172 55580
rect 25340 55412 25396 55450
rect 25340 55346 25396 55356
rect 25228 55298 25284 55310
rect 25228 55246 25230 55298
rect 25282 55246 25284 55298
rect 25228 54964 25284 55246
rect 25228 54898 25284 54908
rect 24556 54626 25284 54628
rect 24556 54574 24558 54626
rect 24610 54574 25284 54626
rect 24556 54572 25284 54574
rect 24556 54562 24612 54572
rect 24332 54462 24334 54514
rect 24386 54462 24388 54514
rect 24332 54450 24388 54462
rect 25116 54404 25172 54414
rect 24668 54290 24724 54302
rect 24668 54238 24670 54290
rect 24722 54238 24724 54290
rect 24668 54180 24724 54238
rect 23884 54124 24724 54180
rect 23548 54068 23604 54078
rect 23548 52836 23604 54012
rect 23548 52770 23604 52780
rect 23548 52612 23604 52622
rect 23604 52556 23716 52612
rect 23548 52546 23604 52556
rect 23324 52274 23492 52276
rect 23324 52222 23326 52274
rect 23378 52222 23492 52274
rect 23324 52220 23492 52222
rect 23324 52210 23380 52220
rect 23436 51602 23492 52220
rect 23660 52162 23716 52556
rect 23660 52110 23662 52162
rect 23714 52110 23716 52162
rect 23660 52098 23716 52110
rect 23884 51940 23940 54124
rect 23996 53956 24052 53966
rect 23996 53862 24052 53900
rect 25116 53844 25172 54348
rect 25228 54402 25284 54572
rect 25228 54350 25230 54402
rect 25282 54350 25284 54402
rect 25228 54338 25284 54350
rect 25452 54292 25508 60508
rect 26236 59444 26292 63200
rect 27580 60114 27636 60126
rect 27580 60062 27582 60114
rect 27634 60062 27636 60114
rect 27356 59892 27412 59902
rect 27356 59798 27412 59836
rect 26348 59778 26404 59790
rect 26348 59726 26350 59778
rect 26402 59726 26404 59778
rect 26348 59668 26404 59726
rect 26348 59602 26404 59612
rect 26236 59378 26292 59388
rect 27468 59444 27524 59454
rect 27468 59350 27524 59388
rect 25564 59220 25620 59230
rect 25564 59126 25620 59164
rect 26460 59218 26516 59230
rect 26460 59166 26462 59218
rect 26514 59166 26516 59218
rect 26124 58996 26180 59006
rect 26124 58902 26180 58940
rect 26460 58100 26516 59166
rect 26796 58996 26852 59006
rect 26460 58034 26516 58044
rect 26684 58210 26740 58222
rect 26684 58158 26686 58210
rect 26738 58158 26740 58210
rect 26684 57876 26740 58158
rect 25900 57820 26740 57876
rect 25676 57652 25732 57662
rect 25900 57652 25956 57820
rect 26796 57764 26852 58940
rect 27020 58436 27076 58446
rect 27020 58342 27076 58380
rect 26684 57708 26852 57764
rect 25676 57650 25956 57652
rect 25676 57598 25678 57650
rect 25730 57598 25956 57650
rect 25676 57596 25956 57598
rect 26012 57652 26068 57662
rect 25676 57586 25732 57596
rect 25676 57090 25732 57102
rect 25676 57038 25678 57090
rect 25730 57038 25732 57090
rect 25676 56980 25732 57038
rect 25676 56914 25732 56924
rect 25676 56308 25732 56318
rect 25564 56196 25620 56206
rect 25564 56102 25620 56140
rect 25676 55298 25732 56252
rect 25788 56082 25844 57596
rect 26012 57558 26068 57596
rect 26124 57538 26180 57550
rect 26124 57486 26126 57538
rect 26178 57486 26180 57538
rect 25788 56030 25790 56082
rect 25842 56030 25844 56082
rect 25788 56018 25844 56030
rect 25900 56084 25956 56094
rect 26124 56084 26180 57486
rect 26460 57316 26516 57326
rect 26460 56978 26516 57260
rect 26460 56926 26462 56978
rect 26514 56926 26516 56978
rect 26460 56914 26516 56926
rect 26684 56866 26740 57708
rect 26684 56814 26686 56866
rect 26738 56814 26740 56866
rect 26684 56802 26740 56814
rect 27020 56868 27076 56878
rect 27020 56194 27076 56812
rect 27580 56868 27636 60062
rect 28588 60002 28644 60014
rect 28588 59950 28590 60002
rect 28642 59950 28644 60002
rect 28140 59780 28196 59790
rect 27804 59220 27860 59230
rect 27692 59164 27804 59220
rect 27692 58322 27748 59164
rect 27804 59154 27860 59164
rect 27916 59108 27972 59118
rect 27804 58996 27860 59006
rect 27804 58436 27860 58940
rect 27804 58342 27860 58380
rect 27692 58270 27694 58322
rect 27746 58270 27748 58322
rect 27692 58258 27748 58270
rect 27916 58212 27972 59052
rect 27804 58156 27972 58212
rect 28028 58660 28084 58670
rect 27580 56774 27636 56812
rect 27692 56980 27748 56990
rect 27468 56196 27524 56206
rect 27020 56142 27022 56194
rect 27074 56142 27076 56194
rect 27020 56130 27076 56142
rect 27244 56194 27524 56196
rect 27244 56142 27470 56194
rect 27522 56142 27524 56194
rect 27244 56140 27524 56142
rect 25956 56028 26180 56084
rect 25900 55990 25956 56028
rect 27244 55468 27300 56140
rect 27468 56130 27524 56140
rect 27692 56196 27748 56924
rect 27804 56532 27860 58156
rect 28028 57764 28084 58604
rect 28028 56754 28084 57708
rect 28140 57650 28196 59724
rect 28364 59778 28420 59790
rect 28364 59726 28366 59778
rect 28418 59726 28420 59778
rect 28364 58772 28420 59726
rect 28364 58706 28420 58716
rect 28588 58436 28644 59950
rect 29596 60004 29652 63200
rect 38332 62188 38388 63200
rect 38332 62132 38612 62188
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 29596 59938 29652 59948
rect 33964 60004 34020 60014
rect 33964 59910 34020 59948
rect 34972 60004 35028 60014
rect 34972 59910 35028 59948
rect 29708 59892 29764 59902
rect 29148 59668 29204 59678
rect 28588 58370 28644 58380
rect 29036 59612 29148 59668
rect 28140 57598 28142 57650
rect 28194 57598 28196 57650
rect 28140 57586 28196 57598
rect 28252 58210 28308 58222
rect 28252 58158 28254 58210
rect 28306 58158 28308 58210
rect 28028 56702 28030 56754
rect 28082 56702 28084 56754
rect 28028 56690 28084 56702
rect 27804 56476 28084 56532
rect 27692 56140 27972 56196
rect 27580 56082 27636 56094
rect 27580 56030 27582 56082
rect 27634 56030 27636 56082
rect 27468 55860 27524 55870
rect 27468 55766 27524 55804
rect 27580 55636 27636 56030
rect 25676 55246 25678 55298
rect 25730 55246 25732 55298
rect 24892 53842 25172 53844
rect 24892 53790 25118 53842
rect 25170 53790 25172 53842
rect 24892 53788 25172 53790
rect 24780 53732 24836 53742
rect 24556 53730 24836 53732
rect 24556 53678 24782 53730
rect 24834 53678 24836 53730
rect 24556 53676 24836 53678
rect 24220 52948 24276 52958
rect 24108 52892 24220 52948
rect 23436 51550 23438 51602
rect 23490 51550 23492 51602
rect 23436 51538 23492 51550
rect 23548 51884 23940 51940
rect 23996 52274 24052 52286
rect 23996 52222 23998 52274
rect 24050 52222 24052 52274
rect 23996 51940 24052 52222
rect 22988 51380 23044 51390
rect 22988 51378 23380 51380
rect 22988 51326 22990 51378
rect 23042 51326 23380 51378
rect 22988 51324 23380 51326
rect 22988 51314 23044 51324
rect 22876 50766 22878 50818
rect 22930 50766 22932 50818
rect 22876 50754 22932 50766
rect 22652 50652 22820 50708
rect 22764 50596 22820 50652
rect 22428 50372 22708 50428
rect 22428 49924 22484 49934
rect 22652 49924 22708 50372
rect 22428 49922 22708 49924
rect 22428 49870 22430 49922
rect 22482 49870 22708 49922
rect 22428 49868 22708 49870
rect 22428 49858 22484 49868
rect 22764 49810 22820 50540
rect 22764 49758 22766 49810
rect 22818 49758 22820 49810
rect 22316 49644 22484 49700
rect 22092 49026 22148 49038
rect 22092 48974 22094 49026
rect 22146 48974 22148 49026
rect 22092 48468 22148 48974
rect 22092 48402 22148 48412
rect 22316 48914 22372 48926
rect 22316 48862 22318 48914
rect 22370 48862 22372 48914
rect 22204 48354 22260 48366
rect 22204 48302 22206 48354
rect 22258 48302 22260 48354
rect 22204 47684 22260 48302
rect 22316 48356 22372 48862
rect 22316 48290 22372 48300
rect 22204 47618 22260 47628
rect 21980 47516 22148 47572
rect 21980 47348 22036 47358
rect 21756 47346 22036 47348
rect 21756 47294 21982 47346
rect 22034 47294 22036 47346
rect 21756 47292 22036 47294
rect 21308 46564 21364 46574
rect 21308 46470 21364 46508
rect 21420 46452 21476 47292
rect 21420 46358 21476 46396
rect 21756 46676 21812 46686
rect 21420 45890 21476 45902
rect 21420 45838 21422 45890
rect 21474 45838 21476 45890
rect 21420 45444 21476 45838
rect 21420 45378 21476 45388
rect 21756 45220 21812 46620
rect 21980 45220 22036 47292
rect 22092 46228 22148 47516
rect 22092 46162 22148 46172
rect 21644 45218 21812 45220
rect 21644 45166 21758 45218
rect 21810 45166 21812 45218
rect 21644 45164 21812 45166
rect 21644 43876 21700 45164
rect 21756 45154 21812 45164
rect 21868 45164 21980 45220
rect 22092 45778 22148 45790
rect 22092 45726 22094 45778
rect 22146 45726 22148 45778
rect 22092 45220 22148 45726
rect 22428 45332 22484 49644
rect 22764 49026 22820 49758
rect 22764 48974 22766 49026
rect 22818 48974 22820 49026
rect 22764 48962 22820 48974
rect 23324 50594 23380 51324
rect 23324 50542 23326 50594
rect 23378 50542 23380 50594
rect 23324 48468 23380 50542
rect 23324 48374 23380 48412
rect 23548 48356 23604 51884
rect 23996 51874 24052 51884
rect 23772 51380 23828 51390
rect 23996 51380 24052 51390
rect 23772 51378 23996 51380
rect 23772 51326 23774 51378
rect 23826 51326 23996 51378
rect 23772 51324 23996 51326
rect 23772 51314 23828 51324
rect 23996 51314 24052 51324
rect 24108 50428 24164 52892
rect 24220 52882 24276 52892
rect 24220 52612 24276 52622
rect 24220 52050 24276 52556
rect 24220 51998 24222 52050
rect 24274 51998 24276 52050
rect 24220 51986 24276 51998
rect 24332 52164 24388 52174
rect 24332 50818 24388 52108
rect 24556 52050 24612 53676
rect 24780 53666 24836 53676
rect 24556 51998 24558 52050
rect 24610 51998 24612 52050
rect 24556 51716 24612 51998
rect 24332 50766 24334 50818
rect 24386 50766 24388 50818
rect 24332 50754 24388 50766
rect 24444 51660 24612 51716
rect 24780 52052 24836 52062
rect 24892 52052 24948 53788
rect 25116 53778 25172 53788
rect 25340 54236 25508 54292
rect 25564 55186 25620 55198
rect 25564 55134 25566 55186
rect 25618 55134 25620 55186
rect 25228 53620 25284 53630
rect 25228 53058 25284 53564
rect 25340 53396 25396 54236
rect 25452 53956 25508 53966
rect 25564 53956 25620 55134
rect 25676 55076 25732 55246
rect 25676 55010 25732 55020
rect 26572 55412 26628 55422
rect 26572 55298 26628 55356
rect 26572 55246 26574 55298
rect 26626 55246 26628 55298
rect 26236 54516 26292 54526
rect 25508 53900 25620 53956
rect 26124 54460 26236 54516
rect 25452 53890 25508 53900
rect 25900 53844 25956 53854
rect 25340 53170 25396 53340
rect 25340 53118 25342 53170
rect 25394 53118 25396 53170
rect 25340 53106 25396 53118
rect 25452 53730 25508 53742
rect 25452 53678 25454 53730
rect 25506 53678 25508 53730
rect 25228 53006 25230 53058
rect 25282 53006 25284 53058
rect 25228 52994 25284 53006
rect 25340 52836 25396 52846
rect 25340 52162 25396 52780
rect 25340 52110 25342 52162
rect 25394 52110 25396 52162
rect 25340 52098 25396 52110
rect 25452 52164 25508 53678
rect 25788 53172 25844 53182
rect 25788 53078 25844 53116
rect 25900 53170 25956 53788
rect 25900 53118 25902 53170
rect 25954 53118 25956 53170
rect 25900 53106 25956 53118
rect 25452 52098 25508 52108
rect 25564 52946 25620 52958
rect 25564 52894 25566 52946
rect 25618 52894 25620 52946
rect 24780 52050 24948 52052
rect 24780 51998 24782 52050
rect 24834 51998 24948 52050
rect 24780 51996 24948 51998
rect 24444 51604 24500 51660
rect 24444 51378 24500 51548
rect 24444 51326 24446 51378
rect 24498 51326 24500 51378
rect 24444 50594 24500 51326
rect 24444 50542 24446 50594
rect 24498 50542 24500 50594
rect 24444 50530 24500 50542
rect 24556 51490 24612 51502
rect 24556 51438 24558 51490
rect 24610 51438 24612 51490
rect 23436 48300 23604 48356
rect 23660 50370 23716 50382
rect 24108 50372 24276 50428
rect 23660 50318 23662 50370
rect 23714 50318 23716 50370
rect 22540 47572 22596 47582
rect 23436 47572 23492 48300
rect 23660 48244 23716 50318
rect 24108 50260 24164 50270
rect 24108 49810 24164 50204
rect 24108 49758 24110 49810
rect 24162 49758 24164 49810
rect 24108 49026 24164 49758
rect 24108 48974 24110 49026
rect 24162 48974 24164 49026
rect 23884 48804 23940 48814
rect 23548 48188 23716 48244
rect 23772 48356 23828 48366
rect 23772 48242 23828 48300
rect 23772 48190 23774 48242
rect 23826 48190 23828 48242
rect 23548 47796 23604 48188
rect 23772 48178 23828 48190
rect 23548 47730 23604 47740
rect 23660 48020 23716 48030
rect 23436 47516 23604 47572
rect 22540 47478 22596 47516
rect 23324 47346 23380 47358
rect 23324 47294 23326 47346
rect 23378 47294 23380 47346
rect 22988 47234 23044 47246
rect 22988 47182 22990 47234
rect 23042 47182 23044 47234
rect 22988 46900 23044 47182
rect 22988 46834 23044 46844
rect 23324 46900 23380 47294
rect 23324 46834 23380 46844
rect 22876 46788 22932 46798
rect 22876 46694 22932 46732
rect 22764 46674 22820 46686
rect 22764 46622 22766 46674
rect 22818 46622 22820 46674
rect 22764 45444 22820 46622
rect 22988 46676 23044 46686
rect 23324 46676 23380 46686
rect 22988 46674 23268 46676
rect 22988 46622 22990 46674
rect 23042 46622 23268 46674
rect 22988 46620 23268 46622
rect 22988 46610 23044 46620
rect 23212 45892 23268 46620
rect 23324 46582 23380 46620
rect 23212 45836 23380 45892
rect 23212 45668 23268 45678
rect 22764 45388 23156 45444
rect 22428 45276 23044 45332
rect 22092 45164 22820 45220
rect 21756 44436 21812 44446
rect 21756 44322 21812 44380
rect 21756 44270 21758 44322
rect 21810 44270 21812 44322
rect 21756 44258 21812 44270
rect 21644 43820 21812 43876
rect 21644 43652 21700 43662
rect 21196 42690 21252 42700
rect 21308 43650 21700 43652
rect 21308 43598 21646 43650
rect 21698 43598 21700 43650
rect 21308 43596 21700 43598
rect 20524 42354 20580 42364
rect 20860 42532 20916 42542
rect 20300 41906 20356 41916
rect 20524 42082 20580 42094
rect 20524 42030 20526 42082
rect 20578 42030 20580 42082
rect 19180 41134 19182 41186
rect 19234 41134 19236 41186
rect 19068 40964 19124 40974
rect 19068 40292 19124 40908
rect 19180 40628 19236 41134
rect 19404 41860 19460 41870
rect 19404 41074 19460 41804
rect 20524 41860 20580 42030
rect 20748 41972 20804 41982
rect 20748 41878 20804 41916
rect 20524 41794 20580 41804
rect 19740 41748 19796 41758
rect 19740 41076 19796 41692
rect 20748 41300 20804 41310
rect 20860 41300 20916 42476
rect 19404 41022 19406 41074
rect 19458 41022 19460 41074
rect 19404 41010 19460 41022
rect 19628 41074 19796 41076
rect 19628 41022 19742 41074
rect 19794 41022 19796 41074
rect 19628 41020 19796 41022
rect 19516 40628 19572 40638
rect 19180 40626 19572 40628
rect 19180 40574 19518 40626
rect 19570 40574 19572 40626
rect 19180 40572 19572 40574
rect 19516 40562 19572 40572
rect 19628 40404 19684 41020
rect 19740 41010 19796 41020
rect 20524 41298 20916 41300
rect 20524 41246 20750 41298
rect 20802 41246 20916 41298
rect 20524 41244 20916 41246
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19068 39620 19124 40236
rect 19516 40348 19684 40404
rect 20188 40402 20244 40414
rect 20188 40350 20190 40402
rect 20242 40350 20244 40402
rect 19292 39620 19348 39630
rect 19068 39618 19348 39620
rect 19068 39566 19294 39618
rect 19346 39566 19348 39618
rect 19068 39564 19348 39566
rect 19292 39554 19348 39564
rect 19404 39284 19460 39294
rect 19180 38836 19236 38846
rect 19180 38742 19236 38780
rect 19404 38834 19460 39228
rect 19404 38782 19406 38834
rect 19458 38782 19460 38834
rect 19404 38770 19460 38782
rect 19516 38668 19572 40348
rect 20188 40292 20244 40350
rect 20188 40226 20244 40236
rect 20412 40404 20468 40414
rect 20412 39618 20468 40348
rect 20412 39566 20414 39618
rect 20466 39566 20468 39618
rect 20412 39554 20468 39566
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20412 39060 20468 39070
rect 20524 39060 20580 41244
rect 20748 41234 20804 41244
rect 20636 41076 20692 41086
rect 20636 40962 20692 41020
rect 20636 40910 20638 40962
rect 20690 40910 20692 40962
rect 20636 40852 20692 40910
rect 20636 40786 20692 40796
rect 21308 39844 21364 43596
rect 21644 43586 21700 43596
rect 21756 43652 21812 43820
rect 21756 43586 21812 43596
rect 21868 43540 21924 45164
rect 21980 45154 22036 45164
rect 22652 44996 22708 45006
rect 22652 44902 22708 44940
rect 22764 44882 22820 45164
rect 22764 44830 22766 44882
rect 22818 44830 22820 44882
rect 22764 44818 22820 44830
rect 22876 45106 22932 45118
rect 22876 45054 22878 45106
rect 22930 45054 22932 45106
rect 22876 44772 22932 45054
rect 22876 44706 22932 44716
rect 21868 43474 21924 43484
rect 21980 44322 22036 44334
rect 21980 44270 21982 44322
rect 22034 44270 22036 44322
rect 21532 43092 21588 43102
rect 21532 42866 21588 43036
rect 21980 42980 22036 44270
rect 22316 44324 22372 44334
rect 22316 44230 22372 44268
rect 22092 44098 22148 44110
rect 22092 44046 22094 44098
rect 22146 44046 22148 44098
rect 22092 43540 22148 44046
rect 22092 43474 22148 43484
rect 22540 44098 22596 44110
rect 22540 44046 22542 44098
rect 22594 44046 22596 44098
rect 21980 42914 22036 42924
rect 21532 42814 21534 42866
rect 21586 42814 21588 42866
rect 21420 42084 21476 42094
rect 21420 41990 21476 42028
rect 21532 41076 21588 42814
rect 21980 42532 22036 42542
rect 21980 42438 22036 42476
rect 21756 42196 21812 42206
rect 21644 41970 21700 41982
rect 21644 41918 21646 41970
rect 21698 41918 21700 41970
rect 21644 41860 21700 41918
rect 21644 41794 21700 41804
rect 21756 41298 21812 42140
rect 22428 41972 22484 41982
rect 22428 41878 22484 41916
rect 21756 41246 21758 41298
rect 21810 41246 21812 41298
rect 21756 41234 21812 41246
rect 21868 41860 21924 41870
rect 21644 41076 21700 41086
rect 21532 41074 21700 41076
rect 21532 41022 21646 41074
rect 21698 41022 21700 41074
rect 21532 41020 21700 41022
rect 21644 40964 21700 41020
rect 21644 40898 21700 40908
rect 21756 41076 21812 41086
rect 21756 40516 21812 41020
rect 21868 41074 21924 41804
rect 22540 41860 22596 44046
rect 22652 42980 22708 42990
rect 22652 42866 22708 42924
rect 22652 42814 22654 42866
rect 22706 42814 22708 42866
rect 22652 42802 22708 42814
rect 22764 41972 22820 41982
rect 22092 41748 22148 41758
rect 22092 41186 22148 41692
rect 22092 41134 22094 41186
rect 22146 41134 22148 41186
rect 22092 41122 22148 41134
rect 22540 41188 22596 41804
rect 22652 41970 22820 41972
rect 22652 41918 22766 41970
rect 22818 41918 22820 41970
rect 22652 41916 22820 41918
rect 22652 41412 22708 41916
rect 22764 41906 22820 41916
rect 22988 41748 23044 45276
rect 23100 45108 23156 45388
rect 23100 45042 23156 45052
rect 23212 45106 23268 45612
rect 23324 45332 23380 45836
rect 23324 45266 23380 45276
rect 23212 45054 23214 45106
rect 23266 45054 23268 45106
rect 23212 45042 23268 45054
rect 23436 45108 23492 45118
rect 23436 45014 23492 45052
rect 23548 44660 23604 47516
rect 23660 47570 23716 47964
rect 23660 47518 23662 47570
rect 23714 47518 23716 47570
rect 23660 47506 23716 47518
rect 23772 46676 23828 46686
rect 23884 46676 23940 48748
rect 23996 48468 24052 48478
rect 23996 48242 24052 48412
rect 23996 48190 23998 48242
rect 24050 48190 24052 48242
rect 23996 48178 24052 48190
rect 23996 47796 24052 47806
rect 23996 47012 24052 47740
rect 24108 47682 24164 48974
rect 24108 47630 24110 47682
rect 24162 47630 24164 47682
rect 24108 47618 24164 47630
rect 23996 46956 24164 47012
rect 23772 46674 23940 46676
rect 23772 46622 23774 46674
rect 23826 46622 23940 46674
rect 23772 46620 23940 46622
rect 23996 46786 24052 46798
rect 23996 46734 23998 46786
rect 24050 46734 24052 46786
rect 23772 46610 23828 46620
rect 23884 46228 23940 46238
rect 23548 44594 23604 44604
rect 23772 46116 23828 46126
rect 23772 44436 23828 46060
rect 23884 45556 23940 46172
rect 23996 45892 24052 46734
rect 23996 45826 24052 45836
rect 23884 45218 23940 45500
rect 23884 45166 23886 45218
rect 23938 45166 23940 45218
rect 23884 45154 23940 45166
rect 24108 45332 24164 46956
rect 24220 46002 24276 50372
rect 24556 50036 24612 51438
rect 24780 51380 24836 51996
rect 25452 51716 25508 51726
rect 25228 51604 25284 51614
rect 25228 51510 25284 51548
rect 24780 51314 24836 51324
rect 25452 51378 25508 51660
rect 25564 51604 25620 52894
rect 26012 52946 26068 52958
rect 26012 52894 26014 52946
rect 26066 52894 26068 52946
rect 26012 52500 26068 52894
rect 26012 52434 26068 52444
rect 26124 52276 26180 54460
rect 26236 54450 26292 54460
rect 26572 53956 26628 55246
rect 27020 55412 27300 55468
rect 27356 55580 27580 55636
rect 26684 55188 26740 55198
rect 26684 55094 26740 55132
rect 26908 55076 26964 55086
rect 26908 54982 26964 55020
rect 26572 53890 26628 53900
rect 26684 53732 26740 53742
rect 27020 53732 27076 55412
rect 26740 53676 27076 53732
rect 27132 55300 27188 55310
rect 27132 53732 27188 55244
rect 27356 54628 27412 55580
rect 27580 55570 27636 55580
rect 27244 54572 27412 54628
rect 27468 55412 27524 55422
rect 27244 54292 27300 54572
rect 27244 54226 27300 54236
rect 27356 54402 27412 54414
rect 27356 54350 27358 54402
rect 27410 54350 27412 54402
rect 27356 53844 27412 54350
rect 27356 53778 27412 53788
rect 27244 53732 27300 53742
rect 27132 53730 27300 53732
rect 27132 53678 27246 53730
rect 27298 53678 27300 53730
rect 27132 53676 27300 53678
rect 26684 53638 26740 53676
rect 27244 53666 27300 53676
rect 27468 53730 27524 55356
rect 27692 55298 27748 56140
rect 27916 56082 27972 56140
rect 27916 56030 27918 56082
rect 27970 56030 27972 56082
rect 27916 56018 27972 56030
rect 27692 55246 27694 55298
rect 27746 55246 27748 55298
rect 27692 55234 27748 55246
rect 27804 55748 27860 55758
rect 27804 55186 27860 55692
rect 27804 55134 27806 55186
rect 27858 55134 27860 55186
rect 27804 55122 27860 55134
rect 27916 55524 27972 55534
rect 28028 55524 28084 56476
rect 28140 56194 28196 56206
rect 28140 56142 28142 56194
rect 28194 56142 28196 56194
rect 28140 55748 28196 56142
rect 28140 55682 28196 55692
rect 28028 55468 28196 55524
rect 27804 54628 27860 54638
rect 27692 54180 27748 54190
rect 27468 53678 27470 53730
rect 27522 53678 27524 53730
rect 27468 53666 27524 53678
rect 27580 54124 27692 54180
rect 26460 53508 26516 53518
rect 26460 52946 26516 53452
rect 27580 53506 27636 54124
rect 27692 54114 27748 54124
rect 27692 53956 27748 53966
rect 27692 53862 27748 53900
rect 27580 53454 27582 53506
rect 27634 53454 27636 53506
rect 27580 53442 27636 53454
rect 27020 53172 27076 53182
rect 27020 53078 27076 53116
rect 26684 53060 26740 53070
rect 26684 53058 26852 53060
rect 26684 53006 26686 53058
rect 26738 53006 26852 53058
rect 26684 53004 26852 53006
rect 26684 52994 26740 53004
rect 26460 52894 26462 52946
rect 26514 52894 26516 52946
rect 26460 52882 26516 52894
rect 26012 52220 26180 52276
rect 26572 52500 26628 52510
rect 26012 51828 26068 52220
rect 26124 52052 26180 52062
rect 26124 52050 26516 52052
rect 26124 51998 26126 52050
rect 26178 51998 26516 52050
rect 26124 51996 26516 51998
rect 26124 51986 26180 51996
rect 26012 51772 26292 51828
rect 25564 51538 25620 51548
rect 25452 51326 25454 51378
rect 25506 51326 25508 51378
rect 25452 51314 25508 51326
rect 25564 51212 25956 51268
rect 25004 50482 25060 50494
rect 25004 50430 25006 50482
rect 25058 50430 25060 50482
rect 25004 50428 25060 50430
rect 25004 50372 25172 50428
rect 24556 49970 24612 49980
rect 25116 49812 25172 50372
rect 25228 49812 25284 49822
rect 25116 49810 25284 49812
rect 25116 49758 25230 49810
rect 25282 49758 25284 49810
rect 25116 49756 25284 49758
rect 24668 49698 24724 49710
rect 24668 49646 24670 49698
rect 24722 49646 24724 49698
rect 24444 49028 24500 49038
rect 24332 49026 24500 49028
rect 24332 48974 24446 49026
rect 24498 48974 24500 49026
rect 24332 48972 24500 48974
rect 24332 48466 24388 48972
rect 24444 48962 24500 48972
rect 24332 48414 24334 48466
rect 24386 48414 24388 48466
rect 24332 48402 24388 48414
rect 24556 48914 24612 48926
rect 24556 48862 24558 48914
rect 24610 48862 24612 48914
rect 24444 47460 24500 47470
rect 24444 47366 24500 47404
rect 24556 47012 24612 48862
rect 24444 46956 24612 47012
rect 24668 47012 24724 49646
rect 24780 48804 24836 48814
rect 24780 47346 24836 48748
rect 24780 47294 24782 47346
rect 24834 47294 24836 47346
rect 24780 47282 24836 47294
rect 25004 47684 25060 47694
rect 25004 47346 25060 47628
rect 25004 47294 25006 47346
rect 25058 47294 25060 47346
rect 25004 47282 25060 47294
rect 24332 46676 24388 46686
rect 24332 46582 24388 46620
rect 24444 46452 24500 46956
rect 24668 46946 24724 46956
rect 24556 46788 24612 46798
rect 24556 46694 24612 46732
rect 24220 45950 24222 46002
rect 24274 45950 24276 46002
rect 24220 45938 24276 45950
rect 24332 46396 24500 46452
rect 24668 46562 24724 46574
rect 24668 46510 24670 46562
rect 24722 46510 24724 46562
rect 24108 45218 24164 45276
rect 24332 45220 24388 46396
rect 24556 45892 24612 45930
rect 24556 45826 24612 45836
rect 24556 45668 24612 45678
rect 24668 45668 24724 46510
rect 25116 46340 25172 49756
rect 25228 49746 25284 49756
rect 25564 49810 25620 51212
rect 25900 51156 25956 51212
rect 26236 51156 26292 51772
rect 26348 51604 26404 51614
rect 26348 51510 26404 51548
rect 26460 51380 26516 51996
rect 26572 51602 26628 52444
rect 26572 51550 26574 51602
rect 26626 51550 26628 51602
rect 26572 51538 26628 51550
rect 26796 51828 26852 53004
rect 26796 51604 26852 51772
rect 27020 52612 27076 52622
rect 26796 51548 26964 51604
rect 26684 51380 26740 51390
rect 26460 51378 26740 51380
rect 26460 51326 26686 51378
rect 26738 51326 26740 51378
rect 26460 51324 26740 51326
rect 26684 51314 26740 51324
rect 26796 51380 26852 51390
rect 26796 51286 26852 51324
rect 26908 51156 26964 51548
rect 25900 51100 26292 51156
rect 25788 51044 25844 51054
rect 25788 50594 25844 50988
rect 25788 50542 25790 50594
rect 25842 50542 25844 50594
rect 25676 50036 25732 50046
rect 25676 49942 25732 49980
rect 25788 49812 25844 50542
rect 26236 50594 26292 51100
rect 26236 50542 26238 50594
rect 26290 50542 26292 50594
rect 26236 50530 26292 50542
rect 26796 51100 26964 51156
rect 26796 50428 26852 51100
rect 25564 49758 25566 49810
rect 25618 49758 25620 49810
rect 25340 49140 25396 49150
rect 25340 48130 25396 49084
rect 25452 48804 25508 48814
rect 25452 48710 25508 48748
rect 25340 48078 25342 48130
rect 25394 48078 25396 48130
rect 25340 47068 25396 48078
rect 25004 46284 25172 46340
rect 25228 47012 25396 47068
rect 25564 47012 25620 49758
rect 24780 46116 24836 46126
rect 24780 46022 24836 46060
rect 24556 45666 24724 45668
rect 24556 45614 24558 45666
rect 24610 45614 24724 45666
rect 24556 45612 24724 45614
rect 24556 45602 24612 45612
rect 24780 45332 24836 45342
rect 24836 45276 24948 45332
rect 24780 45266 24836 45276
rect 24108 45166 24110 45218
rect 24162 45166 24164 45218
rect 24108 45154 24164 45166
rect 24220 45164 24388 45220
rect 23996 45108 24052 45118
rect 23996 45014 24052 45052
rect 23996 44436 24052 44446
rect 23772 44434 24164 44436
rect 23772 44382 23998 44434
rect 24050 44382 24164 44434
rect 23772 44380 24164 44382
rect 23996 44370 24052 44380
rect 23100 44322 23156 44334
rect 23100 44270 23102 44322
rect 23154 44270 23156 44322
rect 23100 43314 23156 44270
rect 23212 44324 23268 44334
rect 23660 44324 23716 44334
rect 24108 44324 24164 44380
rect 23268 44268 23380 44324
rect 23212 44258 23268 44268
rect 23100 43262 23102 43314
rect 23154 43262 23156 43314
rect 23100 42756 23156 43262
rect 23100 42662 23156 42700
rect 23212 43652 23268 43662
rect 23212 42532 23268 43596
rect 22652 41346 22708 41356
rect 22764 41692 23044 41748
rect 23100 42476 23268 42532
rect 21868 41022 21870 41074
rect 21922 41022 21924 41074
rect 21868 41010 21924 41022
rect 22204 40628 22260 40638
rect 21980 40516 22036 40526
rect 21756 40514 22036 40516
rect 21756 40462 21982 40514
rect 22034 40462 22036 40514
rect 21756 40460 22036 40462
rect 21980 40450 22036 40460
rect 22092 40516 22148 40526
rect 20412 39058 20580 39060
rect 20412 39006 20414 39058
rect 20466 39006 20580 39058
rect 20412 39004 20580 39006
rect 21084 39788 21364 39844
rect 21420 40404 21476 40414
rect 21420 39842 21476 40348
rect 22092 40402 22148 40460
rect 22092 40350 22094 40402
rect 22146 40350 22148 40402
rect 22092 40338 22148 40350
rect 21420 39790 21422 39842
rect 21474 39790 21476 39842
rect 20412 38994 20468 39004
rect 20076 38948 20132 38958
rect 19852 38834 19908 38846
rect 19852 38782 19854 38834
rect 19906 38782 19908 38834
rect 19852 38668 19908 38782
rect 19404 38612 19572 38668
rect 19628 38612 19908 38668
rect 19404 37940 19460 38612
rect 19404 37874 19460 37884
rect 19516 38388 19572 38398
rect 19516 37938 19572 38332
rect 19516 37886 19518 37938
rect 19570 37886 19572 37938
rect 19516 37874 19572 37886
rect 19292 36482 19348 36494
rect 19292 36430 19294 36482
rect 19346 36430 19348 36482
rect 19292 36036 19348 36430
rect 19292 35970 19348 35980
rect 19628 36484 19684 38612
rect 20076 38388 20132 38892
rect 20412 38612 20468 38622
rect 20076 38332 20356 38388
rect 20300 38162 20356 38332
rect 20300 38110 20302 38162
rect 20354 38110 20356 38162
rect 20300 38098 20356 38110
rect 19852 38052 19908 38062
rect 19852 37958 19908 37996
rect 20412 38050 20468 38556
rect 20412 37998 20414 38050
rect 20466 37998 20468 38050
rect 20412 37986 20468 37998
rect 20748 38052 20804 38062
rect 20188 37828 20244 37838
rect 20412 37828 20468 37838
rect 20188 37826 20356 37828
rect 20188 37774 20190 37826
rect 20242 37774 20356 37826
rect 20188 37772 20356 37774
rect 20188 37762 20244 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37044 20244 37054
rect 19740 36484 19796 36494
rect 19628 36482 19796 36484
rect 19628 36430 19742 36482
rect 19794 36430 19796 36482
rect 19628 36428 19796 36430
rect 19628 35700 19684 36428
rect 19740 36418 19796 36428
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19628 35606 19684 35644
rect 19964 35588 20020 35598
rect 20188 35588 20244 36988
rect 20300 36708 20356 37772
rect 20300 36484 20356 36652
rect 20300 36418 20356 36428
rect 18956 35532 19460 35588
rect 18508 35420 19236 35476
rect 18620 34916 18676 34926
rect 18284 34802 18340 34814
rect 18284 34750 18286 34802
rect 18338 34750 18340 34802
rect 18172 34244 18228 34254
rect 18172 34150 18228 34188
rect 18284 34020 18340 34750
rect 18396 34692 18452 34702
rect 18396 34242 18452 34636
rect 18396 34190 18398 34242
rect 18450 34190 18452 34242
rect 18396 34178 18452 34190
rect 18508 34242 18564 34254
rect 18508 34190 18510 34242
rect 18562 34190 18564 34242
rect 18396 34020 18452 34030
rect 18284 34018 18452 34020
rect 18284 33966 18398 34018
rect 18450 33966 18452 34018
rect 18284 33964 18452 33966
rect 18396 33954 18452 33964
rect 18172 33908 18228 33918
rect 18228 33852 18340 33908
rect 18172 33842 18228 33852
rect 18060 32162 18116 32172
rect 18172 33124 18228 33134
rect 17500 32060 18004 32116
rect 17500 32002 17556 32060
rect 17500 31950 17502 32002
rect 17554 31950 17556 32002
rect 17500 31444 17556 31950
rect 17836 31780 17892 31790
rect 17836 31686 17892 31724
rect 18060 31780 18116 31790
rect 18172 31780 18228 33068
rect 18060 31778 18228 31780
rect 18060 31726 18062 31778
rect 18114 31726 18228 31778
rect 18060 31724 18228 31726
rect 18060 31714 18116 31724
rect 17500 31378 17556 31388
rect 17500 31220 17556 31230
rect 17276 31218 17556 31220
rect 17276 31166 17502 31218
rect 17554 31166 17556 31218
rect 17276 31164 17556 31166
rect 17500 31154 17556 31164
rect 17836 31108 17892 31118
rect 17836 31014 17892 31052
rect 17948 29540 18004 29550
rect 17948 29538 18116 29540
rect 17948 29486 17950 29538
rect 18002 29486 18116 29538
rect 17948 29484 18116 29486
rect 17948 29474 18004 29484
rect 17388 29426 17444 29438
rect 17388 29374 17390 29426
rect 17442 29374 17444 29426
rect 17276 28980 17332 28990
rect 17276 28642 17332 28924
rect 17388 28756 17444 29374
rect 17388 28690 17444 28700
rect 17724 29426 17780 29438
rect 17724 29374 17726 29426
rect 17778 29374 17780 29426
rect 17276 28590 17278 28642
rect 17330 28590 17332 28642
rect 17276 28532 17332 28590
rect 17276 28466 17332 28476
rect 16940 27022 16942 27074
rect 16994 27022 16996 27074
rect 16940 26964 16996 27022
rect 16940 26898 16996 26908
rect 17052 28364 17220 28420
rect 16716 26684 16884 26740
rect 17052 26740 17108 28364
rect 17500 27860 17556 27870
rect 16716 26292 16772 26684
rect 17052 26674 17108 26684
rect 17164 27858 17556 27860
rect 17164 27806 17502 27858
rect 17554 27806 17556 27858
rect 17164 27804 17556 27806
rect 16828 26516 16884 26526
rect 17164 26516 17220 27804
rect 17500 27794 17556 27804
rect 17612 27074 17668 27086
rect 17612 27022 17614 27074
rect 17666 27022 17668 27074
rect 16828 26514 17220 26516
rect 16828 26462 16830 26514
rect 16882 26462 17220 26514
rect 16828 26460 17220 26462
rect 17276 26628 17332 26638
rect 16828 26450 16884 26460
rect 17276 26404 17332 26572
rect 16940 26348 17332 26404
rect 16716 26236 16884 26292
rect 16156 24894 16158 24946
rect 16210 24894 16212 24946
rect 16156 24882 16212 24894
rect 16380 25116 16660 25172
rect 16828 25172 16884 26236
rect 15820 24722 15988 24724
rect 15820 24670 15822 24722
rect 15874 24670 15988 24722
rect 15820 24668 15988 24670
rect 15820 24658 15876 24668
rect 15596 24558 15598 24610
rect 15650 24558 15652 24610
rect 15596 24500 15652 24558
rect 15372 24444 15596 24500
rect 15372 24162 15428 24444
rect 15596 24434 15652 24444
rect 15372 24110 15374 24162
rect 15426 24110 15428 24162
rect 15372 24098 15428 24110
rect 15372 23266 15428 23278
rect 16044 23268 16100 23278
rect 15372 23214 15374 23266
rect 15426 23214 15428 23266
rect 15372 22932 15428 23214
rect 15372 22372 15428 22876
rect 15932 23266 16100 23268
rect 15932 23214 16046 23266
rect 16098 23214 16100 23266
rect 15932 23212 16100 23214
rect 15820 22596 15876 22606
rect 15708 22372 15764 22382
rect 15372 22370 15764 22372
rect 15372 22318 15374 22370
rect 15426 22318 15710 22370
rect 15762 22318 15764 22370
rect 15372 22316 15764 22318
rect 15372 22306 15428 22316
rect 15708 22306 15764 22316
rect 15260 22194 15316 22204
rect 15820 22146 15876 22540
rect 15820 22094 15822 22146
rect 15874 22094 15876 22146
rect 15820 21924 15876 22094
rect 15484 21868 15876 21924
rect 15484 21586 15540 21868
rect 15596 21700 15652 21710
rect 15932 21700 15988 23212
rect 16044 23202 16100 23212
rect 16156 23154 16212 23166
rect 16156 23102 16158 23154
rect 16210 23102 16212 23154
rect 15596 21606 15652 21644
rect 15708 21644 15988 21700
rect 16044 22930 16100 22942
rect 16044 22878 16046 22930
rect 16098 22878 16100 22930
rect 15484 21534 15486 21586
rect 15538 21534 15540 21586
rect 15484 21140 15540 21534
rect 15596 21140 15652 21150
rect 15484 21084 15596 21140
rect 15596 21074 15652 21084
rect 14700 20972 14812 21028
rect 14588 20804 14644 20814
rect 14700 20804 14756 20972
rect 14812 20962 14868 20972
rect 14924 20972 15092 21028
rect 14588 20802 14756 20804
rect 14588 20750 14590 20802
rect 14642 20750 14756 20802
rect 14588 20748 14756 20750
rect 14588 20738 14644 20748
rect 14476 20692 14532 20702
rect 14476 20598 14532 20636
rect 14924 20692 14980 20972
rect 15596 20916 15652 20926
rect 15708 20916 15764 21644
rect 15932 21364 15988 21374
rect 15596 20914 15764 20916
rect 15596 20862 15598 20914
rect 15650 20862 15764 20914
rect 15596 20860 15764 20862
rect 15820 21308 15932 21364
rect 15596 20850 15652 20860
rect 14924 20626 14980 20636
rect 15036 20804 15092 20814
rect 14364 18386 14420 18396
rect 14476 20356 14532 20366
rect 14364 17780 14420 17790
rect 14364 17686 14420 17724
rect 13916 17054 13918 17106
rect 13970 17054 13972 17106
rect 13916 17042 13972 17054
rect 14140 17554 14196 17566
rect 14140 17502 14142 17554
rect 14194 17502 14196 17554
rect 13804 16996 13860 17006
rect 13692 16940 13804 16996
rect 13244 16146 13300 16156
rect 13580 16884 13636 16894
rect 13580 16210 13636 16828
rect 13580 16158 13582 16210
rect 13634 16158 13636 16210
rect 13580 16146 13636 16158
rect 13468 16100 13524 16110
rect 13468 16006 13524 16044
rect 13692 15988 13748 16940
rect 13804 16930 13860 16940
rect 14140 16884 14196 17502
rect 14140 16818 14196 16828
rect 14252 16996 14308 17006
rect 14252 16882 14308 16940
rect 14252 16830 14254 16882
rect 14306 16830 14308 16882
rect 14252 16818 14308 16830
rect 14476 16994 14532 20300
rect 14700 20132 14756 20142
rect 14700 20018 14756 20076
rect 14700 19966 14702 20018
rect 14754 19966 14756 20018
rect 14700 19954 14756 19966
rect 14700 19796 14756 19806
rect 14588 19460 14644 19470
rect 14588 19234 14644 19404
rect 14588 19182 14590 19234
rect 14642 19182 14644 19234
rect 14588 19170 14644 19182
rect 14700 17890 14756 19740
rect 14924 19124 14980 19134
rect 15036 19124 15092 20748
rect 15484 20804 15540 20814
rect 14924 19122 15092 19124
rect 14924 19070 14926 19122
rect 14978 19070 15092 19122
rect 14924 19068 15092 19070
rect 15148 20690 15204 20702
rect 15148 20638 15150 20690
rect 15202 20638 15204 20690
rect 14924 19058 14980 19068
rect 15036 18676 15092 18686
rect 15036 18338 15092 18620
rect 15036 18286 15038 18338
rect 15090 18286 15092 18338
rect 15036 18274 15092 18286
rect 15148 18452 15204 20638
rect 15372 20692 15428 20702
rect 15372 20598 15428 20636
rect 15484 20690 15540 20748
rect 15484 20638 15486 20690
rect 15538 20638 15540 20690
rect 15484 20626 15540 20638
rect 15708 20692 15764 20702
rect 15820 20692 15876 21308
rect 15932 21298 15988 21308
rect 16044 20804 16100 22878
rect 16156 22372 16212 23102
rect 16156 22306 16212 22316
rect 16268 21364 16324 21374
rect 16268 21270 16324 21308
rect 16044 20738 16100 20748
rect 15708 20690 15876 20692
rect 15708 20638 15710 20690
rect 15762 20638 15876 20690
rect 15708 20636 15876 20638
rect 15708 20626 15764 20636
rect 15596 20580 15652 20590
rect 15484 20132 15540 20142
rect 15372 20020 15428 20030
rect 15372 19926 15428 19964
rect 15372 19124 15428 19134
rect 14700 17838 14702 17890
rect 14754 17838 14756 17890
rect 14700 17826 14756 17838
rect 15148 17556 15204 18396
rect 15260 19122 15428 19124
rect 15260 19070 15374 19122
rect 15426 19070 15428 19122
rect 15260 19068 15428 19070
rect 15260 18228 15316 19068
rect 15372 19058 15428 19068
rect 15484 19122 15540 20076
rect 15596 20020 15652 20524
rect 16380 20356 16436 25116
rect 16828 25106 16884 25116
rect 16604 24948 16660 24958
rect 16604 24854 16660 24892
rect 16828 24724 16884 24762
rect 16828 24658 16884 24668
rect 16604 24612 16660 24622
rect 16492 24498 16548 24510
rect 16492 24446 16494 24498
rect 16546 24446 16548 24498
rect 16492 23716 16548 24446
rect 16492 23650 16548 23660
rect 16604 23154 16660 24556
rect 16716 23716 16772 23726
rect 16716 23380 16772 23660
rect 16716 23314 16772 23324
rect 16604 23102 16606 23154
rect 16658 23102 16660 23154
rect 16604 23090 16660 23102
rect 16828 23266 16884 23278
rect 16828 23214 16830 23266
rect 16882 23214 16884 23266
rect 16828 22260 16884 23214
rect 16940 22932 16996 26348
rect 17612 26292 17668 27022
rect 17724 26908 17780 29374
rect 17948 29314 18004 29326
rect 17948 29262 17950 29314
rect 18002 29262 18004 29314
rect 17724 26852 17892 26908
rect 17612 26226 17668 26236
rect 17724 26516 17780 26526
rect 17052 26180 17108 26190
rect 17052 25508 17108 26124
rect 17052 25414 17108 25452
rect 17612 26068 17668 26078
rect 17724 26068 17780 26460
rect 17668 26012 17780 26068
rect 17612 25506 17668 26012
rect 17612 25454 17614 25506
rect 17666 25454 17668 25506
rect 17612 25442 17668 25454
rect 17724 25620 17780 25630
rect 16940 22866 16996 22876
rect 17164 25282 17220 25294
rect 17164 25230 17166 25282
rect 17218 25230 17220 25282
rect 16940 22484 16996 22494
rect 16996 22428 17108 22484
rect 16940 22418 16996 22428
rect 16828 22194 16884 22204
rect 16940 22148 16996 22158
rect 16940 22054 16996 22092
rect 16604 21364 16660 21374
rect 16604 21362 16772 21364
rect 16604 21310 16606 21362
rect 16658 21310 16772 21362
rect 16604 21308 16772 21310
rect 16604 21298 16660 21308
rect 15596 19954 15652 19964
rect 16156 20300 16436 20356
rect 16492 21140 16548 21150
rect 16492 20580 16548 21084
rect 15708 19236 15764 19246
rect 15708 19142 15764 19180
rect 15484 19070 15486 19122
rect 15538 19070 15540 19122
rect 15484 18676 15540 19070
rect 15932 19012 15988 19022
rect 15484 18610 15540 18620
rect 15596 19010 15988 19012
rect 15596 18958 15934 19010
rect 15986 18958 15988 19010
rect 15596 18956 15988 18958
rect 15372 18452 15428 18462
rect 15596 18452 15652 18956
rect 15932 18946 15988 18956
rect 16044 18562 16100 18574
rect 16044 18510 16046 18562
rect 16098 18510 16100 18562
rect 15372 18450 15764 18452
rect 15372 18398 15374 18450
rect 15426 18398 15764 18450
rect 15372 18396 15764 18398
rect 15372 18386 15428 18396
rect 15260 18172 15428 18228
rect 15260 17892 15316 17902
rect 15260 17798 15316 17836
rect 15260 17556 15316 17566
rect 15148 17554 15316 17556
rect 15148 17502 15262 17554
rect 15314 17502 15316 17554
rect 15148 17500 15316 17502
rect 15260 17490 15316 17500
rect 15372 17556 15428 18172
rect 15708 17892 15764 18396
rect 16044 18228 16100 18510
rect 16044 18162 16100 18172
rect 15820 17892 15876 17902
rect 15708 17890 15876 17892
rect 15708 17838 15822 17890
rect 15874 17838 15876 17890
rect 15708 17836 15876 17838
rect 15820 17826 15876 17836
rect 15596 17556 15652 17566
rect 15372 17554 15596 17556
rect 15372 17502 15374 17554
rect 15426 17502 15596 17554
rect 15372 17500 15596 17502
rect 15372 17490 15428 17500
rect 15596 17490 15652 17500
rect 15484 17108 15540 17118
rect 15484 17014 15540 17052
rect 16044 17108 16100 17118
rect 14476 16942 14478 16994
rect 14530 16942 14532 16994
rect 14476 16436 14532 16942
rect 14476 16370 14532 16380
rect 14924 16994 14980 17006
rect 14924 16942 14926 16994
rect 14978 16942 14980 16994
rect 13916 16324 13972 16334
rect 13916 16230 13972 16268
rect 14028 16100 14084 16110
rect 14028 16006 14084 16044
rect 14476 16098 14532 16110
rect 14700 16100 14756 16110
rect 14476 16046 14478 16098
rect 14530 16046 14532 16098
rect 13020 15538 13188 15540
rect 13020 15486 13022 15538
rect 13074 15486 13188 15538
rect 13020 15484 13188 15486
rect 13580 15932 13748 15988
rect 13020 15474 13076 15484
rect 12908 15262 12910 15314
rect 12962 15262 12964 15314
rect 12908 15250 12964 15262
rect 13244 15314 13300 15326
rect 13244 15262 13246 15314
rect 13298 15262 13300 15314
rect 13132 15202 13188 15214
rect 13132 15150 13134 15202
rect 13186 15150 13188 15202
rect 13132 13860 13188 15150
rect 13244 15148 13300 15262
rect 13244 15092 13524 15148
rect 13132 13794 13188 13804
rect 13132 12292 13188 12302
rect 13132 12198 13188 12236
rect 13020 12178 13076 12190
rect 13020 12126 13022 12178
rect 13074 12126 13076 12178
rect 12796 11732 12964 11788
rect 12684 11554 12740 11564
rect 12796 11618 12852 11630
rect 12796 11566 12798 11618
rect 12850 11566 12852 11618
rect 12572 11442 12628 11452
rect 12684 11284 12740 11294
rect 12460 11282 12740 11284
rect 12460 11230 12686 11282
rect 12738 11230 12740 11282
rect 12460 11228 12740 11230
rect 12460 10836 12516 10846
rect 12460 10742 12516 10780
rect 12460 10612 12516 10622
rect 12460 10518 12516 10556
rect 12236 10386 12292 10444
rect 12236 10334 12238 10386
rect 12290 10334 12292 10386
rect 12236 10322 12292 10334
rect 12124 10210 12180 10220
rect 12012 9996 12404 10052
rect 11564 8932 11620 9996
rect 12012 9826 12068 9838
rect 12012 9774 12014 9826
rect 12066 9774 12068 9826
rect 11564 8866 11620 8876
rect 11676 9714 11732 9726
rect 11676 9662 11678 9714
rect 11730 9662 11732 9714
rect 11004 8260 11060 8270
rect 11004 8166 11060 8204
rect 11564 8260 11620 8270
rect 10892 8082 10948 8092
rect 10556 6862 10558 6914
rect 10610 6862 10612 6914
rect 10556 6850 10612 6862
rect 10892 7586 10948 7598
rect 10892 7534 10894 7586
rect 10946 7534 10948 7586
rect 10892 6804 10948 7534
rect 10892 6710 10948 6748
rect 10108 6638 10110 6690
rect 10162 6638 10164 6690
rect 10108 6626 10164 6638
rect 11564 6578 11620 8204
rect 11676 7364 11732 9662
rect 12012 9268 12068 9774
rect 12012 9202 12068 9212
rect 11676 7298 11732 7308
rect 11788 9154 11844 9166
rect 11788 9102 11790 9154
rect 11842 9102 11844 9154
rect 11788 8146 11844 9102
rect 11788 8094 11790 8146
rect 11842 8094 11844 8146
rect 11788 6804 11844 8094
rect 11788 6738 11844 6748
rect 12236 8146 12292 8158
rect 12236 8094 12238 8146
rect 12290 8094 12292 8146
rect 12236 7250 12292 8094
rect 12236 7198 12238 7250
rect 12290 7198 12292 7250
rect 11676 6692 11732 6702
rect 11676 6598 11732 6636
rect 12236 6692 12292 7198
rect 12348 6692 12404 9996
rect 12572 8372 12628 8382
rect 12460 8260 12516 8270
rect 12460 8166 12516 8204
rect 12572 7476 12628 8316
rect 12684 8036 12740 11228
rect 12796 10610 12852 11566
rect 12796 10558 12798 10610
rect 12850 10558 12852 10610
rect 12796 10546 12852 10558
rect 12908 11618 12964 11732
rect 12908 11566 12910 11618
rect 12962 11566 12964 11618
rect 12908 10388 12964 11566
rect 13020 11060 13076 12126
rect 13244 12178 13300 12190
rect 13244 12126 13246 12178
rect 13298 12126 13300 12178
rect 13020 10994 13076 11004
rect 13132 11396 13188 11406
rect 13020 10836 13076 10846
rect 13020 10610 13076 10780
rect 13020 10558 13022 10610
rect 13074 10558 13076 10610
rect 13020 10546 13076 10558
rect 12796 10332 12964 10388
rect 13132 10500 13188 11340
rect 13244 11172 13300 12126
rect 13356 11396 13412 11406
rect 13356 11302 13412 11340
rect 13244 11106 13300 11116
rect 13244 10948 13300 10958
rect 13244 10834 13300 10892
rect 13244 10782 13246 10834
rect 13298 10782 13300 10834
rect 13244 10770 13300 10782
rect 13468 10834 13524 15092
rect 13580 14756 13636 15932
rect 14476 15764 14532 16046
rect 13580 14662 13636 14700
rect 13692 15708 14532 15764
rect 14588 16098 14756 16100
rect 14588 16046 14702 16098
rect 14754 16046 14756 16098
rect 14588 16044 14756 16046
rect 13692 14642 13748 15708
rect 14588 15652 14644 16044
rect 14700 16034 14756 16044
rect 13916 15596 14644 15652
rect 14812 15874 14868 15886
rect 14812 15822 14814 15874
rect 14866 15822 14868 15874
rect 13916 15538 13972 15596
rect 13916 15486 13918 15538
rect 13970 15486 13972 15538
rect 13916 15474 13972 15486
rect 13804 15428 13860 15438
rect 13804 15148 13860 15372
rect 14812 15426 14868 15822
rect 14812 15374 14814 15426
rect 14866 15374 14868 15426
rect 14812 15362 14868 15374
rect 14924 15204 14980 16942
rect 15484 16884 15540 16894
rect 15932 16884 15988 16894
rect 15484 16790 15540 16828
rect 15708 16882 15988 16884
rect 15708 16830 15934 16882
rect 15986 16830 15988 16882
rect 15708 16828 15988 16830
rect 15372 16772 15428 16782
rect 15372 16322 15428 16716
rect 15372 16270 15374 16322
rect 15426 16270 15428 16322
rect 15372 16258 15428 16270
rect 15708 16098 15764 16828
rect 15932 16818 15988 16828
rect 15708 16046 15710 16098
rect 15762 16046 15764 16098
rect 15708 15428 15764 16046
rect 15708 15362 15764 15372
rect 15820 16658 15876 16670
rect 15820 16606 15822 16658
rect 15874 16606 15876 16658
rect 14812 15148 14980 15204
rect 13804 15092 13972 15148
rect 13692 14590 13694 14642
rect 13746 14590 13748 14642
rect 13692 14578 13748 14590
rect 13804 14980 13860 14990
rect 13804 14420 13860 14924
rect 13804 14326 13860 14364
rect 13916 14308 13972 15092
rect 14028 15090 14084 15102
rect 14028 15038 14030 15090
rect 14082 15038 14084 15090
rect 14028 14756 14084 15038
rect 14812 14980 14868 15148
rect 14588 14924 14868 14980
rect 14588 14756 14644 14924
rect 14028 14700 14644 14756
rect 14700 14756 14756 14766
rect 14252 14308 14308 14318
rect 13916 14306 14308 14308
rect 13916 14254 14254 14306
rect 14306 14254 14308 14306
rect 13916 14252 14308 14254
rect 13692 13524 13748 13534
rect 13580 12292 13636 12302
rect 13580 12198 13636 12236
rect 13468 10782 13470 10834
rect 13522 10782 13524 10834
rect 12796 9940 12852 10332
rect 13020 10276 13076 10286
rect 12796 8428 12852 9884
rect 12908 10220 13020 10276
rect 12908 9154 12964 10220
rect 13020 10210 13076 10220
rect 13020 9268 13076 9278
rect 13020 9174 13076 9212
rect 13132 9266 13188 10444
rect 13132 9214 13134 9266
rect 13186 9214 13188 9266
rect 13132 9202 13188 9214
rect 13356 10498 13412 10510
rect 13356 10446 13358 10498
rect 13410 10446 13412 10498
rect 12908 9102 12910 9154
rect 12962 9102 12964 9154
rect 12908 9090 12964 9102
rect 12796 8372 12964 8428
rect 12796 8260 12852 8270
rect 12796 8166 12852 8204
rect 12684 7980 12852 8036
rect 12684 7476 12740 7486
rect 12572 7474 12740 7476
rect 12572 7422 12686 7474
rect 12738 7422 12740 7474
rect 12572 7420 12740 7422
rect 12460 6692 12516 6702
rect 12348 6690 12516 6692
rect 12348 6638 12462 6690
rect 12514 6638 12516 6690
rect 12348 6636 12516 6638
rect 12236 6626 12292 6636
rect 12460 6626 12516 6636
rect 11564 6526 11566 6578
rect 11618 6526 11620 6578
rect 11564 6514 11620 6526
rect 12460 6132 12516 6142
rect 12572 6132 12628 7420
rect 12684 7410 12740 7420
rect 12796 6580 12852 7980
rect 12796 6514 12852 6524
rect 12908 6468 12964 8372
rect 13356 7588 13412 10446
rect 13468 7924 13524 10782
rect 13580 11060 13636 11070
rect 13580 10388 13636 11004
rect 13692 10836 13748 13468
rect 14252 12964 14308 14252
rect 14364 13524 14420 14700
rect 14476 14532 14532 14542
rect 14476 13634 14532 14476
rect 14588 14306 14644 14318
rect 14588 14254 14590 14306
rect 14642 14254 14644 14306
rect 14588 13748 14644 14254
rect 14588 13682 14644 13692
rect 14476 13582 14478 13634
rect 14530 13582 14532 13634
rect 14476 13570 14532 13582
rect 14364 13458 14420 13468
rect 14252 12898 14308 12908
rect 14028 12852 14084 12862
rect 14028 12758 14084 12796
rect 13804 12180 13860 12190
rect 13804 12086 13860 12124
rect 14252 12178 14308 12190
rect 14252 12126 14254 12178
rect 14306 12126 14308 12178
rect 14028 12066 14084 12078
rect 14028 12014 14030 12066
rect 14082 12014 14084 12066
rect 14028 11620 14084 12014
rect 14028 11554 14084 11564
rect 13692 10770 13748 10780
rect 13916 11396 13972 11406
rect 13580 9042 13636 10332
rect 13916 10498 13972 11340
rect 13916 10446 13918 10498
rect 13970 10446 13972 10498
rect 13804 10164 13860 10174
rect 13916 10164 13972 10446
rect 13860 10108 13972 10164
rect 14140 10386 14196 10398
rect 14140 10334 14142 10386
rect 14194 10334 14196 10386
rect 13804 9938 13860 10108
rect 13804 9886 13806 9938
rect 13858 9886 13860 9938
rect 13804 9874 13860 9886
rect 14028 9828 14084 9838
rect 14140 9828 14196 10334
rect 14028 9826 14196 9828
rect 14028 9774 14030 9826
rect 14082 9774 14196 9826
rect 14028 9772 14196 9774
rect 14028 9762 14084 9772
rect 13580 8990 13582 9042
rect 13634 8990 13636 9042
rect 13580 8978 13636 8990
rect 14140 9042 14196 9772
rect 14252 9268 14308 12126
rect 14588 12180 14644 12190
rect 14588 12086 14644 12124
rect 14476 11954 14532 11966
rect 14476 11902 14478 11954
rect 14530 11902 14532 11954
rect 14476 10612 14532 11902
rect 14476 10546 14532 10556
rect 14476 10386 14532 10398
rect 14476 10334 14478 10386
rect 14530 10334 14532 10386
rect 14364 9604 14420 9614
rect 14364 9510 14420 9548
rect 14252 9202 14308 9212
rect 14140 8990 14142 9042
rect 14194 8990 14196 9042
rect 14140 8372 14196 8990
rect 14476 9042 14532 10334
rect 14700 10164 14756 14700
rect 14924 14532 14980 14542
rect 14924 14438 14980 14476
rect 14812 14420 14868 14430
rect 15596 14420 15652 14430
rect 14812 11788 14868 14364
rect 15372 14364 15596 14420
rect 15260 14308 15316 14318
rect 15260 14214 15316 14252
rect 15036 13748 15092 13758
rect 15036 13654 15092 13692
rect 15260 12292 15316 12302
rect 15260 12198 15316 12236
rect 15036 12180 15092 12190
rect 15036 12086 15092 12124
rect 14812 11732 14980 11788
rect 14476 8990 14478 9042
rect 14530 8990 14532 9042
rect 14476 8978 14532 8990
rect 14588 10108 14756 10164
rect 14140 8306 14196 8316
rect 14140 8036 14196 8046
rect 14140 8034 14420 8036
rect 14140 7982 14142 8034
rect 14194 7982 14420 8034
rect 14140 7980 14420 7982
rect 14140 7970 14196 7980
rect 13468 7868 13636 7924
rect 13468 7588 13524 7598
rect 13356 7586 13524 7588
rect 13356 7534 13470 7586
rect 13522 7534 13524 7586
rect 13356 7532 13524 7534
rect 13468 7522 13524 7532
rect 13580 7028 13636 7868
rect 13468 6972 13748 7028
rect 13468 6916 13524 6972
rect 13356 6860 13524 6916
rect 13020 6692 13076 6702
rect 13356 6692 13412 6860
rect 13580 6804 13636 6814
rect 13020 6690 13412 6692
rect 13020 6638 13022 6690
rect 13074 6638 13412 6690
rect 13020 6636 13412 6638
rect 13468 6692 13524 6702
rect 13020 6626 13076 6636
rect 13468 6598 13524 6636
rect 12908 6412 13300 6468
rect 12460 6130 12628 6132
rect 12460 6078 12462 6130
rect 12514 6078 12628 6130
rect 12460 6076 12628 6078
rect 13244 6130 13300 6412
rect 13244 6078 13246 6130
rect 13298 6078 13300 6130
rect 12460 6066 12516 6076
rect 13244 6066 13300 6078
rect 13468 6132 13524 6142
rect 13580 6132 13636 6748
rect 13468 6130 13636 6132
rect 13468 6078 13470 6130
rect 13522 6078 13636 6130
rect 13468 6076 13636 6078
rect 13468 6066 13524 6076
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 13692 5236 13748 6972
rect 13804 6580 13860 6590
rect 14364 6580 14420 7980
rect 13804 6486 13860 6524
rect 13916 6578 14420 6580
rect 13916 6526 14366 6578
rect 14418 6526 14420 6578
rect 13916 6524 14420 6526
rect 13804 6020 13860 6030
rect 13916 6020 13972 6524
rect 14364 6514 14420 6524
rect 14588 6692 14644 10108
rect 14700 9940 14756 9950
rect 14700 9826 14756 9884
rect 14700 9774 14702 9826
rect 14754 9774 14756 9826
rect 14700 9762 14756 9774
rect 14812 9602 14868 9614
rect 14812 9550 14814 9602
rect 14866 9550 14868 9602
rect 14812 9156 14868 9550
rect 14812 9090 14868 9100
rect 14476 6132 14532 6142
rect 14588 6132 14644 6636
rect 14700 7028 14756 7038
rect 14700 6690 14756 6972
rect 14700 6638 14702 6690
rect 14754 6638 14756 6690
rect 14700 6626 14756 6638
rect 14476 6130 14644 6132
rect 14476 6078 14478 6130
rect 14530 6078 14644 6130
rect 14476 6076 14644 6078
rect 14924 6580 14980 11732
rect 15148 11620 15204 11630
rect 15148 11282 15204 11564
rect 15148 11230 15150 11282
rect 15202 11230 15204 11282
rect 15148 11218 15204 11230
rect 15148 10724 15204 10734
rect 15036 9828 15092 9838
rect 15036 8428 15092 9772
rect 15148 9154 15204 10668
rect 15148 9102 15150 9154
rect 15202 9102 15204 9154
rect 15148 9090 15204 9102
rect 15260 10610 15316 10622
rect 15260 10558 15262 10610
rect 15314 10558 15316 10610
rect 15260 9714 15316 10558
rect 15372 9828 15428 14364
rect 15596 14326 15652 14364
rect 15820 13860 15876 16606
rect 15932 16212 15988 16222
rect 15932 16098 15988 16156
rect 15932 16046 15934 16098
rect 15986 16046 15988 16098
rect 15932 16034 15988 16046
rect 16044 14420 16100 17052
rect 16044 14354 16100 14364
rect 16156 14084 16212 20300
rect 16268 20020 16324 20030
rect 16268 18228 16324 19964
rect 16492 20018 16548 20524
rect 16492 19966 16494 20018
rect 16546 19966 16548 20018
rect 16492 19954 16548 19966
rect 16604 20692 16660 20702
rect 16604 19794 16660 20636
rect 16716 20020 16772 21308
rect 16716 19954 16772 19964
rect 16828 21028 16884 21038
rect 16828 19796 16884 20972
rect 16604 19742 16606 19794
rect 16658 19742 16660 19794
rect 16604 19730 16660 19742
rect 16716 19740 16884 19796
rect 16492 19122 16548 19134
rect 16492 19070 16494 19122
rect 16546 19070 16548 19122
rect 16492 18452 16548 19070
rect 16492 18386 16548 18396
rect 16604 18562 16660 18574
rect 16604 18510 16606 18562
rect 16658 18510 16660 18562
rect 16268 18162 16324 18172
rect 16604 17668 16660 18510
rect 16716 18450 16772 19740
rect 16940 19348 16996 19358
rect 16940 19254 16996 19292
rect 16828 19236 16884 19246
rect 16828 19142 16884 19180
rect 16716 18398 16718 18450
rect 16770 18398 16772 18450
rect 16716 18386 16772 18398
rect 16940 18340 16996 18350
rect 16940 18246 16996 18284
rect 16604 17602 16660 17612
rect 16492 17556 16548 17566
rect 17052 17556 17108 22428
rect 17164 20244 17220 25230
rect 17388 25282 17444 25294
rect 17388 25230 17390 25282
rect 17442 25230 17444 25282
rect 17276 23826 17332 23838
rect 17276 23774 17278 23826
rect 17330 23774 17332 23826
rect 17276 23156 17332 23774
rect 17388 23492 17444 25230
rect 17724 24948 17780 25564
rect 17836 25060 17892 26852
rect 17948 26402 18004 29262
rect 18060 28532 18116 29484
rect 18060 28466 18116 28476
rect 18172 29426 18228 29438
rect 18172 29374 18174 29426
rect 18226 29374 18228 29426
rect 18172 28420 18228 29374
rect 18172 28354 18228 28364
rect 18284 28196 18340 33852
rect 18508 33796 18564 34190
rect 18508 33730 18564 33740
rect 18620 33346 18676 34860
rect 18620 33294 18622 33346
rect 18674 33294 18676 33346
rect 18620 33282 18676 33294
rect 18732 34130 18788 34142
rect 18732 34078 18734 34130
rect 18786 34078 18788 34130
rect 18508 33234 18564 33246
rect 18508 33182 18510 33234
rect 18562 33182 18564 33234
rect 18508 32564 18564 33182
rect 18508 32498 18564 32508
rect 18732 32452 18788 34078
rect 19068 33460 19124 33498
rect 19068 33394 19124 33404
rect 19068 33236 19124 33246
rect 19068 33142 19124 33180
rect 18732 32386 18788 32396
rect 19068 32562 19124 32574
rect 19068 32510 19070 32562
rect 19122 32510 19124 32562
rect 19068 32340 19124 32510
rect 18508 31778 18564 31790
rect 18508 31726 18510 31778
rect 18562 31726 18564 31778
rect 18508 31668 18564 31726
rect 18508 30996 18564 31612
rect 18732 31668 18788 31678
rect 19068 31668 19124 32284
rect 18732 31666 19124 31668
rect 18732 31614 18734 31666
rect 18786 31614 19124 31666
rect 18732 31612 19124 31614
rect 18732 31220 18788 31612
rect 18732 31154 18788 31164
rect 18844 31220 18900 31230
rect 19068 31220 19124 31230
rect 18844 31218 19068 31220
rect 18844 31166 18846 31218
rect 18898 31166 19068 31218
rect 18844 31164 19068 31166
rect 18844 31154 18900 31164
rect 19068 31154 19124 31164
rect 18508 30930 18564 30940
rect 18956 30098 19012 30110
rect 18956 30046 18958 30098
rect 19010 30046 19012 30098
rect 18732 29428 18788 29438
rect 18732 29426 18900 29428
rect 18732 29374 18734 29426
rect 18786 29374 18900 29426
rect 18732 29372 18900 29374
rect 18732 29362 18788 29372
rect 18620 28756 18676 28766
rect 18172 28140 18340 28196
rect 18508 28700 18620 28756
rect 18060 28084 18116 28094
rect 18060 27186 18116 28028
rect 18060 27134 18062 27186
rect 18114 27134 18116 27186
rect 18060 27122 18116 27134
rect 18172 26908 18228 28140
rect 17948 26350 17950 26402
rect 18002 26350 18004 26402
rect 17948 26338 18004 26350
rect 18060 26852 18228 26908
rect 18284 27746 18340 27758
rect 18284 27694 18286 27746
rect 18338 27694 18340 27746
rect 17948 25732 18004 25742
rect 17948 25618 18004 25676
rect 17948 25566 17950 25618
rect 18002 25566 18004 25618
rect 17948 25554 18004 25566
rect 18060 25396 18116 26852
rect 18284 25620 18340 27694
rect 18508 26908 18564 28700
rect 18620 28690 18676 28700
rect 18844 28418 18900 29372
rect 18956 28754 19012 30046
rect 18956 28702 18958 28754
rect 19010 28702 19012 28754
rect 18956 28690 19012 28702
rect 19180 29540 19236 35420
rect 19292 33796 19348 33806
rect 19292 33346 19348 33740
rect 19292 33294 19294 33346
rect 19346 33294 19348 33346
rect 19292 32562 19348 33294
rect 19292 32510 19294 32562
rect 19346 32510 19348 32562
rect 19292 32498 19348 32510
rect 18844 28366 18846 28418
rect 18898 28366 18900 28418
rect 18620 27972 18676 27982
rect 18844 27972 18900 28366
rect 19068 28644 19124 28654
rect 19068 28196 19124 28588
rect 18676 27916 18900 27972
rect 18956 28140 19124 28196
rect 18620 27858 18676 27916
rect 18620 27806 18622 27858
rect 18674 27806 18676 27858
rect 18620 27794 18676 27806
rect 18732 27748 18788 27758
rect 18788 27692 18900 27748
rect 18732 27682 18788 27692
rect 18844 27076 18900 27692
rect 18396 26852 18564 26908
rect 18732 26964 18788 27002
rect 18732 26898 18788 26908
rect 18396 26516 18452 26852
rect 18396 26450 18452 26460
rect 18732 25956 18788 25966
rect 18620 25900 18732 25956
rect 18060 25330 18116 25340
rect 18172 25564 18340 25620
rect 18508 25620 18564 25630
rect 18060 25172 18116 25182
rect 17836 25004 18004 25060
rect 17724 24892 17892 24948
rect 17836 24834 17892 24892
rect 17836 24782 17838 24834
rect 17890 24782 17892 24834
rect 17836 24770 17892 24782
rect 17500 24724 17556 24734
rect 17500 24630 17556 24668
rect 17388 23426 17444 23436
rect 17612 24610 17668 24622
rect 17612 24558 17614 24610
rect 17666 24558 17668 24610
rect 17612 23378 17668 24558
rect 17612 23326 17614 23378
rect 17666 23326 17668 23378
rect 17612 23314 17668 23326
rect 17724 24164 17780 24174
rect 17948 24164 18004 25004
rect 18060 24834 18116 25116
rect 18060 24782 18062 24834
rect 18114 24782 18116 24834
rect 18060 24770 18116 24782
rect 18060 24164 18116 24174
rect 17948 24162 18116 24164
rect 17948 24110 18062 24162
rect 18114 24110 18116 24162
rect 17948 24108 18116 24110
rect 17276 23100 17444 23156
rect 17388 22932 17444 23100
rect 17500 22932 17556 22942
rect 17388 22930 17556 22932
rect 17388 22878 17502 22930
rect 17554 22878 17556 22930
rect 17388 22876 17556 22878
rect 17500 22866 17556 22876
rect 17276 22484 17332 22494
rect 17276 22258 17332 22428
rect 17276 22206 17278 22258
rect 17330 22206 17332 22258
rect 17276 22194 17332 22206
rect 17612 22370 17668 22382
rect 17612 22318 17614 22370
rect 17666 22318 17668 22370
rect 17612 22260 17668 22318
rect 17612 22194 17668 22204
rect 17724 21810 17780 24108
rect 18060 24098 18116 24108
rect 18172 23940 18228 25564
rect 18396 25508 18452 25518
rect 18284 25452 18396 25508
rect 18284 25394 18340 25452
rect 18396 25442 18452 25452
rect 18508 25506 18564 25564
rect 18508 25454 18510 25506
rect 18562 25454 18564 25506
rect 18508 25442 18564 25454
rect 18284 25342 18286 25394
rect 18338 25342 18340 25394
rect 18284 25330 18340 25342
rect 18508 25282 18564 25294
rect 18508 25230 18510 25282
rect 18562 25230 18564 25282
rect 18396 25172 18452 25182
rect 18396 24722 18452 25116
rect 18396 24670 18398 24722
rect 18450 24670 18452 24722
rect 18396 24658 18452 24670
rect 18396 23940 18452 23950
rect 17948 23884 18228 23940
rect 18284 23938 18452 23940
rect 18284 23886 18398 23938
rect 18450 23886 18452 23938
rect 18284 23884 18452 23886
rect 17836 23380 17892 23390
rect 17836 23266 17892 23324
rect 17836 23214 17838 23266
rect 17890 23214 17892 23266
rect 17836 23202 17892 23214
rect 17948 22372 18004 23884
rect 18284 23604 18340 23884
rect 18396 23874 18452 23884
rect 18060 23548 18340 23604
rect 18060 23268 18116 23548
rect 18172 23380 18228 23390
rect 18172 23378 18452 23380
rect 18172 23326 18174 23378
rect 18226 23326 18452 23378
rect 18172 23324 18452 23326
rect 18172 23314 18228 23324
rect 18060 23202 18116 23212
rect 18284 23156 18340 23166
rect 18284 23062 18340 23100
rect 17724 21758 17726 21810
rect 17778 21758 17780 21810
rect 17724 21746 17780 21758
rect 17836 22316 18004 22372
rect 18060 22932 18116 22942
rect 17612 21700 17668 21710
rect 17388 21586 17444 21598
rect 17388 21534 17390 21586
rect 17442 21534 17444 21586
rect 17388 21028 17444 21534
rect 17388 20934 17444 20972
rect 17276 20916 17332 20926
rect 17276 20802 17332 20860
rect 17276 20750 17278 20802
rect 17330 20750 17332 20802
rect 17276 20468 17332 20750
rect 17276 20402 17332 20412
rect 17164 20188 17332 20244
rect 16492 17108 16548 17500
rect 16716 17554 17108 17556
rect 16716 17502 17054 17554
rect 17106 17502 17108 17554
rect 16716 17500 17108 17502
rect 16604 17108 16660 17118
rect 16492 17106 16660 17108
rect 16492 17054 16606 17106
rect 16658 17054 16660 17106
rect 16492 17052 16660 17054
rect 16604 17042 16660 17052
rect 16268 16996 16324 17006
rect 16268 16902 16324 16940
rect 16716 16996 16772 17500
rect 17052 17490 17108 17500
rect 16716 16902 16772 16940
rect 16492 16212 16548 16222
rect 16380 15986 16436 15998
rect 16380 15934 16382 15986
rect 16434 15934 16436 15986
rect 16268 15874 16324 15886
rect 16268 15822 16270 15874
rect 16322 15822 16324 15874
rect 16268 15428 16324 15822
rect 16268 14530 16324 15372
rect 16268 14478 16270 14530
rect 16322 14478 16324 14530
rect 16268 14466 16324 14478
rect 15820 13794 15876 13804
rect 16044 14028 16212 14084
rect 16268 14308 16324 14318
rect 15596 13636 15652 13646
rect 15484 13188 15540 13198
rect 15484 12180 15540 13132
rect 15596 13186 15652 13580
rect 15596 13134 15598 13186
rect 15650 13134 15652 13186
rect 15596 12404 15652 13134
rect 15596 12338 15652 12348
rect 15932 12290 15988 12302
rect 15932 12238 15934 12290
rect 15986 12238 15988 12290
rect 15596 12180 15652 12190
rect 15484 12178 15652 12180
rect 15484 12126 15598 12178
rect 15650 12126 15652 12178
rect 15484 12124 15652 12126
rect 15484 10610 15540 10622
rect 15484 10558 15486 10610
rect 15538 10558 15540 10610
rect 15484 10052 15540 10558
rect 15484 9986 15540 9996
rect 15372 9772 15540 9828
rect 15260 9662 15262 9714
rect 15314 9662 15316 9714
rect 15260 8708 15316 9662
rect 15260 8642 15316 8652
rect 15036 8372 15204 8428
rect 14924 6130 14980 6524
rect 14924 6078 14926 6130
rect 14978 6078 14980 6130
rect 14476 6066 14532 6076
rect 14924 6066 14980 6078
rect 13804 6018 13916 6020
rect 13804 5966 13806 6018
rect 13858 5966 13916 6018
rect 13804 5964 13916 5966
rect 13804 5954 13860 5964
rect 13916 5926 13972 5964
rect 13804 5236 13860 5246
rect 13692 5234 13860 5236
rect 13692 5182 13806 5234
rect 13858 5182 13860 5234
rect 13692 5180 13860 5182
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 7644 3332 7700 3342
rect 7420 3330 7700 3332
rect 7420 3278 7646 3330
rect 7698 3278 7700 3330
rect 7420 3276 7700 3278
rect 7420 800 7476 3276
rect 7644 3266 7700 3276
rect 13804 2996 13860 5180
rect 15148 5124 15204 8372
rect 15260 8372 15316 8382
rect 15260 8034 15316 8316
rect 15260 7982 15262 8034
rect 15314 7982 15316 8034
rect 15260 7476 15316 7982
rect 15260 7410 15316 7420
rect 15372 6580 15428 6590
rect 15372 6486 15428 6524
rect 15372 6132 15428 6142
rect 15484 6132 15540 9772
rect 15596 8428 15652 12124
rect 15932 11956 15988 12238
rect 16044 11956 16100 14028
rect 16268 13858 16324 14252
rect 16268 13806 16270 13858
rect 16322 13806 16324 13858
rect 16268 13794 16324 13806
rect 16380 13748 16436 15934
rect 16492 15540 16548 16156
rect 16492 15538 17220 15540
rect 16492 15486 16494 15538
rect 16546 15486 17220 15538
rect 16492 15484 17220 15486
rect 16492 15474 16548 15484
rect 16380 13682 16436 13692
rect 16940 13860 16996 13870
rect 16380 13524 16436 13534
rect 16380 12402 16436 13468
rect 16828 13186 16884 13198
rect 16828 13134 16830 13186
rect 16882 13134 16884 13186
rect 16604 12964 16660 12974
rect 16604 12870 16660 12908
rect 16380 12350 16382 12402
rect 16434 12350 16436 12402
rect 16380 12338 16436 12350
rect 16492 12852 16548 12862
rect 16492 12292 16548 12796
rect 16268 12180 16324 12190
rect 16268 12086 16324 12124
rect 16492 12178 16548 12236
rect 16828 12516 16884 13134
rect 16940 12738 16996 13804
rect 17164 13748 17220 15484
rect 17276 14308 17332 20188
rect 17388 20018 17444 20030
rect 17388 19966 17390 20018
rect 17442 19966 17444 20018
rect 17388 17892 17444 19966
rect 17612 18340 17668 21644
rect 17836 21364 17892 22316
rect 17836 20914 17892 21308
rect 17836 20862 17838 20914
rect 17890 20862 17892 20914
rect 17836 20850 17892 20862
rect 17948 20802 18004 20814
rect 17948 20750 17950 20802
rect 18002 20750 18004 20802
rect 17948 20580 18004 20750
rect 17948 20514 18004 20524
rect 18060 19908 18116 22876
rect 18396 22482 18452 23324
rect 18508 23154 18564 25230
rect 18508 23102 18510 23154
rect 18562 23102 18564 23154
rect 18508 23090 18564 23102
rect 18396 22430 18398 22482
rect 18450 22430 18452 22482
rect 18396 22418 18452 22430
rect 18620 21812 18676 25900
rect 18732 25890 18788 25900
rect 18844 25506 18900 27020
rect 18956 25732 19012 28140
rect 19180 27860 19236 29484
rect 19292 30098 19348 30110
rect 19292 30046 19294 30098
rect 19346 30046 19348 30098
rect 19292 29428 19348 30046
rect 19292 29362 19348 29372
rect 19068 27188 19124 27198
rect 19068 27094 19124 27132
rect 18956 25666 19012 25676
rect 18844 25454 18846 25506
rect 18898 25454 18900 25506
rect 18844 24948 18900 25454
rect 19180 25284 19236 27804
rect 19292 27076 19348 27086
rect 19292 26962 19348 27020
rect 19292 26910 19294 26962
rect 19346 26910 19348 26962
rect 19292 26898 19348 26910
rect 19404 25956 19460 35532
rect 19964 35586 20244 35588
rect 19964 35534 19966 35586
rect 20018 35534 20244 35586
rect 19964 35532 20244 35534
rect 19964 35028 20020 35532
rect 19964 34962 20020 34972
rect 20412 34916 20468 37772
rect 20636 37826 20692 37838
rect 20636 37774 20638 37826
rect 20690 37774 20692 37826
rect 20524 36596 20580 36606
rect 20524 36502 20580 36540
rect 20636 36372 20692 37774
rect 20748 37154 20804 37996
rect 21084 38052 21140 39788
rect 21420 39778 21476 39790
rect 21308 39618 21364 39630
rect 21308 39566 21310 39618
rect 21362 39566 21364 39618
rect 21308 39508 21364 39566
rect 21308 39442 21364 39452
rect 21532 38946 21588 38958
rect 21532 38894 21534 38946
rect 21586 38894 21588 38946
rect 21084 37986 21140 37996
rect 21196 38836 21252 38846
rect 21196 38050 21252 38780
rect 21532 38388 21588 38894
rect 22204 38724 22260 40572
rect 22540 40402 22596 41132
rect 22652 41186 22708 41198
rect 22652 41134 22654 41186
rect 22706 41134 22708 41186
rect 22652 40852 22708 41134
rect 22652 40786 22708 40796
rect 22540 40350 22542 40402
rect 22594 40350 22596 40402
rect 22540 40338 22596 40350
rect 22428 40068 22484 40078
rect 22316 39508 22372 39518
rect 22316 39414 22372 39452
rect 22428 39284 22484 40012
rect 22204 38658 22260 38668
rect 22316 39228 22484 39284
rect 22652 39506 22708 39518
rect 22652 39454 22654 39506
rect 22706 39454 22708 39506
rect 21588 38332 21700 38388
rect 21532 38322 21588 38332
rect 21196 37998 21198 38050
rect 21250 37998 21252 38050
rect 21196 37986 21252 37998
rect 21532 38052 21588 38062
rect 21420 37940 21476 37950
rect 21420 37846 21476 37884
rect 21532 37716 21588 37996
rect 20748 37102 20750 37154
rect 20802 37102 20804 37154
rect 20748 37090 20804 37102
rect 20860 37660 21588 37716
rect 20748 36932 20804 36942
rect 20748 36482 20804 36876
rect 20748 36430 20750 36482
rect 20802 36430 20804 36482
rect 20748 36418 20804 36430
rect 20636 36306 20692 36316
rect 20860 35588 20916 37660
rect 21644 37378 21700 38332
rect 21644 37326 21646 37378
rect 21698 37326 21700 37378
rect 21644 37314 21700 37326
rect 21868 37940 21924 37950
rect 22316 37940 22372 39228
rect 22652 39060 22708 39454
rect 21868 37938 22372 37940
rect 21868 37886 21870 37938
rect 21922 37886 22372 37938
rect 21868 37884 22372 37886
rect 22428 39004 22708 39060
rect 22428 38050 22484 39004
rect 22540 38722 22596 38734
rect 22540 38670 22542 38722
rect 22594 38670 22596 38722
rect 22540 38388 22596 38670
rect 22652 38724 22708 38762
rect 22652 38658 22708 38668
rect 22540 38322 22596 38332
rect 22428 37998 22430 38050
rect 22482 37998 22484 38050
rect 21644 36484 21700 36494
rect 21644 36390 21700 36428
rect 21532 36260 21588 36270
rect 21532 36166 21588 36204
rect 21084 35810 21140 35822
rect 21084 35758 21086 35810
rect 21138 35758 21140 35810
rect 20412 34860 20580 34916
rect 20076 34692 20132 34730
rect 20076 34626 20132 34636
rect 20412 34690 20468 34702
rect 20412 34638 20414 34690
rect 20466 34638 20468 34690
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19852 34244 19908 34254
rect 20412 34244 20468 34638
rect 19852 34242 20468 34244
rect 19852 34190 19854 34242
rect 19906 34190 20468 34242
rect 19852 34188 20468 34190
rect 19852 33684 19908 34188
rect 19852 33618 19908 33628
rect 20524 33572 20580 34860
rect 20748 34804 20804 34814
rect 20748 34710 20804 34748
rect 20860 34020 20916 35532
rect 20412 33516 20580 33572
rect 20636 33964 20916 34020
rect 20972 35700 21028 35710
rect 20188 33122 20244 33134
rect 20188 33070 20190 33122
rect 20242 33070 20244 33122
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19516 31890 19572 31902
rect 19516 31838 19518 31890
rect 19570 31838 19572 31890
rect 19516 30434 19572 31838
rect 20188 31778 20244 33070
rect 20412 32004 20468 33516
rect 20412 31938 20468 31948
rect 20524 33346 20580 33358
rect 20524 33294 20526 33346
rect 20578 33294 20580 33346
rect 20188 31726 20190 31778
rect 20242 31726 20244 31778
rect 20188 31714 20244 31726
rect 20300 31780 20356 31790
rect 20524 31780 20580 33294
rect 20356 31724 20580 31780
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20188 31220 20244 31230
rect 20300 31220 20356 31724
rect 20188 31218 20356 31220
rect 20188 31166 20190 31218
rect 20242 31166 20356 31218
rect 20188 31164 20356 31166
rect 20188 31154 20244 31164
rect 19516 30382 19518 30434
rect 19570 30382 19572 30434
rect 19516 30324 19572 30382
rect 19516 30258 19572 30268
rect 20300 30548 20356 30558
rect 19852 30212 19908 30222
rect 19852 30118 19908 30156
rect 20300 30210 20356 30492
rect 20300 30158 20302 30210
rect 20354 30158 20356 30210
rect 20300 30146 20356 30158
rect 20524 29986 20580 29998
rect 20524 29934 20526 29986
rect 20578 29934 20580 29986
rect 20524 29876 20580 29934
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20524 29810 20580 29820
rect 19836 29754 20100 29764
rect 19852 29428 19908 29438
rect 19628 29426 19908 29428
rect 19628 29374 19854 29426
rect 19906 29374 19908 29426
rect 19628 29372 19908 29374
rect 19516 28868 19572 28878
rect 19516 28642 19572 28812
rect 19516 28590 19518 28642
rect 19570 28590 19572 28642
rect 19516 28578 19572 28590
rect 19628 28644 19684 29372
rect 19852 29362 19908 29372
rect 20524 29426 20580 29438
rect 20524 29374 20526 29426
rect 20578 29374 20580 29426
rect 19740 29092 19796 29102
rect 19740 28754 19796 29036
rect 20300 28868 20356 28878
rect 20300 28774 20356 28812
rect 20524 28868 20580 29374
rect 20524 28802 20580 28812
rect 19740 28702 19742 28754
rect 19794 28702 19796 28754
rect 19740 28690 19796 28702
rect 19964 28756 20020 28766
rect 19628 27858 19684 28588
rect 19964 28642 20020 28700
rect 19964 28590 19966 28642
rect 20018 28590 20020 28642
rect 19964 28578 20020 28590
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 27806 19630 27858
rect 19682 27806 19684 27858
rect 19628 27794 19684 27806
rect 20636 27746 20692 33964
rect 20748 33346 20804 33358
rect 20748 33294 20750 33346
rect 20802 33294 20804 33346
rect 20748 33124 20804 33294
rect 20748 33058 20804 33068
rect 20860 32452 20916 32462
rect 20860 31218 20916 32396
rect 20972 32116 21028 35644
rect 21084 33684 21140 35758
rect 21868 35588 21924 37884
rect 22428 36932 22484 37998
rect 22764 37828 22820 41692
rect 23100 41636 23156 42476
rect 23212 41972 23268 41982
rect 23324 41972 23380 44268
rect 23716 44268 23940 44324
rect 23660 44230 23716 44268
rect 23660 43652 23716 43662
rect 23660 43650 23828 43652
rect 23660 43598 23662 43650
rect 23714 43598 23828 43650
rect 23660 43596 23828 43598
rect 23660 43586 23716 43596
rect 23548 43538 23604 43550
rect 23548 43486 23550 43538
rect 23602 43486 23604 43538
rect 23436 42644 23492 42654
rect 23436 42550 23492 42588
rect 23548 42084 23604 43486
rect 23660 43314 23716 43326
rect 23660 43262 23662 43314
rect 23714 43262 23716 43314
rect 23660 42756 23716 43262
rect 23772 43092 23828 43596
rect 23772 43026 23828 43036
rect 23884 42866 23940 44268
rect 24108 44258 24164 44268
rect 23884 42814 23886 42866
rect 23938 42814 23940 42866
rect 23884 42802 23940 42814
rect 23996 44210 24052 44222
rect 23996 44158 23998 44210
rect 24050 44158 24052 44210
rect 23996 42980 24052 44158
rect 24108 43538 24164 43550
rect 24108 43486 24110 43538
rect 24162 43486 24164 43538
rect 24108 43316 24164 43486
rect 24108 43250 24164 43260
rect 23996 42756 24052 42924
rect 24108 42756 24164 42766
rect 23660 42700 23828 42756
rect 23996 42754 24164 42756
rect 23996 42702 24110 42754
rect 24162 42702 24164 42754
rect 23996 42700 24164 42702
rect 23548 42028 23716 42084
rect 23212 41970 23380 41972
rect 23212 41918 23214 41970
rect 23266 41918 23380 41970
rect 23212 41916 23380 41918
rect 23436 41972 23492 41982
rect 23492 41916 23604 41972
rect 23212 41906 23268 41916
rect 23436 41878 23492 41916
rect 23100 41580 23268 41636
rect 22988 41412 23044 41422
rect 23100 41412 23156 41422
rect 22988 41410 23100 41412
rect 22988 41358 22990 41410
rect 23042 41358 23100 41410
rect 22988 41356 23100 41358
rect 22988 41346 23044 41356
rect 22988 41076 23044 41086
rect 22988 40982 23044 41020
rect 23100 39618 23156 41356
rect 23212 40068 23268 41580
rect 23212 40002 23268 40012
rect 23100 39566 23102 39618
rect 23154 39566 23156 39618
rect 23100 39554 23156 39566
rect 23548 39618 23604 41916
rect 23660 40628 23716 42028
rect 23772 41524 23828 42700
rect 24108 42196 24164 42700
rect 24108 42130 24164 42140
rect 24220 41748 24276 45164
rect 24668 45108 24724 45118
rect 24668 45014 24724 45052
rect 24444 44882 24500 44894
rect 24444 44830 24446 44882
rect 24498 44830 24500 44882
rect 24444 44324 24500 44830
rect 24780 44660 24836 44670
rect 24556 44436 24612 44446
rect 24556 44342 24612 44380
rect 24444 44258 24500 44268
rect 24556 43428 24612 43438
rect 24556 42308 24612 43372
rect 24556 42242 24612 42252
rect 24668 41970 24724 41982
rect 24668 41918 24670 41970
rect 24722 41918 24724 41970
rect 24332 41860 24388 41870
rect 24332 41858 24612 41860
rect 24332 41806 24334 41858
rect 24386 41806 24612 41858
rect 24332 41804 24612 41806
rect 24332 41794 24388 41804
rect 23884 41524 23940 41534
rect 23772 41468 23884 41524
rect 23884 41458 23940 41468
rect 24220 41298 24276 41692
rect 24220 41246 24222 41298
rect 24274 41246 24276 41298
rect 24220 41234 24276 41246
rect 24444 41636 24500 41646
rect 24332 41188 24388 41198
rect 24332 41094 24388 41132
rect 23660 40562 23716 40572
rect 23996 40964 24052 40974
rect 23884 40290 23940 40302
rect 23884 40238 23886 40290
rect 23938 40238 23940 40290
rect 23884 40180 23940 40238
rect 23884 40114 23940 40124
rect 23548 39566 23550 39618
rect 23602 39566 23604 39618
rect 23548 39554 23604 39566
rect 23996 39620 24052 40908
rect 24108 40852 24164 40862
rect 24108 40514 24164 40796
rect 24108 40462 24110 40514
rect 24162 40462 24164 40514
rect 24108 40450 24164 40462
rect 24220 40740 24276 40750
rect 24108 39620 24164 39630
rect 23996 39618 24164 39620
rect 23996 39566 24110 39618
rect 24162 39566 24164 39618
rect 23996 39564 24164 39566
rect 22876 39394 22932 39406
rect 22876 39342 22878 39394
rect 22930 39342 22932 39394
rect 22876 37940 22932 39342
rect 23548 38948 23604 38958
rect 23548 38854 23604 38892
rect 23996 38946 24052 38958
rect 23996 38894 23998 38946
rect 24050 38894 24052 38946
rect 23996 38836 24052 38894
rect 23324 38612 23380 38622
rect 22988 38164 23044 38174
rect 22988 38162 23156 38164
rect 22988 38110 22990 38162
rect 23042 38110 23156 38162
rect 22988 38108 23156 38110
rect 22988 38098 23044 38108
rect 22876 37938 23044 37940
rect 22876 37886 22878 37938
rect 22930 37886 23044 37938
rect 22876 37884 23044 37886
rect 22876 37874 22932 37884
rect 22764 37762 22820 37772
rect 22428 36866 22484 36876
rect 22652 37156 22708 37166
rect 22316 36484 22372 36494
rect 21980 36372 22036 36382
rect 21980 36258 22036 36316
rect 21980 36206 21982 36258
rect 22034 36206 22036 36258
rect 21980 36194 22036 36206
rect 22316 35924 22372 36428
rect 22540 36370 22596 36382
rect 22540 36318 22542 36370
rect 22594 36318 22596 36370
rect 22428 35924 22484 35934
rect 22316 35922 22484 35924
rect 22316 35870 22430 35922
rect 22482 35870 22484 35922
rect 22316 35868 22484 35870
rect 22428 35700 22484 35868
rect 22428 35634 22484 35644
rect 21308 34972 21588 35028
rect 21308 33908 21364 34972
rect 21532 34914 21588 34972
rect 21532 34862 21534 34914
rect 21586 34862 21588 34914
rect 21532 34850 21588 34862
rect 21420 34802 21476 34814
rect 21420 34750 21422 34802
rect 21474 34750 21476 34802
rect 21420 34692 21476 34750
rect 21476 34636 21588 34692
rect 21420 34626 21476 34636
rect 21420 33908 21476 33918
rect 21308 33906 21476 33908
rect 21308 33854 21422 33906
rect 21474 33854 21476 33906
rect 21308 33852 21476 33854
rect 21084 33618 21140 33628
rect 21420 32676 21476 33852
rect 21420 32610 21476 32620
rect 21532 32562 21588 34636
rect 21644 33460 21700 33470
rect 21868 33460 21924 35532
rect 22540 35252 22596 36318
rect 22428 35196 22596 35252
rect 22204 34914 22260 34926
rect 22204 34862 22206 34914
rect 22258 34862 22260 34914
rect 22092 33908 22148 33918
rect 21644 33458 21924 33460
rect 21644 33406 21646 33458
rect 21698 33406 21924 33458
rect 21644 33404 21924 33406
rect 21980 33852 22092 33908
rect 21980 33458 22036 33852
rect 22092 33842 22148 33852
rect 21980 33406 21982 33458
rect 22034 33406 22036 33458
rect 21644 33394 21700 33404
rect 21980 33394 22036 33406
rect 21532 32510 21534 32562
rect 21586 32510 21588 32562
rect 21532 32498 21588 32510
rect 21868 33236 21924 33246
rect 21196 32340 21252 32350
rect 21196 32246 21252 32284
rect 20972 32060 21252 32116
rect 20860 31166 20862 31218
rect 20914 31166 20916 31218
rect 20860 31154 20916 31166
rect 20748 30994 20804 31006
rect 21084 30996 21140 31006
rect 20748 30942 20750 30994
rect 20802 30942 20804 30994
rect 20748 30772 20804 30942
rect 20748 30706 20804 30716
rect 20860 30940 21084 30996
rect 20860 30324 20916 30940
rect 21084 30902 21140 30940
rect 20748 30268 20916 30324
rect 20748 30098 20804 30268
rect 20748 30046 20750 30098
rect 20802 30046 20804 30098
rect 20748 30034 20804 30046
rect 20860 29988 20916 29998
rect 20860 29894 20916 29932
rect 20748 29428 20804 29438
rect 20748 29334 20804 29372
rect 20860 28644 20916 28654
rect 20860 28550 20916 28588
rect 21084 27972 21140 27982
rect 20636 27694 20638 27746
rect 20690 27694 20692 27746
rect 20524 27300 20580 27310
rect 19404 25890 19460 25900
rect 19516 27188 19572 27198
rect 19516 25396 19572 27132
rect 20524 27074 20580 27244
rect 20524 27022 20526 27074
rect 20578 27022 20580 27074
rect 20524 27010 20580 27022
rect 19628 26962 19684 26974
rect 19628 26910 19630 26962
rect 19682 26910 19684 26962
rect 19628 26514 19684 26910
rect 20636 26908 20692 27694
rect 20972 27858 21028 27870
rect 20972 27806 20974 27858
rect 21026 27806 21028 27858
rect 20524 26852 20692 26908
rect 20748 26962 20804 26974
rect 20748 26910 20750 26962
rect 20802 26910 20804 26962
rect 20748 26908 20804 26910
rect 20972 26908 21028 27806
rect 20748 26852 21028 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26462 19630 26514
rect 19682 26462 19684 26514
rect 19628 25732 19684 26462
rect 19628 25666 19684 25676
rect 20076 26066 20132 26078
rect 20076 26014 20078 26066
rect 20130 26014 20132 26066
rect 19516 25302 19572 25340
rect 19628 25508 19684 25518
rect 20076 25508 20132 26014
rect 20300 25732 20356 25742
rect 20300 25638 20356 25676
rect 19628 25506 20132 25508
rect 19628 25454 19630 25506
rect 19682 25454 20132 25506
rect 19628 25452 20132 25454
rect 19180 25228 19348 25284
rect 18844 24882 18900 24892
rect 18844 24722 18900 24734
rect 18844 24670 18846 24722
rect 18898 24670 18900 24722
rect 18732 24498 18788 24510
rect 18732 24446 18734 24498
rect 18786 24446 18788 24498
rect 18732 23940 18788 24446
rect 18732 23874 18788 23884
rect 18844 23828 18900 24670
rect 19180 24722 19236 24734
rect 19180 24670 19182 24722
rect 19234 24670 19236 24722
rect 19068 24610 19124 24622
rect 19068 24558 19070 24610
rect 19122 24558 19124 24610
rect 18844 23762 18900 23772
rect 18956 24164 19012 24174
rect 18956 23826 19012 24108
rect 18956 23774 18958 23826
rect 19010 23774 19012 23826
rect 18956 23604 19012 23774
rect 18956 23538 19012 23548
rect 18956 23154 19012 23166
rect 18956 23102 18958 23154
rect 19010 23102 19012 23154
rect 18956 22708 19012 23102
rect 19068 23156 19124 24558
rect 19180 24164 19236 24670
rect 19292 24388 19348 25228
rect 19628 25060 19684 25452
rect 19516 25004 19684 25060
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19292 24322 19348 24332
rect 19404 24948 19460 24958
rect 19180 24098 19236 24108
rect 19404 24052 19460 24892
rect 19180 23938 19236 23950
rect 19180 23886 19182 23938
rect 19234 23886 19236 23938
rect 19180 23828 19236 23886
rect 19180 23762 19236 23772
rect 19180 23492 19236 23502
rect 19236 23436 19348 23492
rect 19180 23426 19236 23436
rect 19068 23090 19124 23100
rect 18620 21746 18676 21756
rect 18732 22148 18788 22158
rect 18060 19814 18116 19852
rect 18396 21698 18452 21710
rect 18396 21646 18398 21698
rect 18450 21646 18452 21698
rect 18396 19684 18452 21646
rect 18620 19908 18676 19918
rect 18396 19628 18564 19684
rect 18284 19124 18340 19134
rect 18060 18450 18116 18462
rect 18060 18398 18062 18450
rect 18114 18398 18116 18450
rect 17612 18338 17780 18340
rect 17612 18286 17614 18338
rect 17666 18286 17780 18338
rect 17612 18284 17780 18286
rect 17612 18274 17668 18284
rect 17388 17826 17444 17836
rect 17612 17108 17668 17118
rect 17612 17014 17668 17052
rect 17388 16996 17444 17006
rect 17388 15986 17444 16940
rect 17388 15934 17390 15986
rect 17442 15934 17444 15986
rect 17388 15922 17444 15934
rect 17388 15428 17444 15438
rect 17388 15334 17444 15372
rect 17276 14242 17332 14252
rect 17388 13748 17444 13758
rect 17164 13746 17444 13748
rect 17164 13694 17390 13746
rect 17442 13694 17444 13746
rect 17164 13692 17444 13694
rect 17388 13682 17444 13692
rect 17612 13748 17668 13758
rect 17612 13654 17668 13692
rect 17052 12962 17108 12974
rect 17052 12910 17054 12962
rect 17106 12910 17108 12962
rect 17052 12852 17108 12910
rect 17052 12786 17108 12796
rect 17388 12850 17444 12862
rect 17388 12798 17390 12850
rect 17442 12798 17444 12850
rect 16940 12686 16942 12738
rect 16994 12686 16996 12738
rect 16940 12674 16996 12686
rect 17388 12628 17444 12798
rect 17724 12852 17780 18284
rect 18060 17892 18116 18398
rect 18060 17826 18116 17836
rect 18172 17668 18228 17678
rect 18172 17574 18228 17612
rect 17948 16996 18004 17006
rect 17948 16902 18004 16940
rect 18172 16882 18228 16894
rect 18172 16830 18174 16882
rect 18226 16830 18228 16882
rect 18172 16100 18228 16830
rect 18284 16770 18340 19068
rect 18508 18228 18564 19628
rect 18508 18134 18564 18172
rect 18620 17780 18676 19852
rect 18732 19796 18788 22092
rect 18844 21586 18900 21598
rect 18844 21534 18846 21586
rect 18898 21534 18900 21586
rect 18844 20916 18900 21534
rect 18844 20850 18900 20860
rect 18732 19730 18788 19740
rect 18956 18676 19012 22652
rect 19068 22930 19124 22942
rect 19068 22878 19070 22930
rect 19122 22878 19124 22930
rect 19068 21028 19124 22878
rect 19068 20962 19124 20972
rect 19180 21586 19236 21598
rect 19180 21534 19182 21586
rect 19234 21534 19236 21586
rect 18844 18620 19012 18676
rect 18732 17892 18788 17902
rect 18732 17798 18788 17836
rect 18620 17108 18676 17724
rect 18732 17108 18788 17118
rect 18620 17106 18788 17108
rect 18620 17054 18734 17106
rect 18786 17054 18788 17106
rect 18620 17052 18788 17054
rect 18732 17042 18788 17052
rect 18284 16718 18286 16770
rect 18338 16718 18340 16770
rect 18284 16706 18340 16718
rect 18396 16882 18452 16894
rect 18844 16884 18900 18620
rect 18956 18452 19012 18462
rect 19180 18452 19236 21534
rect 19292 21476 19348 23436
rect 19404 23378 19460 23996
rect 19404 23326 19406 23378
rect 19458 23326 19460 23378
rect 19404 23314 19460 23326
rect 19516 23156 19572 25004
rect 19628 24834 19684 24846
rect 19628 24782 19630 24834
rect 19682 24782 19684 24834
rect 19628 24388 19684 24782
rect 19964 24724 20020 24734
rect 19964 24630 20020 24668
rect 20412 24500 20468 24510
rect 19628 24322 19684 24332
rect 20300 24498 20468 24500
rect 20300 24446 20414 24498
rect 20466 24446 20468 24498
rect 20300 24444 20468 24446
rect 19628 24164 19684 24174
rect 19628 23938 19684 24108
rect 20188 24052 20244 24062
rect 19628 23886 19630 23938
rect 19682 23886 19684 23938
rect 19628 23874 19684 23886
rect 19964 23938 20020 23950
rect 19964 23886 19966 23938
rect 20018 23886 20020 23938
rect 19964 23828 20020 23886
rect 20076 23940 20132 23950
rect 20076 23846 20132 23884
rect 20188 23938 20244 23996
rect 20188 23886 20190 23938
rect 20242 23886 20244 23938
rect 20188 23874 20244 23886
rect 19964 23762 20020 23772
rect 19740 23716 19796 23726
rect 19628 23714 19796 23716
rect 19628 23662 19742 23714
rect 19794 23662 19796 23714
rect 19628 23660 19796 23662
rect 19628 23380 19684 23660
rect 19740 23650 19796 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23314 19684 23324
rect 19628 23156 19684 23166
rect 19516 23154 19684 23156
rect 19516 23102 19630 23154
rect 19682 23102 19684 23154
rect 19516 23100 19684 23102
rect 19628 23090 19684 23100
rect 19516 22372 19572 22382
rect 19516 21810 19572 22316
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19516 21758 19518 21810
rect 19570 21758 19572 21810
rect 19516 21746 19572 21758
rect 19628 21812 19684 21822
rect 19628 21718 19684 21756
rect 20076 21812 20132 21822
rect 20132 21756 20244 21812
rect 20076 21746 20132 21756
rect 19404 21700 19460 21710
rect 19404 21606 19460 21644
rect 19964 21700 20020 21710
rect 19964 21606 20020 21644
rect 19292 21410 19348 21420
rect 20076 21476 20132 21486
rect 19628 20916 19684 20926
rect 19516 19460 19572 19470
rect 19516 19346 19572 19404
rect 19516 19294 19518 19346
rect 19570 19294 19572 19346
rect 19516 19282 19572 19294
rect 19628 19234 19684 20860
rect 20076 20802 20132 21420
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20738 20132 20750
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20244 20244 21756
rect 20300 21810 20356 24444
rect 20412 24434 20468 24444
rect 20524 23716 20580 26852
rect 20748 25620 20804 26852
rect 20748 25554 20804 25564
rect 20860 25508 20916 25518
rect 20636 25284 20692 25294
rect 20636 25282 20804 25284
rect 20636 25230 20638 25282
rect 20690 25230 20804 25282
rect 20636 25228 20804 25230
rect 20636 25218 20692 25228
rect 20524 23650 20580 23660
rect 20748 24498 20804 25228
rect 20748 24446 20750 24498
rect 20802 24446 20804 24498
rect 20524 23268 20580 23278
rect 20748 23268 20804 24446
rect 20524 23266 20804 23268
rect 20524 23214 20526 23266
rect 20578 23214 20804 23266
rect 20524 23212 20804 23214
rect 20524 23202 20580 23212
rect 20300 21758 20302 21810
rect 20354 21758 20356 21810
rect 20300 21746 20356 21758
rect 20524 22482 20580 22494
rect 20524 22430 20526 22482
rect 20578 22430 20580 22482
rect 20524 21812 20580 22430
rect 20860 21812 20916 25452
rect 20972 24724 21028 24734
rect 20972 24388 21028 24668
rect 21084 24612 21140 27916
rect 21196 27076 21252 32060
rect 21868 32004 21924 33180
rect 21868 31938 21924 31948
rect 22092 33122 22148 33134
rect 22092 33070 22094 33122
rect 22146 33070 22148 33122
rect 22092 31948 22148 33070
rect 22204 32674 22260 34862
rect 22428 34132 22484 35196
rect 22540 35028 22596 35038
rect 22540 34934 22596 34972
rect 22652 34354 22708 37100
rect 22876 36260 22932 36270
rect 22876 36166 22932 36204
rect 22988 35810 23044 37884
rect 22988 35758 22990 35810
rect 23042 35758 23044 35810
rect 22988 35746 23044 35758
rect 23100 35140 23156 38108
rect 23324 38050 23380 38556
rect 23324 37998 23326 38050
rect 23378 37998 23380 38050
rect 23324 36596 23380 37998
rect 23548 37268 23604 37278
rect 23324 36594 23492 36596
rect 23324 36542 23326 36594
rect 23378 36542 23492 36594
rect 23324 36540 23492 36542
rect 23324 36530 23380 36540
rect 23212 35700 23268 35710
rect 23268 35644 23380 35700
rect 23212 35606 23268 35644
rect 23100 35084 23268 35140
rect 23100 34914 23156 34926
rect 23100 34862 23102 34914
rect 23154 34862 23156 34914
rect 23100 34356 23156 34862
rect 22652 34302 22654 34354
rect 22706 34302 22708 34354
rect 22652 34290 22708 34302
rect 22876 34300 23156 34356
rect 22876 34132 22932 34300
rect 23212 34244 23268 35084
rect 23324 35138 23380 35644
rect 23436 35252 23492 36540
rect 23548 35700 23604 37212
rect 23660 37042 23716 37054
rect 23660 36990 23662 37042
rect 23714 36990 23716 37042
rect 23660 36932 23716 36990
rect 23660 35700 23716 36876
rect 23996 36596 24052 38780
rect 24108 38050 24164 39564
rect 24220 38834 24276 40684
rect 24444 40626 24500 41580
rect 24444 40574 24446 40626
rect 24498 40574 24500 40626
rect 24444 40562 24500 40574
rect 24332 40514 24388 40526
rect 24332 40462 24334 40514
rect 24386 40462 24388 40514
rect 24332 40404 24388 40462
rect 24332 40348 24500 40404
rect 24220 38782 24222 38834
rect 24274 38782 24276 38834
rect 24220 38500 24276 38782
rect 24444 38668 24500 40348
rect 24556 39730 24612 41804
rect 24668 40852 24724 41918
rect 24668 40786 24724 40796
rect 24780 40740 24836 44604
rect 24892 44324 24948 45276
rect 24892 44230 24948 44268
rect 24892 42754 24948 42766
rect 24892 42702 24894 42754
rect 24946 42702 24948 42754
rect 24892 41972 24948 42702
rect 24892 41906 24948 41916
rect 24780 40674 24836 40684
rect 24668 40628 24724 40638
rect 24668 40534 24724 40572
rect 24556 39678 24558 39730
rect 24610 39678 24612 39730
rect 24556 39058 24612 39678
rect 24556 39006 24558 39058
rect 24610 39006 24612 39058
rect 24556 38994 24612 39006
rect 25004 38668 25060 46284
rect 25116 45778 25172 45790
rect 25116 45726 25118 45778
rect 25170 45726 25172 45778
rect 25116 45332 25172 45726
rect 25116 45266 25172 45276
rect 25228 44996 25284 47012
rect 25452 46956 25620 47012
rect 25676 49810 25844 49812
rect 25676 49758 25790 49810
rect 25842 49758 25844 49810
rect 25676 49756 25844 49758
rect 25452 46564 25508 46956
rect 25564 46788 25620 46798
rect 25564 46694 25620 46732
rect 25452 46508 25620 46564
rect 25340 45778 25396 45790
rect 25340 45726 25342 45778
rect 25394 45726 25396 45778
rect 25340 45556 25396 45726
rect 25340 45332 25396 45500
rect 25452 45332 25508 45342
rect 25340 45276 25452 45332
rect 25452 45266 25508 45276
rect 25116 44940 25284 44996
rect 25116 44660 25172 44940
rect 25452 44660 25508 44670
rect 25116 44604 25284 44660
rect 25116 44436 25172 44446
rect 25116 42532 25172 44380
rect 25228 42980 25284 44604
rect 25340 44324 25396 44334
rect 25340 43538 25396 44268
rect 25452 43650 25508 44604
rect 25452 43598 25454 43650
rect 25506 43598 25508 43650
rect 25452 43586 25508 43598
rect 25340 43486 25342 43538
rect 25394 43486 25396 43538
rect 25340 43474 25396 43486
rect 25452 43428 25508 43438
rect 25228 42924 25396 42980
rect 25228 42756 25284 42766
rect 25228 42662 25284 42700
rect 25228 42532 25284 42542
rect 25116 42530 25284 42532
rect 25116 42478 25230 42530
rect 25282 42478 25284 42530
rect 25116 42476 25284 42478
rect 25228 42466 25284 42476
rect 25340 42084 25396 42924
rect 25228 42028 25396 42084
rect 25228 40628 25284 42028
rect 25340 41860 25396 41870
rect 25452 41860 25508 43372
rect 25340 41858 25508 41860
rect 25340 41806 25342 41858
rect 25394 41806 25508 41858
rect 25340 41804 25508 41806
rect 25340 41636 25396 41804
rect 25340 41570 25396 41580
rect 25340 40628 25396 40638
rect 25284 40626 25396 40628
rect 25284 40574 25342 40626
rect 25394 40574 25396 40626
rect 25284 40572 25396 40574
rect 25228 40534 25284 40572
rect 25340 40562 25396 40572
rect 25564 40180 25620 46508
rect 25676 45332 25732 49756
rect 25788 49746 25844 49756
rect 26572 50372 26852 50428
rect 25900 48020 25956 48030
rect 25900 47926 25956 47964
rect 26572 47684 26628 50372
rect 27020 49252 27076 52556
rect 27804 52500 27860 54572
rect 27916 53730 27972 55468
rect 27916 53678 27918 53730
rect 27970 53678 27972 53730
rect 27916 53666 27972 53678
rect 28028 54514 28084 54526
rect 28028 54462 28030 54514
rect 28082 54462 28084 54514
rect 28028 52724 28084 54462
rect 28140 54404 28196 55468
rect 28252 55412 28308 58158
rect 28588 58210 28644 58222
rect 28588 58158 28590 58210
rect 28642 58158 28644 58210
rect 28476 57876 28532 57886
rect 28476 57540 28532 57820
rect 28476 57446 28532 57484
rect 28252 55346 28308 55356
rect 28476 57204 28532 57214
rect 28476 55298 28532 57148
rect 28588 56308 28644 58158
rect 28588 56242 28644 56252
rect 28812 58212 28868 58222
rect 28812 56420 28868 58156
rect 28812 56194 28868 56364
rect 28812 56142 28814 56194
rect 28866 56142 28868 56194
rect 28812 56130 28868 56142
rect 28476 55246 28478 55298
rect 28530 55246 28532 55298
rect 28476 55234 28532 55246
rect 28252 55076 28308 55086
rect 28252 54982 28308 55020
rect 28476 54628 28532 54638
rect 28476 54534 28532 54572
rect 28700 54514 28756 54526
rect 28700 54462 28702 54514
rect 28754 54462 28756 54514
rect 28140 54348 28532 54404
rect 28140 53620 28196 53630
rect 28140 53172 28196 53564
rect 28476 53618 28532 54348
rect 28476 53566 28478 53618
rect 28530 53566 28532 53618
rect 28476 53554 28532 53566
rect 28588 53732 28644 53742
rect 28588 53618 28644 53676
rect 28588 53566 28590 53618
rect 28642 53566 28644 53618
rect 28252 53508 28308 53518
rect 28252 53414 28308 53452
rect 28140 53170 28308 53172
rect 28140 53118 28142 53170
rect 28194 53118 28308 53170
rect 28140 53116 28308 53118
rect 28140 53106 28196 53116
rect 28028 52658 28084 52668
rect 27244 52444 27860 52500
rect 27132 52164 27188 52174
rect 27132 50034 27188 52108
rect 27132 49982 27134 50034
rect 27186 49982 27188 50034
rect 27132 49970 27188 49982
rect 27020 49186 27076 49196
rect 27132 49812 27188 49822
rect 26684 48916 26740 48926
rect 26684 48822 26740 48860
rect 26572 47590 26628 47628
rect 25788 47458 25844 47470
rect 25788 47406 25790 47458
rect 25842 47406 25844 47458
rect 25788 45890 25844 47406
rect 26012 47460 26068 47470
rect 26012 47348 26068 47404
rect 26908 47348 26964 47358
rect 26012 47346 26180 47348
rect 26012 47294 26014 47346
rect 26066 47294 26180 47346
rect 26012 47292 26180 47294
rect 26012 47282 26068 47292
rect 25788 45838 25790 45890
rect 25842 45838 25844 45890
rect 25788 45780 25844 45838
rect 25788 45714 25844 45724
rect 25900 47236 25956 47246
rect 25900 45444 25956 47180
rect 26012 45892 26068 45902
rect 26012 45798 26068 45836
rect 26012 45668 26068 45678
rect 26012 45574 26068 45612
rect 25900 45388 26068 45444
rect 25676 45266 25732 45276
rect 25900 45220 25956 45230
rect 25676 44994 25732 45006
rect 25676 44942 25678 44994
rect 25730 44942 25732 44994
rect 25676 44772 25732 44942
rect 25676 44706 25732 44716
rect 25900 44772 25956 45164
rect 26012 45106 26068 45388
rect 26124 45332 26180 47292
rect 26908 47254 26964 47292
rect 26236 46676 26292 46686
rect 26236 45556 26292 46620
rect 26348 45890 26404 45902
rect 26348 45838 26350 45890
rect 26402 45838 26404 45890
rect 26348 45780 26404 45838
rect 26796 45892 26852 45902
rect 26796 45798 26852 45836
rect 27020 45890 27076 45902
rect 27020 45838 27022 45890
rect 27074 45838 27076 45890
rect 26572 45780 26628 45790
rect 26348 45778 26628 45780
rect 26348 45726 26574 45778
rect 26626 45726 26628 45778
rect 26348 45724 26628 45726
rect 26236 45490 26292 45500
rect 26348 45332 26404 45342
rect 26124 45330 26404 45332
rect 26124 45278 26350 45330
rect 26402 45278 26404 45330
rect 26124 45276 26404 45278
rect 26348 45266 26404 45276
rect 26572 45220 26628 45724
rect 26908 45780 26964 45790
rect 26684 45666 26740 45678
rect 26684 45614 26686 45666
rect 26738 45614 26740 45666
rect 26684 45556 26740 45614
rect 26684 45490 26740 45500
rect 26796 45668 26852 45678
rect 26572 45154 26628 45164
rect 26012 45054 26014 45106
rect 26066 45054 26068 45106
rect 26012 44996 26068 45054
rect 26012 44930 26068 44940
rect 25900 44706 25956 44716
rect 26236 44660 26292 44670
rect 25676 44322 25732 44334
rect 25676 44270 25678 44322
rect 25730 44270 25732 44322
rect 25676 42754 25732 44270
rect 25900 44212 25956 44222
rect 25900 44210 26068 44212
rect 25900 44158 25902 44210
rect 25954 44158 26068 44210
rect 25900 44156 26068 44158
rect 25900 44146 25956 44156
rect 25676 42702 25678 42754
rect 25730 42702 25732 42754
rect 25676 41412 25732 42702
rect 26012 42644 26068 44156
rect 26236 44210 26292 44604
rect 26796 44434 26852 45612
rect 26796 44382 26798 44434
rect 26850 44382 26852 44434
rect 26796 44370 26852 44382
rect 26236 44158 26238 44210
rect 26290 44158 26292 44210
rect 26124 43540 26180 43550
rect 26124 43446 26180 43484
rect 26236 43428 26292 44158
rect 26460 44212 26516 44222
rect 26460 43650 26516 44156
rect 26460 43598 26462 43650
rect 26514 43598 26516 43650
rect 26460 43586 26516 43598
rect 26908 43650 26964 45724
rect 27020 45108 27076 45838
rect 27132 45444 27188 49756
rect 27244 48916 27300 52444
rect 27580 52276 27636 52286
rect 28252 52276 28308 53116
rect 28588 53060 28644 53566
rect 28700 53172 28756 54462
rect 28700 53106 28756 53116
rect 28588 52994 28644 53004
rect 27580 50428 27636 52220
rect 27804 52274 28308 52276
rect 27804 52222 28254 52274
rect 28306 52222 28308 52274
rect 27804 52220 28308 52222
rect 27804 52164 27860 52220
rect 28252 52210 28308 52220
rect 27804 51602 27860 52108
rect 28924 52052 28980 52062
rect 28924 51604 28980 51996
rect 27804 51550 27806 51602
rect 27858 51550 27860 51602
rect 27804 51538 27860 51550
rect 28588 51602 28980 51604
rect 28588 51550 28926 51602
rect 28978 51550 28980 51602
rect 28588 51548 28980 51550
rect 28028 50596 28084 50606
rect 28028 50502 28084 50540
rect 28588 50594 28644 51548
rect 28924 51538 28980 51548
rect 28588 50542 28590 50594
rect 28642 50542 28644 50594
rect 28588 50530 28644 50542
rect 29036 50428 29092 59612
rect 29148 59602 29204 59612
rect 29596 59106 29652 59118
rect 29596 59054 29598 59106
rect 29650 59054 29652 59106
rect 29148 58772 29204 58782
rect 29148 57204 29204 58716
rect 29596 58772 29652 59054
rect 29596 58706 29652 58716
rect 29484 58660 29540 58670
rect 29484 58566 29540 58604
rect 29596 58436 29652 58446
rect 29596 58342 29652 58380
rect 29260 57652 29316 57662
rect 29260 57558 29316 57596
rect 29596 57652 29652 57662
rect 29708 57652 29764 59836
rect 31164 59892 31220 59902
rect 31164 59798 31220 59836
rect 32732 59892 32788 59902
rect 29820 59778 29876 59790
rect 29820 59726 29822 59778
rect 29874 59726 29876 59778
rect 29820 59332 29876 59726
rect 30044 59780 30100 59790
rect 30044 59442 30100 59724
rect 30044 59390 30046 59442
rect 30098 59390 30100 59442
rect 30044 59378 30100 59390
rect 32172 59778 32228 59790
rect 32172 59726 32174 59778
rect 32226 59726 32228 59778
rect 29820 59108 29876 59276
rect 29820 59042 29876 59052
rect 30828 59330 30884 59342
rect 30828 59278 30830 59330
rect 30882 59278 30884 59330
rect 30268 58884 30324 58894
rect 30156 58436 30212 58446
rect 30156 58322 30212 58380
rect 30156 58270 30158 58322
rect 30210 58270 30212 58322
rect 30156 58258 30212 58270
rect 29596 57650 29764 57652
rect 29596 57598 29598 57650
rect 29650 57598 29764 57650
rect 29596 57596 29764 57598
rect 30156 57652 30212 57662
rect 29596 57586 29652 57596
rect 30156 57558 30212 57596
rect 29148 56756 29204 57148
rect 29484 57540 29540 57550
rect 29260 56756 29316 56766
rect 29148 56754 29428 56756
rect 29148 56702 29262 56754
rect 29314 56702 29428 56754
rect 29148 56700 29428 56702
rect 29260 56690 29316 56700
rect 29148 56308 29204 56318
rect 29148 56194 29204 56252
rect 29148 56142 29150 56194
rect 29202 56142 29204 56194
rect 29148 56130 29204 56142
rect 29372 56082 29428 56700
rect 29372 56030 29374 56082
rect 29426 56030 29428 56082
rect 29372 56018 29428 56030
rect 29484 55468 29540 57484
rect 29820 57538 29876 57550
rect 29820 57486 29822 57538
rect 29874 57486 29876 57538
rect 29820 57204 29876 57486
rect 29820 57138 29876 57148
rect 29596 56866 29652 56878
rect 29596 56814 29598 56866
rect 29650 56814 29652 56866
rect 29596 56196 29652 56814
rect 29932 56756 29988 56766
rect 29932 56754 30100 56756
rect 29932 56702 29934 56754
rect 29986 56702 30100 56754
rect 29932 56700 30100 56702
rect 29932 56690 29988 56700
rect 29596 56082 29652 56140
rect 29596 56030 29598 56082
rect 29650 56030 29652 56082
rect 29596 56018 29652 56030
rect 29708 56532 29764 56542
rect 29148 55412 29540 55468
rect 29596 55412 29652 55422
rect 29708 55412 29764 56476
rect 29932 56084 29988 56094
rect 29932 55990 29988 56028
rect 29148 54516 29204 55412
rect 29596 55410 29764 55412
rect 29596 55358 29598 55410
rect 29650 55358 29764 55410
rect 29596 55356 29764 55358
rect 29596 55346 29652 55356
rect 29260 55298 29316 55310
rect 29260 55246 29262 55298
rect 29314 55246 29316 55298
rect 29260 54852 29316 55246
rect 29484 55298 29540 55310
rect 29484 55246 29486 55298
rect 29538 55246 29540 55298
rect 29484 54964 29540 55246
rect 29820 55300 29876 55310
rect 29820 55298 29988 55300
rect 29820 55246 29822 55298
rect 29874 55246 29988 55298
rect 29820 55244 29988 55246
rect 29820 55234 29876 55244
rect 29484 54908 29876 54964
rect 29260 54796 29540 54852
rect 29484 54740 29540 54796
rect 29484 54646 29540 54684
rect 29148 54450 29204 54460
rect 29260 54514 29316 54526
rect 29260 54462 29262 54514
rect 29314 54462 29316 54514
rect 29260 53730 29316 54462
rect 29260 53678 29262 53730
rect 29314 53678 29316 53730
rect 29260 53172 29316 53678
rect 29484 54514 29540 54526
rect 29484 54462 29486 54514
rect 29538 54462 29540 54514
rect 29484 53396 29540 54462
rect 29708 54514 29764 54526
rect 29708 54462 29710 54514
rect 29762 54462 29764 54514
rect 29708 53732 29764 54462
rect 29820 53844 29876 54908
rect 29932 54516 29988 55244
rect 29932 54450 29988 54460
rect 30044 55298 30100 56700
rect 30268 56308 30324 58828
rect 30380 58772 30436 58782
rect 30380 56866 30436 58716
rect 30828 56980 30884 59278
rect 31164 58996 31220 59006
rect 31164 58434 31220 58940
rect 32172 58996 32228 59726
rect 32284 59778 32340 59790
rect 32284 59726 32286 59778
rect 32338 59726 32340 59778
rect 32284 59220 32340 59726
rect 32284 59154 32340 59164
rect 32396 59780 32452 59790
rect 32620 59780 32676 59790
rect 32172 58930 32228 58940
rect 31164 58382 31166 58434
rect 31218 58382 31220 58434
rect 31164 57650 31220 58382
rect 31164 57598 31166 57650
rect 31218 57598 31220 57650
rect 31164 57586 31220 57598
rect 31276 58772 31332 58782
rect 31276 58434 31332 58716
rect 31276 58382 31278 58434
rect 31330 58382 31332 58434
rect 31164 56980 31220 56990
rect 30828 56978 31220 56980
rect 30828 56926 31166 56978
rect 31218 56926 31220 56978
rect 30828 56924 31220 56926
rect 31164 56914 31220 56924
rect 30380 56814 30382 56866
rect 30434 56814 30436 56866
rect 30380 56802 30436 56814
rect 30604 56866 30660 56878
rect 30604 56814 30606 56866
rect 30658 56814 30660 56866
rect 30492 56644 30548 56654
rect 30380 56308 30436 56318
rect 30268 56306 30436 56308
rect 30268 56254 30382 56306
rect 30434 56254 30436 56306
rect 30268 56252 30436 56254
rect 30380 56242 30436 56252
rect 30492 56194 30548 56588
rect 30492 56142 30494 56194
rect 30546 56142 30548 56194
rect 30492 56130 30548 56142
rect 30604 56196 30660 56814
rect 31276 56754 31332 58382
rect 32172 58436 32228 58446
rect 31724 57538 31780 57550
rect 31724 57486 31726 57538
rect 31778 57486 31780 57538
rect 31276 56702 31278 56754
rect 31330 56702 31332 56754
rect 31052 56642 31108 56654
rect 31052 56590 31054 56642
rect 31106 56590 31108 56642
rect 31052 56532 31108 56590
rect 31276 56644 31332 56702
rect 31388 56756 31444 56766
rect 31388 56662 31444 56700
rect 31500 56754 31556 56766
rect 31500 56702 31502 56754
rect 31554 56702 31556 56754
rect 31276 56578 31332 56588
rect 31052 56466 31108 56476
rect 30380 55858 30436 55870
rect 30380 55806 30382 55858
rect 30434 55806 30436 55858
rect 30156 55412 30212 55422
rect 30156 55318 30212 55356
rect 30044 55246 30046 55298
rect 30098 55246 30100 55298
rect 30044 53956 30100 55246
rect 30380 55300 30436 55806
rect 30380 55244 30548 55300
rect 30268 55188 30324 55198
rect 30268 55186 30436 55188
rect 30268 55134 30270 55186
rect 30322 55134 30436 55186
rect 30268 55132 30436 55134
rect 30268 55122 30324 55132
rect 30156 54740 30212 54750
rect 30156 54514 30212 54684
rect 30156 54462 30158 54514
rect 30210 54462 30212 54514
rect 30156 54450 30212 54462
rect 30380 54292 30436 55132
rect 30156 53956 30212 53966
rect 30044 53954 30212 53956
rect 30044 53902 30158 53954
rect 30210 53902 30212 53954
rect 30044 53900 30212 53902
rect 30156 53890 30212 53900
rect 30380 53954 30436 54236
rect 30380 53902 30382 53954
rect 30434 53902 30436 53954
rect 30380 53890 30436 53902
rect 29820 53788 30100 53844
rect 29708 53676 29988 53732
rect 29708 53508 29764 53518
rect 29708 53414 29764 53452
rect 29484 53340 29652 53396
rect 29260 53078 29316 53116
rect 29372 52836 29428 52846
rect 29260 52164 29316 52174
rect 29148 52052 29204 52062
rect 29148 51958 29204 51996
rect 29260 51938 29316 52108
rect 29260 51886 29262 51938
rect 29314 51886 29316 51938
rect 29260 51874 29316 51886
rect 29372 51602 29428 52780
rect 29372 51550 29374 51602
rect 29426 51550 29428 51602
rect 29372 51538 29428 51550
rect 29596 51602 29652 53340
rect 29708 53172 29764 53210
rect 29708 53106 29764 53116
rect 29596 51550 29598 51602
rect 29650 51550 29652 51602
rect 29372 50482 29428 50494
rect 29372 50430 29374 50482
rect 29426 50430 29428 50482
rect 29372 50428 29428 50430
rect 27580 50372 27860 50428
rect 29036 50372 29316 50428
rect 29372 50372 29540 50428
rect 27804 49812 27860 50372
rect 27804 49746 27860 49756
rect 27692 49700 27748 49710
rect 27692 49140 27748 49644
rect 29036 49588 29092 49598
rect 29036 49494 29092 49532
rect 27692 49138 27972 49140
rect 27692 49086 27694 49138
rect 27746 49086 27972 49138
rect 27692 49084 27972 49086
rect 27692 49074 27748 49084
rect 27244 48466 27300 48860
rect 27244 48414 27246 48466
rect 27298 48414 27300 48466
rect 27244 48402 27300 48414
rect 27804 47570 27860 47582
rect 27804 47518 27806 47570
rect 27858 47518 27860 47570
rect 27580 47236 27636 47246
rect 27132 45378 27188 45388
rect 27244 47234 27636 47236
rect 27244 47182 27582 47234
rect 27634 47182 27636 47234
rect 27244 47180 27636 47182
rect 27020 43762 27076 45052
rect 27020 43710 27022 43762
rect 27074 43710 27076 43762
rect 27020 43698 27076 43710
rect 26908 43598 26910 43650
rect 26962 43598 26964 43650
rect 26908 43586 26964 43598
rect 26236 43362 26292 43372
rect 26796 43316 26852 43326
rect 26236 42644 26292 42654
rect 26012 42642 26292 42644
rect 26012 42590 26238 42642
rect 26290 42590 26292 42642
rect 26012 42588 26292 42590
rect 26124 42196 26180 42206
rect 26124 42102 26180 42140
rect 26236 42084 26292 42588
rect 26348 42084 26404 42094
rect 26236 42082 26516 42084
rect 26236 42030 26350 42082
rect 26402 42030 26516 42082
rect 26236 42028 26516 42030
rect 26348 42018 26404 42028
rect 25676 41346 25732 41356
rect 25788 41970 25844 41982
rect 25788 41918 25790 41970
rect 25842 41918 25844 41970
rect 25676 40516 25732 40526
rect 25676 40422 25732 40460
rect 25788 40292 25844 41918
rect 26012 41972 26068 41982
rect 26012 41878 26068 41916
rect 26348 41524 26404 41534
rect 26012 40740 26068 40750
rect 25340 40124 25620 40180
rect 25676 40236 25844 40292
rect 25900 40626 25956 40638
rect 25900 40574 25902 40626
rect 25954 40574 25956 40626
rect 24444 38612 24612 38668
rect 24220 38434 24276 38444
rect 24108 37998 24110 38050
rect 24162 37998 24164 38050
rect 24108 37986 24164 37998
rect 24556 37938 24612 38612
rect 24556 37886 24558 37938
rect 24610 37886 24612 37938
rect 24556 36708 24612 37886
rect 24780 38612 25060 38668
rect 25228 39508 25284 39518
rect 24668 37156 24724 37166
rect 24668 37062 24724 37100
rect 24668 36708 24724 36718
rect 24556 36706 24724 36708
rect 24556 36654 24670 36706
rect 24722 36654 24724 36706
rect 24556 36652 24724 36654
rect 24668 36642 24724 36652
rect 23996 36482 24052 36540
rect 23996 36430 23998 36482
rect 24050 36430 24052 36482
rect 23996 36418 24052 36430
rect 24332 36372 24388 36382
rect 24332 36278 24388 36316
rect 24108 35700 24164 35710
rect 23660 35698 24164 35700
rect 23660 35646 24110 35698
rect 24162 35646 24164 35698
rect 23660 35644 24164 35646
rect 23548 35634 23604 35644
rect 24108 35634 24164 35644
rect 24444 35588 24500 35598
rect 24444 35494 24500 35532
rect 23548 35476 23604 35486
rect 23548 35382 23604 35420
rect 23436 35196 23604 35252
rect 23324 35086 23326 35138
rect 23378 35086 23380 35138
rect 23324 35074 23380 35086
rect 23548 34692 23604 35196
rect 23660 34916 23716 34926
rect 23996 34916 24052 34926
rect 23660 34914 24052 34916
rect 23660 34862 23662 34914
rect 23714 34862 23998 34914
rect 24050 34862 24052 34914
rect 23660 34860 24052 34862
rect 23660 34850 23716 34860
rect 23996 34850 24052 34860
rect 23548 34636 23940 34692
rect 23100 34188 23268 34244
rect 23324 34244 23380 34254
rect 22428 34076 22932 34132
rect 22988 34130 23044 34142
rect 22988 34078 22990 34130
rect 23042 34078 23044 34130
rect 22428 33124 22484 34076
rect 22876 33908 22932 33918
rect 22876 33814 22932 33852
rect 22988 33460 23044 34078
rect 22540 33404 23044 33460
rect 22540 33346 22596 33404
rect 22540 33294 22542 33346
rect 22594 33294 22596 33346
rect 22540 33282 22596 33294
rect 22428 33068 22708 33124
rect 22204 32622 22206 32674
rect 22258 32622 22260 32674
rect 22204 32340 22260 32622
rect 22316 32676 22372 32686
rect 22316 32562 22372 32620
rect 22316 32510 22318 32562
rect 22370 32510 22372 32562
rect 22316 32498 22372 32510
rect 22204 32284 22596 32340
rect 22316 32004 22372 32014
rect 22092 31892 22260 31948
rect 22316 31910 22372 31948
rect 22540 32004 22596 32284
rect 22540 31938 22596 31948
rect 21532 31780 21588 31818
rect 21532 31714 21588 31724
rect 22092 31780 22148 31790
rect 22204 31780 22260 31892
rect 22540 31780 22596 31790
rect 22204 31778 22596 31780
rect 22204 31726 22542 31778
rect 22594 31726 22596 31778
rect 22204 31724 22596 31726
rect 21308 31668 21364 31678
rect 21308 31574 21364 31612
rect 21980 31668 22036 31678
rect 21308 30994 21364 31006
rect 21308 30942 21310 30994
rect 21362 30942 21364 30994
rect 21308 30884 21364 30942
rect 21308 30818 21364 30828
rect 21420 30324 21476 30334
rect 21420 30210 21476 30268
rect 21420 30158 21422 30210
rect 21474 30158 21476 30210
rect 21420 28082 21476 30158
rect 21868 30100 21924 30110
rect 21420 28030 21422 28082
rect 21474 28030 21476 28082
rect 21420 28018 21476 28030
rect 21644 29428 21700 29438
rect 21644 28082 21700 29372
rect 21756 29204 21812 29214
rect 21868 29204 21924 30044
rect 21756 29202 21924 29204
rect 21756 29150 21758 29202
rect 21810 29150 21924 29202
rect 21756 29148 21924 29150
rect 21756 29138 21812 29148
rect 21644 28030 21646 28082
rect 21698 28030 21700 28082
rect 21644 28018 21700 28030
rect 21756 28642 21812 28654
rect 21756 28590 21758 28642
rect 21810 28590 21812 28642
rect 21756 27972 21812 28590
rect 21756 27906 21812 27916
rect 21868 27858 21924 29148
rect 21868 27806 21870 27858
rect 21922 27806 21924 27858
rect 21868 27794 21924 27806
rect 21196 27010 21252 27020
rect 21756 27746 21812 27758
rect 21756 27694 21758 27746
rect 21810 27694 21812 27746
rect 21644 26962 21700 26974
rect 21644 26910 21646 26962
rect 21698 26910 21700 26962
rect 21308 26402 21364 26414
rect 21308 26350 21310 26402
rect 21362 26350 21364 26402
rect 21308 25060 21364 26350
rect 21644 25844 21700 26910
rect 21644 25778 21700 25788
rect 21532 25396 21588 25406
rect 21532 25302 21588 25340
rect 21308 25004 21588 25060
rect 21308 24834 21364 24846
rect 21308 24782 21310 24834
rect 21362 24782 21364 24834
rect 21308 24724 21364 24782
rect 21308 24658 21364 24668
rect 21420 24722 21476 24734
rect 21420 24670 21422 24722
rect 21474 24670 21476 24722
rect 21084 24546 21140 24556
rect 20972 22932 21028 24332
rect 21420 23828 21476 24670
rect 21084 23156 21140 23166
rect 21084 23154 21252 23156
rect 21084 23102 21086 23154
rect 21138 23102 21252 23154
rect 21084 23100 21252 23102
rect 21084 23090 21140 23100
rect 20972 22876 21140 22932
rect 20524 21756 20916 21812
rect 20412 21700 20468 21710
rect 20412 20802 20468 21644
rect 20636 21588 20692 21598
rect 20636 21494 20692 21532
rect 20412 20750 20414 20802
rect 20466 20750 20468 20802
rect 20412 20738 20468 20750
rect 20636 20804 20692 20814
rect 20636 20710 20692 20748
rect 20524 20578 20580 20590
rect 20524 20526 20526 20578
rect 20578 20526 20580 20578
rect 20524 20244 20580 20526
rect 20524 20188 20692 20244
rect 20076 19906 20132 19918
rect 20076 19854 20078 19906
rect 20130 19854 20132 19906
rect 20076 19460 20132 19854
rect 20076 19394 20132 19404
rect 19628 19182 19630 19234
rect 19682 19182 19684 19234
rect 19628 19170 19684 19182
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19852 18452 19908 18462
rect 19180 18450 19908 18452
rect 19180 18398 19854 18450
rect 19906 18398 19908 18450
rect 19180 18396 19908 18398
rect 18956 18358 19012 18396
rect 19068 18340 19124 18350
rect 18396 16830 18398 16882
rect 18450 16830 18452 16882
rect 18396 16772 18452 16830
rect 18396 16706 18452 16716
rect 18508 16828 18900 16884
rect 18956 17668 19012 17678
rect 18956 17106 19012 17612
rect 18956 17054 18958 17106
rect 19010 17054 19012 17106
rect 17836 15202 17892 15214
rect 17836 15150 17838 15202
rect 17890 15150 17892 15202
rect 17836 14532 17892 15150
rect 17836 14466 17892 14476
rect 17948 14530 18004 14542
rect 17948 14478 17950 14530
rect 18002 14478 18004 14530
rect 17836 14306 17892 14318
rect 17836 14254 17838 14306
rect 17890 14254 17892 14306
rect 17836 13076 17892 14254
rect 17948 13970 18004 14478
rect 17948 13918 17950 13970
rect 18002 13918 18004 13970
rect 17948 13906 18004 13918
rect 17836 13010 17892 13020
rect 17948 13076 18004 13086
rect 18172 13076 18228 16044
rect 18396 14308 18452 14318
rect 17948 13074 18228 13076
rect 17948 13022 17950 13074
rect 18002 13022 18228 13074
rect 17948 13020 18228 13022
rect 18284 14196 18340 14206
rect 17948 13010 18004 13020
rect 18172 12852 18228 12862
rect 18284 12852 18340 14140
rect 17724 12796 18116 12852
rect 17388 12572 17780 12628
rect 16828 12460 17668 12516
rect 16828 12290 16884 12460
rect 17612 12402 17668 12460
rect 17612 12350 17614 12402
rect 17666 12350 17668 12402
rect 17612 12338 17668 12350
rect 16828 12238 16830 12290
rect 16882 12238 16884 12290
rect 16828 12226 16884 12238
rect 16492 12126 16494 12178
rect 16546 12126 16548 12178
rect 16044 11900 16324 11956
rect 15932 11890 15988 11900
rect 16268 11506 16324 11900
rect 16268 11454 16270 11506
rect 16322 11454 16324 11506
rect 16268 11442 16324 11454
rect 16492 11396 16548 12126
rect 17388 12178 17444 12190
rect 17388 12126 17390 12178
rect 17442 12126 17444 12178
rect 16492 11282 16548 11340
rect 16716 11732 16772 11742
rect 16716 11394 16772 11676
rect 16828 11620 16884 11630
rect 16828 11526 16884 11564
rect 16716 11342 16718 11394
rect 16770 11342 16772 11394
rect 16716 11330 16772 11342
rect 17052 11396 17108 11406
rect 17388 11396 17444 12126
rect 17724 12180 17780 12572
rect 17052 11394 17444 11396
rect 17052 11342 17054 11394
rect 17106 11342 17444 11394
rect 17052 11340 17444 11342
rect 17500 12068 17556 12078
rect 17052 11330 17108 11340
rect 16492 11230 16494 11282
rect 16546 11230 16548 11282
rect 16492 11218 16548 11230
rect 16604 11172 16660 11182
rect 16156 10724 16212 10734
rect 16044 10500 16100 10510
rect 16044 10406 16100 10444
rect 16044 9940 16100 9950
rect 16156 9940 16212 10668
rect 16044 9938 16212 9940
rect 16044 9886 16046 9938
rect 16098 9886 16212 9938
rect 16044 9884 16212 9886
rect 16380 10722 16436 10734
rect 16380 10670 16382 10722
rect 16434 10670 16436 10722
rect 16044 9874 16100 9884
rect 16380 9828 16436 10670
rect 16380 9762 16436 9772
rect 16492 10610 16548 10622
rect 16492 10558 16494 10610
rect 16546 10558 16548 10610
rect 16492 10052 16548 10558
rect 15708 9602 15764 9614
rect 15708 9550 15710 9602
rect 15762 9550 15764 9602
rect 15708 9492 15764 9550
rect 15708 8596 15764 9436
rect 15932 9602 15988 9614
rect 15932 9550 15934 9602
rect 15986 9550 15988 9602
rect 15932 9044 15988 9550
rect 16156 9602 16212 9614
rect 16156 9550 16158 9602
rect 16210 9550 16212 9602
rect 16156 9156 16212 9550
rect 16380 9156 16436 9166
rect 16156 9154 16436 9156
rect 16156 9102 16382 9154
rect 16434 9102 16436 9154
rect 16156 9100 16436 9102
rect 15932 9042 16100 9044
rect 15932 8990 15934 9042
rect 15986 8990 16100 9042
rect 15932 8988 16100 8990
rect 15932 8978 15988 8988
rect 15708 8530 15764 8540
rect 15596 8372 15764 8428
rect 15596 7362 15652 7374
rect 15596 7310 15598 7362
rect 15650 7310 15652 7362
rect 15596 7028 15652 7310
rect 15596 6962 15652 6972
rect 15372 6130 15540 6132
rect 15372 6078 15374 6130
rect 15426 6078 15540 6130
rect 15372 6076 15540 6078
rect 15708 6132 15764 8372
rect 16044 8260 16100 8988
rect 15932 8036 15988 8046
rect 15932 7942 15988 7980
rect 16044 7698 16100 8204
rect 16044 7646 16046 7698
rect 16098 7646 16100 7698
rect 16044 7634 16100 7646
rect 16156 8932 16212 8942
rect 15932 7476 15988 7486
rect 15932 7382 15988 7420
rect 15820 6692 15876 6702
rect 15820 6598 15876 6636
rect 15820 6132 15876 6142
rect 15708 6130 15876 6132
rect 15708 6078 15822 6130
rect 15874 6078 15876 6130
rect 15708 6076 15876 6078
rect 15372 6066 15428 6076
rect 15820 6066 15876 6076
rect 16044 6132 16100 6142
rect 16044 5234 16100 6076
rect 16156 5796 16212 8876
rect 16380 8372 16436 9100
rect 16492 8932 16548 9996
rect 16492 8866 16548 8876
rect 16268 8260 16324 8270
rect 16380 8260 16436 8316
rect 16268 8258 16436 8260
rect 16268 8206 16270 8258
rect 16322 8206 16436 8258
rect 16268 8204 16436 8206
rect 16492 8708 16548 8718
rect 16268 8194 16324 8204
rect 16268 6692 16324 6702
rect 16268 6598 16324 6636
rect 16492 6132 16548 8652
rect 16604 7586 16660 11116
rect 17052 10276 17108 10286
rect 16940 10052 16996 10062
rect 16828 9996 16940 10052
rect 16716 8372 16772 8382
rect 16716 7698 16772 8316
rect 16716 7646 16718 7698
rect 16770 7646 16772 7698
rect 16716 7634 16772 7646
rect 16604 7534 16606 7586
rect 16658 7534 16660 7586
rect 16604 6690 16660 7534
rect 16716 7252 16772 7262
rect 16828 7252 16884 9996
rect 16940 9986 16996 9996
rect 16940 9828 16996 9838
rect 16940 9602 16996 9772
rect 17052 9826 17108 10220
rect 17052 9774 17054 9826
rect 17106 9774 17108 9826
rect 17052 9762 17108 9774
rect 16940 9550 16942 9602
rect 16994 9550 16996 9602
rect 16940 9538 16996 9550
rect 17164 9604 17220 11340
rect 17500 10500 17556 12012
rect 17612 11620 17668 11630
rect 17612 11394 17668 11564
rect 17612 11342 17614 11394
rect 17666 11342 17668 11394
rect 17612 11330 17668 11342
rect 17724 11508 17780 12124
rect 17836 12178 17892 12190
rect 17836 12126 17838 12178
rect 17890 12126 17892 12178
rect 17836 11732 17892 12126
rect 17948 12178 18004 12190
rect 17948 12126 17950 12178
rect 18002 12126 18004 12178
rect 17948 12068 18004 12126
rect 17948 12002 18004 12012
rect 17836 11666 17892 11676
rect 17836 11508 17892 11518
rect 17724 11506 17892 11508
rect 17724 11454 17838 11506
rect 17890 11454 17892 11506
rect 17724 11452 17892 11454
rect 18060 11508 18116 12796
rect 18172 12850 18340 12852
rect 18172 12798 18174 12850
rect 18226 12798 18340 12850
rect 18172 12796 18340 12798
rect 18172 12786 18228 12796
rect 18396 12404 18452 14252
rect 18508 13076 18564 16828
rect 18956 16098 19012 17054
rect 19068 17666 19124 18284
rect 19852 18116 19908 18396
rect 20188 18450 20244 20188
rect 20636 20132 20692 20188
rect 20636 20066 20692 20076
rect 20188 18398 20190 18450
rect 20242 18398 20244 18450
rect 20188 18386 20244 18398
rect 20300 20018 20356 20030
rect 20524 20020 20580 20030
rect 20300 19966 20302 20018
rect 20354 19966 20356 20018
rect 20300 18452 20356 19966
rect 20412 19964 20524 20020
rect 20412 19234 20468 19964
rect 20524 19926 20580 19964
rect 20412 19182 20414 19234
rect 20466 19182 20468 19234
rect 20412 19170 20468 19182
rect 20300 18386 20356 18396
rect 20524 18452 20580 18462
rect 19852 18060 20356 18116
rect 19628 17778 19684 17790
rect 19628 17726 19630 17778
rect 19682 17726 19684 17778
rect 19068 17614 19070 17666
rect 19122 17614 19124 17666
rect 19068 16994 19124 17614
rect 19068 16942 19070 16994
rect 19122 16942 19124 16994
rect 19068 16930 19124 16942
rect 19292 17666 19348 17678
rect 19292 17614 19294 17666
rect 19346 17614 19348 17666
rect 18956 16046 18958 16098
rect 19010 16046 19012 16098
rect 18956 16034 19012 16046
rect 19068 16770 19124 16782
rect 19068 16718 19070 16770
rect 19122 16718 19124 16770
rect 18732 15202 18788 15214
rect 18732 15150 18734 15202
rect 18786 15150 18788 15202
rect 18732 15092 18788 15150
rect 18620 14756 18676 14766
rect 18620 14642 18676 14700
rect 18620 14590 18622 14642
rect 18674 14590 18676 14642
rect 18620 14578 18676 14590
rect 18732 14196 18788 15036
rect 18732 14130 18788 14140
rect 18956 14420 19012 14430
rect 18956 13970 19012 14364
rect 18956 13918 18958 13970
rect 19010 13918 19012 13970
rect 18956 13906 19012 13918
rect 18620 13860 18676 13870
rect 18620 13766 18676 13804
rect 19068 13748 19124 16718
rect 19292 15092 19348 17614
rect 19516 16882 19572 16894
rect 19516 16830 19518 16882
rect 19570 16830 19572 16882
rect 19516 16212 19572 16830
rect 19516 16146 19572 16156
rect 19292 15026 19348 15036
rect 19516 14980 19572 14990
rect 19516 14418 19572 14924
rect 19516 14366 19518 14418
rect 19570 14366 19572 14418
rect 19516 14354 19572 14366
rect 19068 13682 19124 13692
rect 19628 13412 19684 17726
rect 20076 17780 20132 17790
rect 20076 17686 20132 17724
rect 20188 17668 20244 17678
rect 20188 17574 20244 17612
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20300 16658 20356 18060
rect 20524 17892 20580 18396
rect 20412 16996 20468 17006
rect 20412 16902 20468 16940
rect 20524 16882 20580 17836
rect 20636 17780 20692 17790
rect 20636 17220 20692 17724
rect 20748 17332 20804 21756
rect 20972 21700 21028 21710
rect 20972 21606 21028 21644
rect 21084 21588 21140 22876
rect 21084 21522 21140 21532
rect 21196 20916 21252 23100
rect 21420 22482 21476 23772
rect 21420 22430 21422 22482
rect 21474 22430 21476 22482
rect 21420 22418 21476 22430
rect 21532 23716 21588 25004
rect 21420 22036 21476 22046
rect 21308 21812 21364 21822
rect 21308 21698 21364 21756
rect 21308 21646 21310 21698
rect 21362 21646 21364 21698
rect 21308 21634 21364 21646
rect 21308 20916 21364 20926
rect 21196 20914 21364 20916
rect 21196 20862 21310 20914
rect 21362 20862 21364 20914
rect 21196 20860 21364 20862
rect 21308 20850 21364 20860
rect 21420 20802 21476 21980
rect 21420 20750 21422 20802
rect 21474 20750 21476 20802
rect 21420 20738 21476 20750
rect 21420 20020 21476 20030
rect 21420 19926 21476 19964
rect 21420 19460 21476 19470
rect 21420 19366 21476 19404
rect 21308 17556 21364 17566
rect 21532 17556 21588 23660
rect 21644 23042 21700 23054
rect 21644 22990 21646 23042
rect 21698 22990 21700 23042
rect 21644 22484 21700 22990
rect 21644 22418 21700 22428
rect 21756 22372 21812 27694
rect 21980 26962 22036 31612
rect 22092 30994 22148 31724
rect 22540 31106 22596 31724
rect 22540 31054 22542 31106
rect 22594 31054 22596 31106
rect 22540 31042 22596 31054
rect 22092 30942 22094 30994
rect 22146 30942 22148 30994
rect 22092 30930 22148 30942
rect 22428 30884 22484 30894
rect 22428 30790 22484 30828
rect 22652 30660 22708 33068
rect 22764 32786 22820 33404
rect 22764 32734 22766 32786
rect 22818 32734 22820 32786
rect 22764 32452 22820 32734
rect 22876 32676 22932 32686
rect 22876 32582 22932 32620
rect 22764 32396 22932 32452
rect 22764 31780 22820 31790
rect 22764 31686 22820 31724
rect 22876 31778 22932 32396
rect 23100 31892 23156 34188
rect 23212 34018 23268 34030
rect 23212 33966 23214 34018
rect 23266 33966 23268 34018
rect 23212 33234 23268 33966
rect 23212 33182 23214 33234
rect 23266 33182 23268 33234
rect 23212 33170 23268 33182
rect 23324 32788 23380 34188
rect 23436 34132 23492 34142
rect 23436 34038 23492 34076
rect 23660 33908 23716 33918
rect 23660 33814 23716 33852
rect 23436 33684 23492 33694
rect 23436 33012 23492 33628
rect 23436 32956 23604 33012
rect 23436 32788 23492 32798
rect 23324 32786 23492 32788
rect 23324 32734 23438 32786
rect 23490 32734 23492 32786
rect 23324 32732 23492 32734
rect 23436 32722 23492 32732
rect 22876 31726 22878 31778
rect 22930 31726 22932 31778
rect 22876 31714 22932 31726
rect 22988 31836 23156 31892
rect 23212 31892 23268 31902
rect 22428 30604 22708 30660
rect 22204 29988 22260 29998
rect 22204 29426 22260 29932
rect 22204 29374 22206 29426
rect 22258 29374 22260 29426
rect 22204 29362 22260 29374
rect 22316 29204 22372 29214
rect 22428 29204 22484 30604
rect 22988 30436 23044 31836
rect 23100 31666 23156 31678
rect 23100 31614 23102 31666
rect 23154 31614 23156 31666
rect 23100 31556 23156 31614
rect 23100 31490 23156 31500
rect 23212 31220 23268 31836
rect 23548 31668 23604 32956
rect 23772 32338 23828 32350
rect 23772 32286 23774 32338
rect 23826 32286 23828 32338
rect 23772 32116 23828 32286
rect 23772 32050 23828 32060
rect 23548 31574 23604 31612
rect 23660 31668 23716 31678
rect 23660 31666 23828 31668
rect 23660 31614 23662 31666
rect 23714 31614 23828 31666
rect 23660 31612 23828 31614
rect 23660 31602 23716 31612
rect 23212 31154 23268 31164
rect 23324 31554 23380 31566
rect 23324 31502 23326 31554
rect 23378 31502 23380 31554
rect 22372 29148 22484 29204
rect 22540 30380 23044 30436
rect 23100 31106 23156 31118
rect 23100 31054 23102 31106
rect 23154 31054 23156 31106
rect 23100 30996 23156 31054
rect 22316 29138 22372 29148
rect 22204 29092 22260 29102
rect 22204 27858 22260 29036
rect 22540 28980 22596 30380
rect 23100 30324 23156 30940
rect 23212 30994 23268 31006
rect 23212 30942 23214 30994
rect 23266 30942 23268 30994
rect 23212 30772 23268 30942
rect 23212 30706 23268 30716
rect 23212 30324 23268 30334
rect 23100 30268 23212 30324
rect 22652 30210 22708 30222
rect 22652 30158 22654 30210
rect 22706 30158 22708 30210
rect 22652 29428 22708 30158
rect 22652 29362 22708 29372
rect 23100 29426 23156 30268
rect 23212 30258 23268 30268
rect 23100 29374 23102 29426
rect 23154 29374 23156 29426
rect 23100 29362 23156 29374
rect 22204 27806 22206 27858
rect 22258 27806 22260 27858
rect 22204 27794 22260 27806
rect 22316 28924 22596 28980
rect 22764 29202 22820 29214
rect 22764 29150 22766 29202
rect 22818 29150 22820 29202
rect 21980 26910 21982 26962
rect 22034 26910 22036 26962
rect 21980 26898 22036 26910
rect 22316 26908 22372 28924
rect 22428 28532 22484 28542
rect 22428 28530 22708 28532
rect 22428 28478 22430 28530
rect 22482 28478 22708 28530
rect 22428 28476 22708 28478
rect 22428 28466 22484 28476
rect 22652 28082 22708 28476
rect 22652 28030 22654 28082
rect 22706 28030 22708 28082
rect 22652 28018 22708 28030
rect 22764 28084 22820 29150
rect 22764 28028 22932 28084
rect 22540 27858 22596 27870
rect 22540 27806 22542 27858
rect 22594 27806 22596 27858
rect 22428 27076 22484 27114
rect 22428 27010 22484 27020
rect 22540 26908 22596 27806
rect 22764 27860 22820 27870
rect 22764 27766 22820 27804
rect 22316 26852 22484 26908
rect 22540 26852 22708 26908
rect 22316 26402 22372 26414
rect 22316 26350 22318 26402
rect 22370 26350 22372 26402
rect 22204 26292 22260 26302
rect 22204 26198 22260 26236
rect 22092 25620 22148 25630
rect 21868 25508 21924 25518
rect 21868 25414 21924 25452
rect 22092 24724 22148 25564
rect 22316 25620 22372 26350
rect 22316 25554 22372 25564
rect 22428 25506 22484 26852
rect 22428 25454 22430 25506
rect 22482 25454 22484 25506
rect 22428 25442 22484 25454
rect 22540 26290 22596 26302
rect 22540 26238 22542 26290
rect 22594 26238 22596 26290
rect 22540 25508 22596 26238
rect 22540 25442 22596 25452
rect 22204 25396 22260 25406
rect 22204 25302 22260 25340
rect 22204 24724 22260 24734
rect 22092 24722 22260 24724
rect 22092 24670 22206 24722
rect 22258 24670 22260 24722
rect 22092 24668 22260 24670
rect 21868 23826 21924 23838
rect 21868 23774 21870 23826
rect 21922 23774 21924 23826
rect 21868 23716 21924 23774
rect 21868 23650 21924 23660
rect 21980 23604 22036 23614
rect 21756 22306 21812 22316
rect 21868 22372 21924 22382
rect 21980 22372 22036 23548
rect 21868 22370 22036 22372
rect 21868 22318 21870 22370
rect 21922 22318 22036 22370
rect 21868 22316 22036 22318
rect 21868 22036 21924 22316
rect 21868 21970 21924 21980
rect 21980 22148 22036 22158
rect 21644 21698 21700 21710
rect 21980 21700 22036 22092
rect 21644 21646 21646 21698
rect 21698 21646 21700 21698
rect 21644 21476 21700 21646
rect 21644 21410 21700 21420
rect 21868 21644 22036 21700
rect 21868 20802 21924 21644
rect 21980 21474 22036 21486
rect 21980 21422 21982 21474
rect 22034 21422 22036 21474
rect 21980 21364 22036 21422
rect 21980 21298 22036 21308
rect 21868 20750 21870 20802
rect 21922 20750 21924 20802
rect 21756 20244 21812 20254
rect 21756 19458 21812 20188
rect 21756 19406 21758 19458
rect 21810 19406 21812 19458
rect 21756 18340 21812 19406
rect 21756 18274 21812 18284
rect 21868 20020 21924 20750
rect 22204 20692 22260 24668
rect 22652 24612 22708 26852
rect 22764 26404 22820 26414
rect 22764 25730 22820 26348
rect 22764 25678 22766 25730
rect 22818 25678 22820 25730
rect 22764 25666 22820 25678
rect 22764 25284 22820 25294
rect 22764 24834 22820 25228
rect 22764 24782 22766 24834
rect 22818 24782 22820 24834
rect 22764 24770 22820 24782
rect 22876 24836 22932 28028
rect 23212 27860 23268 27870
rect 23324 27860 23380 31502
rect 23548 30994 23604 31006
rect 23548 30942 23550 30994
rect 23602 30942 23604 30994
rect 23436 30772 23492 30782
rect 23436 29314 23492 30716
rect 23548 30548 23604 30942
rect 23772 30996 23828 31612
rect 23884 31556 23940 34636
rect 24668 34356 24724 34366
rect 24780 34356 24836 38612
rect 25228 38274 25284 39452
rect 25228 38222 25230 38274
rect 25282 38222 25284 38274
rect 25228 38210 25284 38222
rect 25340 38052 25396 40124
rect 25676 39172 25732 40236
rect 25900 39508 25956 40574
rect 26012 40514 26068 40684
rect 26012 40462 26014 40514
rect 26066 40462 26068 40514
rect 26012 40450 26068 40462
rect 26236 40402 26292 40414
rect 26236 40350 26238 40402
rect 26290 40350 26292 40402
rect 26124 40068 26180 40078
rect 26124 39730 26180 40012
rect 26124 39678 26126 39730
rect 26178 39678 26180 39730
rect 26124 39666 26180 39678
rect 25900 39452 26068 39508
rect 25676 39116 25844 39172
rect 25564 39058 25620 39070
rect 25564 39006 25566 39058
rect 25618 39006 25620 39058
rect 25564 38948 25620 39006
rect 25564 38882 25620 38892
rect 25788 38836 25844 39116
rect 25676 38724 25732 38762
rect 25676 38658 25732 38668
rect 25564 38500 25620 38510
rect 25340 37996 25508 38052
rect 25340 37828 25396 37838
rect 25452 37828 25508 37996
rect 25564 38050 25620 38444
rect 25564 37998 25566 38050
rect 25618 37998 25620 38050
rect 25564 37986 25620 37998
rect 25676 38388 25732 38398
rect 25452 37772 25620 37828
rect 25340 37490 25396 37772
rect 25340 37438 25342 37490
rect 25394 37438 25396 37490
rect 25340 37426 25396 37438
rect 25452 36708 25508 36718
rect 25452 36484 25508 36652
rect 25116 36482 25508 36484
rect 25116 36430 25454 36482
rect 25506 36430 25508 36482
rect 25116 36428 25508 36430
rect 25116 34914 25172 36428
rect 25452 36418 25508 36428
rect 25116 34862 25118 34914
rect 25170 34862 25172 34914
rect 25116 34850 25172 34862
rect 25228 35700 25284 35710
rect 24668 34354 24836 34356
rect 24668 34302 24670 34354
rect 24722 34302 24836 34354
rect 24668 34300 24836 34302
rect 24892 34802 24948 34814
rect 24892 34750 24894 34802
rect 24946 34750 24948 34802
rect 24668 34290 24724 34300
rect 24556 34244 24612 34254
rect 24444 34188 24556 34244
rect 24108 34018 24164 34030
rect 24108 33966 24110 34018
rect 24162 33966 24164 34018
rect 24108 33124 24164 33966
rect 24332 34020 24388 34030
rect 24332 33926 24388 33964
rect 24108 33058 24164 33068
rect 24444 33796 24500 34188
rect 24556 34178 24612 34188
rect 24444 32562 24500 33740
rect 24780 33684 24836 33694
rect 24556 32676 24612 32686
rect 24780 32676 24836 33628
rect 24556 32674 24836 32676
rect 24556 32622 24558 32674
rect 24610 32622 24836 32674
rect 24556 32620 24836 32622
rect 24556 32610 24612 32620
rect 24444 32510 24446 32562
rect 24498 32510 24500 32562
rect 24444 32498 24500 32510
rect 24668 32004 24724 32014
rect 24332 31892 24388 31902
rect 23996 31780 24052 31790
rect 23996 31686 24052 31724
rect 24332 31778 24388 31836
rect 24332 31726 24334 31778
rect 24386 31726 24388 31778
rect 24332 31714 24388 31726
rect 24444 31666 24500 31678
rect 24444 31614 24446 31666
rect 24498 31614 24500 31666
rect 24332 31556 24388 31566
rect 24444 31556 24500 31614
rect 24556 31668 24612 31678
rect 24556 31574 24612 31612
rect 23884 31500 24052 31556
rect 23660 30884 23716 30894
rect 23660 30790 23716 30828
rect 23548 30482 23604 30492
rect 23436 29262 23438 29314
rect 23490 29262 23492 29314
rect 23436 29250 23492 29262
rect 23436 27972 23492 27982
rect 23436 27878 23492 27916
rect 23212 27858 23380 27860
rect 23212 27806 23214 27858
rect 23266 27806 23380 27858
rect 23212 27804 23380 27806
rect 23660 27858 23716 27870
rect 23660 27806 23662 27858
rect 23714 27806 23716 27858
rect 23212 27794 23268 27804
rect 23660 27524 23716 27806
rect 23660 27458 23716 27468
rect 23660 27300 23716 27310
rect 22876 24770 22932 24780
rect 22988 27074 23044 27086
rect 22988 27022 22990 27074
rect 23042 27022 23044 27074
rect 22988 24612 23044 27022
rect 23324 27076 23380 27086
rect 23324 26962 23380 27020
rect 23660 27074 23716 27244
rect 23660 27022 23662 27074
rect 23714 27022 23716 27074
rect 23660 27010 23716 27022
rect 23324 26910 23326 26962
rect 23378 26910 23380 26962
rect 23324 26898 23380 26910
rect 23324 26404 23380 26414
rect 23324 26310 23380 26348
rect 23772 26180 23828 30940
rect 23884 30994 23940 31006
rect 23884 30942 23886 30994
rect 23938 30942 23940 30994
rect 23884 30436 23940 30942
rect 23996 30660 24052 31500
rect 24388 31500 24500 31556
rect 24668 31554 24724 31948
rect 24668 31502 24670 31554
rect 24722 31502 24724 31554
rect 24332 31490 24388 31500
rect 24668 31444 24724 31502
rect 24444 31388 24724 31444
rect 24108 31108 24164 31118
rect 24108 31106 24276 31108
rect 24108 31054 24110 31106
rect 24162 31054 24276 31106
rect 24108 31052 24276 31054
rect 24108 31042 24164 31052
rect 23996 30604 24164 30660
rect 23996 30436 24052 30446
rect 23884 30380 23996 30436
rect 23884 30100 23940 30110
rect 23884 30006 23940 30044
rect 23884 29876 23940 29886
rect 23996 29876 24052 30380
rect 23940 29820 24052 29876
rect 23884 29810 23940 29820
rect 23996 29428 24052 29438
rect 23996 29334 24052 29372
rect 24108 29204 24164 30604
rect 24220 29428 24276 31052
rect 24332 30994 24388 31006
rect 24332 30942 24334 30994
rect 24386 30942 24388 30994
rect 24332 29652 24388 30942
rect 24332 29586 24388 29596
rect 24220 29334 24276 29372
rect 23772 26114 23828 26124
rect 23996 29148 24164 29204
rect 23996 25844 24052 29148
rect 24220 27860 24276 27870
rect 24220 27766 24276 27804
rect 24332 27858 24388 27870
rect 24332 27806 24334 27858
rect 24386 27806 24388 27858
rect 24332 27748 24388 27806
rect 24108 27074 24164 27086
rect 24108 27022 24110 27074
rect 24162 27022 24164 27074
rect 24108 26740 24164 27022
rect 24332 26962 24388 27692
rect 24444 27412 24500 31388
rect 24556 31220 24612 31230
rect 24556 31126 24612 31164
rect 24668 30996 24724 31006
rect 24668 30902 24724 30940
rect 24668 30548 24724 30558
rect 24668 30434 24724 30492
rect 24668 30382 24670 30434
rect 24722 30382 24724 30434
rect 24556 30212 24612 30222
rect 24556 30118 24612 30156
rect 24668 29316 24724 30382
rect 24668 29250 24724 29260
rect 24556 28756 24612 28766
rect 24556 28662 24612 28700
rect 24780 28532 24836 32620
rect 24556 28476 24836 28532
rect 24556 28082 24612 28476
rect 24556 28030 24558 28082
rect 24610 28030 24612 28082
rect 24556 28018 24612 28030
rect 24668 27972 24724 27982
rect 24668 27878 24724 27916
rect 24444 27346 24500 27356
rect 24332 26910 24334 26962
rect 24386 26910 24388 26962
rect 24332 26898 24388 26910
rect 24668 26962 24724 26974
rect 24668 26910 24670 26962
rect 24722 26910 24724 26962
rect 24668 26908 24724 26910
rect 24556 26852 24724 26908
rect 24556 26740 24612 26852
rect 24108 26684 24612 26740
rect 23660 25788 24052 25844
rect 24220 26292 24276 26302
rect 22316 24556 22708 24612
rect 22764 24556 23044 24612
rect 23548 25508 23604 25518
rect 23660 25508 23716 25788
rect 24220 25732 24276 26236
rect 24556 26068 24612 26684
rect 24892 26404 24948 34750
rect 25004 33684 25060 33694
rect 25004 33124 25060 33628
rect 25228 33572 25284 35644
rect 25564 34244 25620 37772
rect 25676 37378 25732 38332
rect 25788 38050 25844 38780
rect 25788 37998 25790 38050
rect 25842 37998 25844 38050
rect 25788 37986 25844 37998
rect 25900 38948 25956 38958
rect 25676 37326 25678 37378
rect 25730 37326 25732 37378
rect 25676 37314 25732 37326
rect 25900 37266 25956 38892
rect 25900 37214 25902 37266
rect 25954 37214 25956 37266
rect 25900 37202 25956 37214
rect 25676 36482 25732 36494
rect 25676 36430 25678 36482
rect 25730 36430 25732 36482
rect 25676 36260 25732 36430
rect 25676 34914 25732 36204
rect 26012 35810 26068 39452
rect 26124 39284 26180 39294
rect 26124 39058 26180 39228
rect 26124 39006 26126 39058
rect 26178 39006 26180 39058
rect 26124 38612 26180 39006
rect 26236 38724 26292 40350
rect 26348 39618 26404 41468
rect 26348 39566 26350 39618
rect 26402 39566 26404 39618
rect 26348 39554 26404 39566
rect 26460 39508 26516 42028
rect 26572 41970 26628 41982
rect 26572 41918 26574 41970
rect 26626 41918 26628 41970
rect 26572 41412 26628 41918
rect 26796 41860 26852 43260
rect 26908 42868 26964 42878
rect 27244 42868 27300 47180
rect 27580 47170 27636 47180
rect 27468 47012 27524 47022
rect 27804 47012 27860 47518
rect 27468 46898 27524 46956
rect 27468 46846 27470 46898
rect 27522 46846 27524 46898
rect 27468 46834 27524 46846
rect 27692 46956 27860 47012
rect 27468 46116 27524 46126
rect 27468 45890 27524 46060
rect 27468 45838 27470 45890
rect 27522 45838 27524 45890
rect 27468 45826 27524 45838
rect 27580 45668 27636 45678
rect 27356 45666 27636 45668
rect 27356 45614 27582 45666
rect 27634 45614 27636 45666
rect 27356 45612 27636 45614
rect 27356 43092 27412 45612
rect 27580 45602 27636 45612
rect 27692 44210 27748 46956
rect 27804 46676 27860 46686
rect 27804 46582 27860 46620
rect 27916 46228 27972 49084
rect 28252 49028 28308 49038
rect 28252 49026 28420 49028
rect 28252 48974 28254 49026
rect 28306 48974 28420 49026
rect 28252 48972 28420 48974
rect 28252 48962 28308 48972
rect 27916 46162 27972 46172
rect 28028 48914 28084 48926
rect 28028 48862 28030 48914
rect 28082 48862 28084 48914
rect 28028 48356 28084 48862
rect 28028 47124 28084 48300
rect 28252 48244 28308 48254
rect 28364 48244 28420 48972
rect 28588 48804 28644 48814
rect 28588 48802 29204 48804
rect 28588 48750 28590 48802
rect 28642 48750 29204 48802
rect 28588 48748 29204 48750
rect 28588 48738 28644 48748
rect 28588 48244 28644 48254
rect 28364 48242 28644 48244
rect 28364 48190 28590 48242
rect 28642 48190 28644 48242
rect 28364 48188 28644 48190
rect 28028 46002 28084 47068
rect 28028 45950 28030 46002
rect 28082 45950 28084 46002
rect 28028 45938 28084 45950
rect 28140 47572 28196 47582
rect 28140 47346 28196 47516
rect 28140 47294 28142 47346
rect 28194 47294 28196 47346
rect 28140 46562 28196 47294
rect 28252 47346 28308 48188
rect 28476 48020 28532 48188
rect 28588 48178 28644 48188
rect 29036 48244 29092 48254
rect 29036 48150 29092 48188
rect 28252 47294 28254 47346
rect 28306 47294 28308 47346
rect 28252 47282 28308 47294
rect 28364 47908 28420 47918
rect 28364 47346 28420 47852
rect 28364 47294 28366 47346
rect 28418 47294 28420 47346
rect 28364 47282 28420 47294
rect 28140 46510 28142 46562
rect 28194 46510 28196 46562
rect 27804 45666 27860 45678
rect 27804 45614 27806 45666
rect 27858 45614 27860 45666
rect 27804 44436 27860 45614
rect 28140 45444 28196 46510
rect 28252 46116 28308 46126
rect 28476 46116 28532 47964
rect 28924 48018 28980 48030
rect 28924 47966 28926 48018
rect 28978 47966 28980 48018
rect 28700 47460 28756 47470
rect 28588 47404 28700 47460
rect 28588 47346 28644 47404
rect 28700 47394 28756 47404
rect 28588 47294 28590 47346
rect 28642 47294 28644 47346
rect 28588 47282 28644 47294
rect 28812 46786 28868 46798
rect 28812 46734 28814 46786
rect 28866 46734 28868 46786
rect 28252 46114 28532 46116
rect 28252 46062 28254 46114
rect 28306 46062 28532 46114
rect 28252 46060 28532 46062
rect 28588 46674 28644 46686
rect 28588 46622 28590 46674
rect 28642 46622 28644 46674
rect 28588 46114 28644 46622
rect 28588 46062 28590 46114
rect 28642 46062 28644 46114
rect 28252 46050 28308 46060
rect 28588 46050 28644 46062
rect 27804 44370 27860 44380
rect 27916 45388 28196 45444
rect 27692 44158 27694 44210
rect 27746 44158 27748 44210
rect 27692 44146 27748 44158
rect 27804 44212 27860 44222
rect 27804 44118 27860 44156
rect 27916 44098 27972 45388
rect 28140 45218 28196 45230
rect 28140 45166 28142 45218
rect 28194 45166 28196 45218
rect 28028 44436 28084 44446
rect 28140 44436 28196 45166
rect 28028 44434 28196 44436
rect 28028 44382 28030 44434
rect 28082 44382 28196 44434
rect 28028 44380 28196 44382
rect 28252 45220 28308 45230
rect 28028 44370 28084 44380
rect 27916 44046 27918 44098
rect 27970 44046 27972 44098
rect 27916 43988 27972 44046
rect 27692 43932 27972 43988
rect 28140 44098 28196 44110
rect 28140 44046 28142 44098
rect 28194 44046 28196 44098
rect 27468 43650 27524 43662
rect 27468 43598 27470 43650
rect 27522 43598 27524 43650
rect 27468 43316 27524 43598
rect 27692 43538 27748 43932
rect 27692 43486 27694 43538
rect 27746 43486 27748 43538
rect 27692 43474 27748 43486
rect 27804 43540 27860 43550
rect 27580 43316 27636 43326
rect 27468 43260 27580 43316
rect 27580 43250 27636 43260
rect 27356 43036 27748 43092
rect 27244 42812 27636 42868
rect 26908 42530 26964 42812
rect 27244 42642 27300 42654
rect 27244 42590 27246 42642
rect 27298 42590 27300 42642
rect 26908 42478 26910 42530
rect 26962 42478 26964 42530
rect 26908 42082 26964 42478
rect 27020 42530 27076 42542
rect 27020 42478 27022 42530
rect 27074 42478 27076 42530
rect 27020 42196 27076 42478
rect 27132 42530 27188 42542
rect 27132 42478 27134 42530
rect 27186 42478 27188 42530
rect 27132 42308 27188 42478
rect 27132 42242 27188 42252
rect 27244 42420 27300 42590
rect 27020 42130 27076 42140
rect 26908 42030 26910 42082
rect 26962 42030 26964 42082
rect 26908 42018 26964 42030
rect 27244 42084 27300 42364
rect 27244 42018 27300 42028
rect 27356 42642 27412 42654
rect 27356 42590 27358 42642
rect 27410 42590 27412 42642
rect 27132 41970 27188 41982
rect 27132 41918 27134 41970
rect 27186 41918 27188 41970
rect 27132 41860 27188 41918
rect 26796 41804 27188 41860
rect 27356 41748 27412 42590
rect 27356 41682 27412 41692
rect 27468 42532 27524 42542
rect 27468 41524 27524 42476
rect 26572 41346 26628 41356
rect 27244 41468 27524 41524
rect 27132 40962 27188 40974
rect 27132 40910 27134 40962
rect 27186 40910 27188 40962
rect 27020 40628 27076 40638
rect 26460 39442 26516 39452
rect 26796 40402 26852 40414
rect 26796 40350 26798 40402
rect 26850 40350 26852 40402
rect 26796 39284 26852 40350
rect 26796 39218 26852 39228
rect 26908 38836 26964 38846
rect 26236 38668 26628 38724
rect 26124 38546 26180 38556
rect 26572 37378 26628 38668
rect 26572 37326 26574 37378
rect 26626 37326 26628 37378
rect 26572 37314 26628 37326
rect 26796 37716 26852 37726
rect 26236 37268 26292 37278
rect 26236 37154 26292 37212
rect 26236 37102 26238 37154
rect 26290 37102 26292 37154
rect 26236 37090 26292 37102
rect 26684 37044 26740 37054
rect 26796 37044 26852 37660
rect 26908 37492 26964 38780
rect 26908 37426 26964 37436
rect 27020 37266 27076 40572
rect 27132 39060 27188 40910
rect 27244 39284 27300 41468
rect 27580 40516 27636 42812
rect 27580 40450 27636 40460
rect 27692 40514 27748 43036
rect 27804 42082 27860 43484
rect 28028 43428 28084 43438
rect 27916 43316 27972 43326
rect 27916 42532 27972 43260
rect 27916 42466 27972 42476
rect 28028 42530 28084 43372
rect 28140 42866 28196 44046
rect 28252 43650 28308 45164
rect 28700 44100 28756 44110
rect 28700 44006 28756 44044
rect 28252 43598 28254 43650
rect 28306 43598 28308 43650
rect 28252 43586 28308 43598
rect 28588 43538 28644 43550
rect 28588 43486 28590 43538
rect 28642 43486 28644 43538
rect 28364 43428 28420 43438
rect 28364 43334 28420 43372
rect 28140 42814 28142 42866
rect 28194 42814 28196 42866
rect 28140 42802 28196 42814
rect 28028 42478 28030 42530
rect 28082 42478 28084 42530
rect 27804 42030 27806 42082
rect 27858 42030 27860 42082
rect 27804 42018 27860 42030
rect 27916 42084 27972 42094
rect 27916 41990 27972 42028
rect 28028 41524 28084 42478
rect 28252 42530 28308 42542
rect 28252 42478 28254 42530
rect 28306 42478 28308 42530
rect 28252 42084 28308 42478
rect 28476 42532 28532 42542
rect 28476 42438 28532 42476
rect 28588 42084 28644 43486
rect 28812 42644 28868 46734
rect 28924 45892 28980 47966
rect 28924 45826 28980 45836
rect 29148 47236 29204 48748
rect 29148 45890 29204 47180
rect 29148 45838 29150 45890
rect 29202 45838 29204 45890
rect 29148 45826 29204 45838
rect 29260 45668 29316 50372
rect 29484 49028 29540 50372
rect 29596 49252 29652 51550
rect 29708 52948 29764 52958
rect 29708 51266 29764 52892
rect 29932 52612 29988 53676
rect 30044 52836 30100 53788
rect 30380 53508 30436 53518
rect 30156 52836 30212 52846
rect 30044 52780 30156 52836
rect 30156 52742 30212 52780
rect 29708 51214 29710 51266
rect 29762 51214 29764 51266
rect 29708 51202 29764 51214
rect 29820 52556 29988 52612
rect 29820 51378 29876 52556
rect 30380 52276 30436 53452
rect 30492 53284 30548 55244
rect 30604 55076 30660 56140
rect 30716 56420 30772 56430
rect 30716 55524 30772 56364
rect 31276 56420 31332 56430
rect 30828 56082 30884 56094
rect 30828 56030 30830 56082
rect 30882 56030 30884 56082
rect 30828 55748 30884 56030
rect 31276 56082 31332 56364
rect 31276 56030 31278 56082
rect 31330 56030 31332 56082
rect 31276 56018 31332 56030
rect 31388 56306 31444 56318
rect 31388 56254 31390 56306
rect 31442 56254 31444 56306
rect 31164 55860 31220 55870
rect 30828 55682 30884 55692
rect 30940 55858 31220 55860
rect 30940 55806 31166 55858
rect 31218 55806 31220 55858
rect 30940 55804 31220 55806
rect 30716 55458 30772 55468
rect 30940 55412 30996 55804
rect 31164 55794 31220 55804
rect 31052 55524 31108 55534
rect 31388 55468 31444 56254
rect 31052 55430 31108 55468
rect 30828 55356 30996 55412
rect 31276 55412 31444 55468
rect 31500 55524 31556 56702
rect 31500 55458 31556 55468
rect 31612 56532 31668 56542
rect 31612 56194 31668 56476
rect 31612 56142 31614 56194
rect 31666 56142 31668 56194
rect 30604 55010 30660 55020
rect 30716 55300 30772 55310
rect 30604 54628 30660 54638
rect 30604 54514 30660 54572
rect 30604 54462 30606 54514
rect 30658 54462 30660 54514
rect 30604 54450 30660 54462
rect 30492 53218 30548 53228
rect 30604 53732 30660 53742
rect 30492 52948 30548 52958
rect 30492 52854 30548 52892
rect 29820 51326 29822 51378
rect 29874 51326 29876 51378
rect 29596 49186 29652 49196
rect 29708 50594 29764 50606
rect 29708 50542 29710 50594
rect 29762 50542 29764 50594
rect 29708 49588 29764 50542
rect 29820 50484 29876 51326
rect 29932 52162 29988 52174
rect 29932 52110 29934 52162
rect 29986 52110 29988 52162
rect 29932 50596 29988 52110
rect 30156 52164 30212 52174
rect 30156 51828 30212 52108
rect 30268 52052 30324 52062
rect 30268 51958 30324 51996
rect 30380 52050 30436 52220
rect 30380 51998 30382 52050
rect 30434 51998 30436 52050
rect 30380 51986 30436 51998
rect 30604 52388 30660 53676
rect 30716 53730 30772 55244
rect 30828 54180 30884 55356
rect 31276 55076 31332 55412
rect 31388 55300 31444 55310
rect 31612 55300 31668 56142
rect 31388 55298 31668 55300
rect 31388 55246 31390 55298
rect 31442 55246 31668 55298
rect 31388 55244 31668 55246
rect 31388 55234 31444 55244
rect 31276 55020 31556 55076
rect 30940 54626 30996 54638
rect 30940 54574 30942 54626
rect 30994 54574 30996 54626
rect 30940 54292 30996 54574
rect 31388 54626 31444 54638
rect 31388 54574 31390 54626
rect 31442 54574 31444 54626
rect 31276 54516 31332 54526
rect 31276 54422 31332 54460
rect 30940 54226 30996 54236
rect 30828 54114 30884 54124
rect 30828 53956 30884 53966
rect 30828 53862 30884 53900
rect 31276 53956 31332 53966
rect 31276 53862 31332 53900
rect 30716 53678 30718 53730
rect 30770 53678 30772 53730
rect 30716 53666 30772 53678
rect 30940 53618 30996 53630
rect 30940 53566 30942 53618
rect 30994 53566 30996 53618
rect 30940 53284 30996 53566
rect 30940 53218 30996 53228
rect 31276 52948 31332 52958
rect 31388 52948 31444 54574
rect 31500 53842 31556 55020
rect 31500 53790 31502 53842
rect 31554 53790 31556 53842
rect 31500 53778 31556 53790
rect 31612 54516 31668 54526
rect 31612 52948 31668 54460
rect 31724 53732 31780 57486
rect 32172 57090 32228 58380
rect 32396 57650 32452 59724
rect 32508 59778 32676 59780
rect 32508 59726 32622 59778
rect 32674 59726 32676 59778
rect 32508 59724 32676 59726
rect 32508 58436 32564 59724
rect 32620 59714 32676 59724
rect 32620 58994 32676 59006
rect 32620 58942 32622 58994
rect 32674 58942 32676 58994
rect 32620 58772 32676 58942
rect 32620 58706 32676 58716
rect 32508 58370 32564 58380
rect 32732 57652 32788 59836
rect 33068 59892 33124 59902
rect 33068 59798 33124 59836
rect 38556 59890 38612 62132
rect 47740 60228 47796 63200
rect 47740 60162 47796 60172
rect 47964 60004 48020 60014
rect 38556 59838 38558 59890
rect 38610 59838 38612 59890
rect 38556 59826 38612 59838
rect 47740 60002 48020 60004
rect 47740 59950 47966 60002
rect 48018 59950 48020 60002
rect 47740 59948 48020 59950
rect 33180 59780 33236 59790
rect 33180 59686 33236 59724
rect 33740 59778 33796 59790
rect 34636 59780 34692 59790
rect 33740 59726 33742 59778
rect 33794 59726 33796 59778
rect 33740 59668 33796 59726
rect 33740 59602 33796 59612
rect 34524 59778 34692 59780
rect 34524 59726 34638 59778
rect 34690 59726 34692 59778
rect 34524 59724 34692 59726
rect 33740 59330 33796 59342
rect 33740 59278 33742 59330
rect 33794 59278 33796 59330
rect 33180 58996 33236 59006
rect 33180 58902 33236 58940
rect 33516 58994 33572 59006
rect 33516 58942 33518 58994
rect 33570 58942 33572 58994
rect 33516 58772 33572 58942
rect 33572 58716 33684 58772
rect 33516 58706 33572 58716
rect 33628 57762 33684 58716
rect 33628 57710 33630 57762
rect 33682 57710 33684 57762
rect 33628 57698 33684 57710
rect 33740 58658 33796 59278
rect 34188 59332 34244 59342
rect 34244 59276 34356 59332
rect 34188 59238 34244 59276
rect 33740 58606 33742 58658
rect 33794 58606 33796 58658
rect 32396 57598 32398 57650
rect 32450 57598 32452 57650
rect 32396 57586 32452 57598
rect 32508 57596 32788 57652
rect 32844 57652 32900 57662
rect 32172 57038 32174 57090
rect 32226 57038 32228 57090
rect 32172 57026 32228 57038
rect 32508 57090 32564 57596
rect 32508 57038 32510 57090
rect 32562 57038 32564 57090
rect 32060 56756 32116 56766
rect 32060 56306 32116 56700
rect 32060 56254 32062 56306
rect 32114 56254 32116 56306
rect 32060 56242 32116 56254
rect 32396 56644 32452 56654
rect 32396 56306 32452 56588
rect 32396 56254 32398 56306
rect 32450 56254 32452 56306
rect 32396 56242 32452 56254
rect 32172 56196 32228 56206
rect 32172 56102 32228 56140
rect 31948 56084 32004 56094
rect 31948 55990 32004 56028
rect 32172 55972 32228 55982
rect 32172 55298 32228 55916
rect 32172 55246 32174 55298
rect 32226 55246 32228 55298
rect 32172 55234 32228 55246
rect 31948 55188 32004 55198
rect 31948 55094 32004 55132
rect 32508 54852 32564 57038
rect 32732 57204 32788 57214
rect 32732 56980 32788 57148
rect 32620 56978 32788 56980
rect 32620 56926 32734 56978
rect 32786 56926 32788 56978
rect 32620 56924 32788 56926
rect 32620 55524 32676 56924
rect 32732 56914 32788 56924
rect 32844 56756 32900 57596
rect 33740 57652 33796 58606
rect 33740 57558 33796 57596
rect 34076 59108 34132 59118
rect 33404 56980 33460 56990
rect 33404 56978 33684 56980
rect 33404 56926 33406 56978
rect 33458 56926 33684 56978
rect 33404 56924 33684 56926
rect 33404 56914 33460 56924
rect 32620 55458 32676 55468
rect 32732 56700 32900 56756
rect 33068 56754 33124 56766
rect 33068 56702 33070 56754
rect 33122 56702 33124 56754
rect 32732 55748 32788 56700
rect 33068 56644 33124 56702
rect 33068 56578 33124 56588
rect 33292 56642 33348 56654
rect 33292 56590 33294 56642
rect 33346 56590 33348 56642
rect 33180 56082 33236 56094
rect 33180 56030 33182 56082
rect 33234 56030 33236 56082
rect 32732 55410 32788 55692
rect 32732 55358 32734 55410
rect 32786 55358 32788 55410
rect 32732 55346 32788 55358
rect 33068 55858 33124 55870
rect 33068 55806 33070 55858
rect 33122 55806 33124 55858
rect 33068 55412 33124 55806
rect 33068 55346 33124 55356
rect 32620 55300 32676 55310
rect 32620 55206 32676 55244
rect 33180 55300 33236 56030
rect 33292 55972 33348 56590
rect 33628 56082 33684 56924
rect 33628 56030 33630 56082
rect 33682 56030 33684 56082
rect 33628 56018 33684 56030
rect 33740 56754 33796 56766
rect 33740 56702 33742 56754
rect 33794 56702 33796 56754
rect 33292 55906 33348 55916
rect 33404 55970 33460 55982
rect 33404 55918 33406 55970
rect 33458 55918 33460 55970
rect 33180 55234 33236 55244
rect 33292 55412 33348 55422
rect 32508 54786 32564 54796
rect 32172 54628 32228 54638
rect 32172 54534 32228 54572
rect 32508 54626 32564 54638
rect 32508 54574 32510 54626
rect 32562 54574 32564 54626
rect 32508 54516 32564 54574
rect 33180 54516 33236 54526
rect 32508 54514 33236 54516
rect 32508 54462 33182 54514
rect 33234 54462 33236 54514
rect 32508 54460 33236 54462
rect 31836 54404 31892 54414
rect 31836 53842 31892 54348
rect 31836 53790 31838 53842
rect 31890 53790 31892 53842
rect 31836 53778 31892 53790
rect 31948 54180 32004 54190
rect 31724 53666 31780 53676
rect 31948 53730 32004 54124
rect 33180 53844 33236 54460
rect 33180 53778 33236 53788
rect 31948 53678 31950 53730
rect 32002 53678 32004 53730
rect 31724 53508 31780 53518
rect 31724 53414 31780 53452
rect 31276 52946 31444 52948
rect 31276 52894 31278 52946
rect 31330 52894 31444 52946
rect 31276 52892 31444 52894
rect 31500 52892 31668 52948
rect 31276 52836 31332 52892
rect 31276 52770 31332 52780
rect 31500 52834 31556 52892
rect 31500 52782 31502 52834
rect 31554 52782 31556 52834
rect 30604 52050 30660 52332
rect 30604 51998 30606 52050
rect 30658 51998 30660 52050
rect 30604 51986 30660 51998
rect 30492 51938 30548 51950
rect 30492 51886 30494 51938
rect 30546 51886 30548 51938
rect 30156 51772 30324 51828
rect 30268 51490 30324 51772
rect 30492 51604 30548 51886
rect 30492 51538 30548 51548
rect 30268 51438 30270 51490
rect 30322 51438 30324 51490
rect 29932 50530 29988 50540
rect 30156 50708 30212 50718
rect 29820 50418 29876 50428
rect 29932 50148 29988 50158
rect 29820 49700 29876 49710
rect 29820 49606 29876 49644
rect 29596 49028 29652 49038
rect 29484 49026 29652 49028
rect 29484 48974 29598 49026
rect 29650 48974 29652 49026
rect 29484 48972 29652 48974
rect 29596 48804 29652 48972
rect 29596 48738 29652 48748
rect 29708 48468 29764 49532
rect 29932 48692 29988 50092
rect 30044 49028 30100 49038
rect 30044 48934 30100 48972
rect 29932 48626 29988 48636
rect 29820 48468 29876 48478
rect 29708 48412 29820 48468
rect 29596 48356 29652 48366
rect 29372 47458 29428 47470
rect 29372 47406 29374 47458
rect 29426 47406 29428 47458
rect 29372 47348 29428 47406
rect 29372 47282 29428 47292
rect 29596 46002 29652 48300
rect 29820 48242 29876 48412
rect 29820 48190 29822 48242
rect 29874 48190 29876 48242
rect 29820 47908 29876 48190
rect 29820 47842 29876 47852
rect 30044 48356 30100 48366
rect 30156 48356 30212 50652
rect 30268 49922 30324 51438
rect 31500 51492 31556 52782
rect 31948 52836 32004 53678
rect 32620 53732 32676 53742
rect 32844 53732 32900 53742
rect 32676 53676 32788 53732
rect 32620 53666 32676 53676
rect 32396 53620 32452 53630
rect 32396 53526 32452 53564
rect 32508 53508 32564 53518
rect 32396 53060 32452 53070
rect 32284 53058 32452 53060
rect 32284 53006 32398 53058
rect 32450 53006 32452 53058
rect 32284 53004 32452 53006
rect 32172 52948 32228 52958
rect 31948 52770 32004 52780
rect 32060 52946 32228 52948
rect 32060 52894 32174 52946
rect 32226 52894 32228 52946
rect 32060 52892 32228 52894
rect 31612 52724 31668 52734
rect 31612 52630 31668 52668
rect 31612 52388 31668 52398
rect 31668 52332 31780 52388
rect 31612 52322 31668 52332
rect 31612 51492 31668 51502
rect 31500 51490 31668 51492
rect 31500 51438 31614 51490
rect 31666 51438 31668 51490
rect 31500 51436 31668 51438
rect 31612 51426 31668 51436
rect 31276 51380 31332 51390
rect 31276 51378 31444 51380
rect 31276 51326 31278 51378
rect 31330 51326 31444 51378
rect 31276 51324 31444 51326
rect 31276 51314 31332 51324
rect 30604 51154 30660 51166
rect 30604 51102 30606 51154
rect 30658 51102 30660 51154
rect 30492 50932 30548 50942
rect 30492 50428 30548 50876
rect 30604 50596 30660 51102
rect 31388 50706 31444 51324
rect 31724 51268 31780 52332
rect 31948 52276 32004 52286
rect 31836 52052 31892 52062
rect 31836 51958 31892 51996
rect 31388 50654 31390 50706
rect 31442 50654 31444 50706
rect 30940 50596 30996 50634
rect 30604 50594 30884 50596
rect 30604 50542 30606 50594
rect 30658 50542 30884 50594
rect 30604 50540 30884 50542
rect 30604 50530 30660 50540
rect 30828 50428 30884 50540
rect 30940 50530 30996 50540
rect 30492 50372 30772 50428
rect 30828 50372 31332 50428
rect 30716 50034 30772 50372
rect 30716 49982 30718 50034
rect 30770 49982 30772 50034
rect 30716 49970 30772 49982
rect 30828 50148 30884 50158
rect 30828 50034 30884 50092
rect 30828 49982 30830 50034
rect 30882 49982 30884 50034
rect 30828 49970 30884 49982
rect 31164 50148 31220 50158
rect 30268 49870 30270 49922
rect 30322 49870 30324 49922
rect 30268 49858 30324 49870
rect 30380 49924 30436 49934
rect 30044 48354 30212 48356
rect 30044 48302 30046 48354
rect 30098 48302 30212 48354
rect 30044 48300 30212 48302
rect 30044 47460 30100 48300
rect 30380 48132 30436 49868
rect 30492 49922 30548 49934
rect 30492 49870 30494 49922
rect 30546 49870 30548 49922
rect 30492 48804 30548 49870
rect 30604 49922 30660 49934
rect 30604 49870 30606 49922
rect 30658 49870 30660 49922
rect 30604 49028 30660 49870
rect 30940 49252 30996 49262
rect 30940 49158 30996 49196
rect 30604 48962 30660 48972
rect 30940 48914 30996 48926
rect 30940 48862 30942 48914
rect 30994 48862 30996 48914
rect 30940 48804 30996 48862
rect 30492 48748 30996 48804
rect 30604 48356 30660 48366
rect 30604 48262 30660 48300
rect 30380 48066 30436 48076
rect 30940 47682 30996 48748
rect 30940 47630 30942 47682
rect 30994 47630 30996 47682
rect 30940 47618 30996 47630
rect 31052 48804 31108 48814
rect 31052 48354 31108 48748
rect 31052 48302 31054 48354
rect 31106 48302 31108 48354
rect 30044 47394 30100 47404
rect 30604 47572 30660 47582
rect 30604 47458 30660 47516
rect 30604 47406 30606 47458
rect 30658 47406 30660 47458
rect 30604 47394 30660 47406
rect 31052 47460 31108 48302
rect 31164 48244 31220 50092
rect 31276 50034 31332 50372
rect 31276 49982 31278 50034
rect 31330 49982 31332 50034
rect 31276 49970 31332 49982
rect 31388 48468 31444 50654
rect 31612 51212 31780 51268
rect 31500 50596 31556 50606
rect 31500 49924 31556 50540
rect 31500 49026 31556 49868
rect 31612 49810 31668 51212
rect 31612 49758 31614 49810
rect 31666 49758 31668 49810
rect 31612 49746 31668 49758
rect 31724 50484 31780 50494
rect 31500 48974 31502 49026
rect 31554 48974 31556 49026
rect 31500 48962 31556 48974
rect 31612 48468 31668 48478
rect 31388 48466 31668 48468
rect 31388 48414 31614 48466
rect 31666 48414 31668 48466
rect 31388 48412 31668 48414
rect 31612 48402 31668 48412
rect 31276 48244 31332 48254
rect 31724 48244 31780 50428
rect 31948 49922 32004 52220
rect 32060 51378 32116 52892
rect 32172 52882 32228 52892
rect 32172 52164 32228 52174
rect 32284 52164 32340 53004
rect 32396 52994 32452 53004
rect 32508 52948 32564 53452
rect 32508 52946 32676 52948
rect 32508 52894 32510 52946
rect 32562 52894 32676 52946
rect 32508 52892 32676 52894
rect 32508 52882 32564 52892
rect 32228 52108 32340 52164
rect 32396 52836 32452 52846
rect 32172 52070 32228 52108
rect 32396 52052 32452 52780
rect 32284 51996 32452 52052
rect 32508 52162 32564 52174
rect 32508 52110 32510 52162
rect 32562 52110 32564 52162
rect 32060 51326 32062 51378
rect 32114 51326 32116 51378
rect 32060 51314 32116 51326
rect 32172 51380 32228 51390
rect 32172 51286 32228 51324
rect 31948 49870 31950 49922
rect 32002 49870 32004 49922
rect 31948 49858 32004 49870
rect 32060 50820 32116 50830
rect 31948 49700 32004 49710
rect 31164 48242 31332 48244
rect 31164 48190 31278 48242
rect 31330 48190 31332 48242
rect 31164 48188 31332 48190
rect 31276 48178 31332 48188
rect 31388 48188 31780 48244
rect 31836 49588 31892 49598
rect 31836 49252 31892 49532
rect 31052 47394 31108 47404
rect 29596 45950 29598 46002
rect 29650 45950 29652 46002
rect 29596 45938 29652 45950
rect 29708 47348 29764 47358
rect 29708 46674 29764 47292
rect 30940 47012 30996 47022
rect 29708 46622 29710 46674
rect 29762 46622 29764 46674
rect 29484 45892 29540 45902
rect 29484 45798 29540 45836
rect 29708 45890 29764 46622
rect 29708 45838 29710 45890
rect 29762 45838 29764 45890
rect 29708 45826 29764 45838
rect 29932 46676 29988 46686
rect 29932 45892 29988 46620
rect 29932 45826 29988 45836
rect 30380 46228 30436 46238
rect 30380 46002 30436 46172
rect 30380 45950 30382 46002
rect 30434 45950 30436 46002
rect 29036 45612 29316 45668
rect 29036 44660 29092 45612
rect 30268 45556 30324 45566
rect 29260 45444 29316 45454
rect 29260 45106 29316 45388
rect 29260 45054 29262 45106
rect 29314 45054 29316 45106
rect 29260 45042 29316 45054
rect 29484 45444 29540 45454
rect 29036 44604 29316 44660
rect 29260 44546 29316 44604
rect 29260 44494 29262 44546
rect 29314 44494 29316 44546
rect 29036 44436 29092 44446
rect 29092 44380 29204 44436
rect 29036 44370 29092 44380
rect 28812 42578 28868 42588
rect 29036 44100 29092 44110
rect 28252 42028 28868 42084
rect 28140 41970 28196 41982
rect 28140 41918 28142 41970
rect 28194 41918 28196 41970
rect 28140 41748 28196 41918
rect 28140 41682 28196 41692
rect 28028 41468 28420 41524
rect 27692 40462 27694 40514
rect 27746 40462 27748 40514
rect 27356 40292 27412 40302
rect 27356 40198 27412 40236
rect 27468 39620 27524 39630
rect 27468 39526 27524 39564
rect 27356 39508 27412 39518
rect 27356 39414 27412 39452
rect 27244 39228 27524 39284
rect 27244 39060 27300 39070
rect 27132 39058 27300 39060
rect 27132 39006 27246 39058
rect 27298 39006 27300 39058
rect 27132 39004 27300 39006
rect 27244 37940 27300 39004
rect 27468 38668 27524 39228
rect 27244 37874 27300 37884
rect 27356 38612 27524 38668
rect 27020 37214 27022 37266
rect 27074 37214 27076 37266
rect 27020 37202 27076 37214
rect 27132 37604 27188 37614
rect 26740 36988 26852 37044
rect 26684 36950 26740 36988
rect 26012 35758 26014 35810
rect 26066 35758 26068 35810
rect 26012 35746 26068 35758
rect 26572 36932 26628 36942
rect 25676 34862 25678 34914
rect 25730 34862 25732 34914
rect 25676 34850 25732 34862
rect 26572 35028 26628 36876
rect 26796 36820 26852 36988
rect 26908 37044 26964 37054
rect 26908 37042 27076 37044
rect 26908 36990 26910 37042
rect 26962 36990 27076 37042
rect 26908 36988 27076 36990
rect 26908 36978 26964 36988
rect 26796 36764 26964 36820
rect 25676 34244 25732 34254
rect 25564 34188 25676 34244
rect 25676 34018 25732 34188
rect 26124 34132 26180 34142
rect 26124 34130 26292 34132
rect 26124 34078 26126 34130
rect 26178 34078 26292 34130
rect 26124 34076 26292 34078
rect 26124 34066 26180 34076
rect 25676 33966 25678 34018
rect 25730 33966 25732 34018
rect 25676 33954 25732 33966
rect 25788 34020 25844 34030
rect 25452 33572 25508 33582
rect 25004 33030 25060 33068
rect 25116 33516 25284 33572
rect 25340 33570 25508 33572
rect 25340 33518 25454 33570
rect 25506 33518 25508 33570
rect 25340 33516 25508 33518
rect 25116 32452 25172 33516
rect 25228 33346 25284 33358
rect 25228 33294 25230 33346
rect 25282 33294 25284 33346
rect 25228 32676 25284 33294
rect 25228 32610 25284 32620
rect 25116 32396 25284 32452
rect 25228 31778 25284 32396
rect 25228 31726 25230 31778
rect 25282 31726 25284 31778
rect 25228 31714 25284 31726
rect 25228 30324 25284 30334
rect 25228 30230 25284 30268
rect 25340 30100 25396 33516
rect 25452 33506 25508 33516
rect 25788 33234 25844 33964
rect 25788 33182 25790 33234
rect 25842 33182 25844 33234
rect 25564 33122 25620 33134
rect 25564 33070 25566 33122
rect 25618 33070 25620 33122
rect 25564 31892 25620 33070
rect 25564 31826 25620 31836
rect 25788 32788 25844 33182
rect 25788 31444 25844 32732
rect 26012 33236 26068 33246
rect 26012 32116 26068 33180
rect 26012 32050 26068 32060
rect 26236 32562 26292 34076
rect 26460 34018 26516 34030
rect 26460 33966 26462 34018
rect 26514 33966 26516 34018
rect 26460 33684 26516 33966
rect 26460 33618 26516 33628
rect 26572 32676 26628 34972
rect 26684 33906 26740 33918
rect 26684 33854 26686 33906
rect 26738 33854 26740 33906
rect 26684 33460 26740 33854
rect 26684 33394 26740 33404
rect 26236 32510 26238 32562
rect 26290 32510 26292 32562
rect 26236 31892 26292 32510
rect 26460 32620 26628 32676
rect 26460 32562 26516 32620
rect 26460 32510 26462 32562
rect 26514 32510 26516 32562
rect 26460 32498 26516 32510
rect 26236 31826 26292 31836
rect 26684 32450 26740 32462
rect 26684 32398 26686 32450
rect 26738 32398 26740 32450
rect 25900 31668 25956 31678
rect 25900 31574 25956 31612
rect 26012 31556 26068 31566
rect 25788 31388 25956 31444
rect 25788 30994 25844 31006
rect 25788 30942 25790 30994
rect 25842 30942 25844 30994
rect 25676 30772 25732 30782
rect 25676 30678 25732 30716
rect 25228 30044 25396 30100
rect 25452 30324 25508 30334
rect 25004 29428 25060 29438
rect 25004 28866 25060 29372
rect 25004 28814 25006 28866
rect 25058 28814 25060 28866
rect 25004 28802 25060 28814
rect 25228 28082 25284 30044
rect 25452 29538 25508 30268
rect 25564 30212 25620 30222
rect 25564 29764 25620 30156
rect 25564 29650 25620 29708
rect 25564 29598 25566 29650
rect 25618 29598 25620 29650
rect 25564 29586 25620 29598
rect 25676 29986 25732 29998
rect 25676 29934 25678 29986
rect 25730 29934 25732 29986
rect 25452 29486 25454 29538
rect 25506 29486 25508 29538
rect 25452 29474 25508 29486
rect 25564 29428 25620 29438
rect 25676 29428 25732 29934
rect 25788 29650 25844 30942
rect 25788 29598 25790 29650
rect 25842 29598 25844 29650
rect 25788 29586 25844 29598
rect 25620 29372 25732 29428
rect 25564 29362 25620 29372
rect 25900 29204 25956 31388
rect 26012 30324 26068 31500
rect 26124 30884 26180 30894
rect 26124 30882 26292 30884
rect 26124 30830 26126 30882
rect 26178 30830 26292 30882
rect 26124 30828 26292 30830
rect 26124 30818 26180 30828
rect 26012 30210 26068 30268
rect 26012 30158 26014 30210
rect 26066 30158 26068 30210
rect 26012 30146 26068 30158
rect 26236 30100 26292 30828
rect 25452 29148 25956 29204
rect 26124 29986 26180 29998
rect 26124 29934 26126 29986
rect 26178 29934 26180 29986
rect 25452 28084 25508 29148
rect 26124 29092 26180 29934
rect 26236 29426 26292 30044
rect 26236 29374 26238 29426
rect 26290 29374 26292 29426
rect 26236 29362 26292 29374
rect 26348 29986 26404 29998
rect 26348 29934 26350 29986
rect 26402 29934 26404 29986
rect 26348 29428 26404 29934
rect 26348 29362 26404 29372
rect 26124 29026 26180 29036
rect 26236 28756 26292 28766
rect 26124 28644 26180 28654
rect 25676 28532 25732 28542
rect 25228 28030 25230 28082
rect 25282 28030 25284 28082
rect 25228 28018 25284 28030
rect 25340 28028 25508 28084
rect 25564 28476 25676 28532
rect 25340 27858 25396 28028
rect 25340 27806 25342 27858
rect 25394 27806 25396 27858
rect 25340 27794 25396 27806
rect 25452 27860 25508 27870
rect 25452 27636 25508 27804
rect 25116 27634 25508 27636
rect 25116 27582 25454 27634
rect 25506 27582 25508 27634
rect 25116 27580 25508 27582
rect 25116 27186 25172 27580
rect 25452 27570 25508 27580
rect 25116 27134 25118 27186
rect 25170 27134 25172 27186
rect 25116 27122 25172 27134
rect 25228 27188 25284 27198
rect 25004 27074 25060 27086
rect 25004 27022 25006 27074
rect 25058 27022 25060 27074
rect 25004 26964 25060 27022
rect 25228 26964 25284 27132
rect 25004 26908 25284 26964
rect 24892 26348 25060 26404
rect 23548 25506 23716 25508
rect 23548 25454 23550 25506
rect 23602 25454 23716 25506
rect 23548 25452 23716 25454
rect 23772 25730 24276 25732
rect 23772 25678 24222 25730
rect 24274 25678 24276 25730
rect 23772 25676 24276 25678
rect 22316 22594 22372 24556
rect 22428 24052 22484 24062
rect 22428 23154 22484 23996
rect 22764 23604 22820 24556
rect 23100 24498 23156 24510
rect 23100 24446 23102 24498
rect 23154 24446 23156 24498
rect 22988 24164 23044 24174
rect 22428 23102 22430 23154
rect 22482 23102 22484 23154
rect 22428 23090 22484 23102
rect 22540 23548 22820 23604
rect 22876 23828 22932 23838
rect 22316 22542 22318 22594
rect 22370 22542 22372 22594
rect 22316 22530 22372 22542
rect 22428 22372 22484 22382
rect 22428 22278 22484 22316
rect 22316 22260 22372 22270
rect 22316 22166 22372 22204
rect 22316 21588 22372 21598
rect 22316 21494 22372 21532
rect 22428 21140 22484 21150
rect 22540 21140 22596 23548
rect 22876 23492 22932 23772
rect 22652 23436 22932 23492
rect 22652 21810 22708 23436
rect 22988 23154 23044 24108
rect 23100 24052 23156 24446
rect 23436 24498 23492 24510
rect 23436 24446 23438 24498
rect 23490 24446 23492 24498
rect 23324 24052 23380 24062
rect 23100 23986 23156 23996
rect 23212 23996 23324 24052
rect 23100 23714 23156 23726
rect 23100 23662 23102 23714
rect 23154 23662 23156 23714
rect 23100 23604 23156 23662
rect 23100 23538 23156 23548
rect 23212 23380 23268 23996
rect 23324 23986 23380 23996
rect 23324 23716 23380 23726
rect 23436 23716 23492 24446
rect 23548 24500 23604 25452
rect 23660 24724 23716 24734
rect 23660 24630 23716 24668
rect 23660 24500 23716 24510
rect 23548 24444 23660 24500
rect 23660 24434 23716 24444
rect 23660 24052 23716 24062
rect 23380 23660 23492 23716
rect 23548 23828 23604 23838
rect 23324 23650 23380 23660
rect 23548 23604 23604 23772
rect 23436 23548 23604 23604
rect 22988 23102 22990 23154
rect 23042 23102 23044 23154
rect 22988 23090 23044 23102
rect 23100 23324 23268 23380
rect 23324 23492 23380 23502
rect 22652 21758 22654 21810
rect 22706 21758 22708 21810
rect 22652 21746 22708 21758
rect 23100 21812 23156 23324
rect 23212 23156 23268 23166
rect 23212 23062 23268 23100
rect 23324 22372 23380 23436
rect 23436 23266 23492 23548
rect 23436 23214 23438 23266
rect 23490 23214 23492 23266
rect 23436 23202 23492 23214
rect 23660 23266 23716 23996
rect 23660 23214 23662 23266
rect 23714 23214 23716 23266
rect 23660 23202 23716 23214
rect 23772 23044 23828 25676
rect 24220 25666 24276 25676
rect 24444 26066 24612 26068
rect 24444 26014 24558 26066
rect 24610 26014 24612 26066
rect 24444 26012 24612 26014
rect 23884 25396 23940 25406
rect 24332 25396 24388 25406
rect 23884 25394 24052 25396
rect 23884 25342 23886 25394
rect 23938 25342 24052 25394
rect 23884 25340 24052 25342
rect 23884 25330 23940 25340
rect 23324 22306 23380 22316
rect 23548 22988 23828 23044
rect 23884 23604 23940 23614
rect 23100 21746 23156 21756
rect 23436 22146 23492 22158
rect 23436 22094 23438 22146
rect 23490 22094 23492 22146
rect 22876 21700 22932 21710
rect 22876 21586 22932 21644
rect 23436 21700 23492 22094
rect 22876 21534 22878 21586
rect 22930 21534 22932 21586
rect 22484 21084 22596 21140
rect 22764 21474 22820 21486
rect 22764 21422 22766 21474
rect 22818 21422 22820 21474
rect 22428 21074 22484 21084
rect 22764 21028 22820 21422
rect 22540 20972 22820 21028
rect 22540 20914 22596 20972
rect 22540 20862 22542 20914
rect 22594 20862 22596 20914
rect 22540 20850 22596 20862
rect 22204 20636 22596 20692
rect 22092 20132 22148 20142
rect 22092 20038 22148 20076
rect 21868 17668 21924 19964
rect 21980 19122 22036 19134
rect 21980 19070 21982 19122
rect 22034 19070 22036 19122
rect 21980 18452 22036 19070
rect 22316 19124 22372 19134
rect 22316 19030 22372 19068
rect 22428 18564 22484 18574
rect 22428 18470 22484 18508
rect 21980 18386 22036 18396
rect 22204 18452 22260 18462
rect 22540 18452 22596 20636
rect 22764 18452 22820 18462
rect 22540 18450 22820 18452
rect 22540 18398 22766 18450
rect 22818 18398 22820 18450
rect 22540 18396 22820 18398
rect 22204 18358 22260 18396
rect 21980 17668 22036 17678
rect 21868 17666 22036 17668
rect 21868 17614 21982 17666
rect 22034 17614 22036 17666
rect 21868 17612 22036 17614
rect 21980 17602 22036 17612
rect 21308 17554 21588 17556
rect 21308 17502 21310 17554
rect 21362 17502 21588 17554
rect 21308 17500 21588 17502
rect 21644 17554 21700 17566
rect 21644 17502 21646 17554
rect 21698 17502 21700 17554
rect 21308 17490 21364 17500
rect 21644 17332 21700 17502
rect 20748 17276 21700 17332
rect 20636 17164 20916 17220
rect 20524 16830 20526 16882
rect 20578 16830 20580 16882
rect 20524 16818 20580 16830
rect 20300 16606 20302 16658
rect 20354 16606 20356 16658
rect 20300 16594 20356 16606
rect 20636 16212 20692 16222
rect 20636 16118 20692 16156
rect 20300 16100 20356 16110
rect 20300 16006 20356 16044
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15426 20244 15438
rect 20188 15374 20190 15426
rect 20242 15374 20244 15426
rect 20188 15148 20244 15374
rect 20076 15092 20244 15148
rect 20524 15316 20580 15326
rect 20076 14980 20132 15092
rect 20076 14914 20132 14924
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13346 19684 13356
rect 19740 13858 19796 13870
rect 19740 13806 19742 13858
rect 19794 13806 19796 13858
rect 19740 13300 19796 13806
rect 19740 13234 19796 13244
rect 20412 13188 20468 13198
rect 18956 13076 19012 13086
rect 19852 13076 19908 13086
rect 18508 13020 18900 13076
rect 18284 12402 18452 12404
rect 18284 12350 18398 12402
rect 18450 12350 18452 12402
rect 18284 12348 18452 12350
rect 18060 11452 18228 11508
rect 17612 10724 17668 10734
rect 17612 10630 17668 10668
rect 17500 10444 17668 10500
rect 17164 9538 17220 9548
rect 17500 10276 17556 10286
rect 17276 9044 17332 9054
rect 16716 7250 16884 7252
rect 16716 7198 16718 7250
rect 16770 7198 16884 7250
rect 16716 7196 16884 7198
rect 16940 9042 17332 9044
rect 16940 8990 17278 9042
rect 17330 8990 17332 9042
rect 16940 8988 17332 8990
rect 16716 7186 16772 7196
rect 16604 6638 16606 6690
rect 16658 6638 16660 6690
rect 16604 6626 16660 6638
rect 16940 6690 16996 8988
rect 17276 8978 17332 8988
rect 17388 8260 17444 8270
rect 17388 8166 17444 8204
rect 17388 7700 17444 7710
rect 17388 7252 17444 7644
rect 17500 7476 17556 10220
rect 17612 7700 17668 10444
rect 17724 9154 17780 11452
rect 17836 11442 17892 11452
rect 17948 11396 18004 11406
rect 17948 11302 18004 11340
rect 18172 10948 18228 11452
rect 17724 9102 17726 9154
rect 17778 9102 17780 9154
rect 17724 9090 17780 9102
rect 17836 10892 18228 10948
rect 17612 7634 17668 7644
rect 17500 7420 17668 7476
rect 17500 7252 17556 7262
rect 17388 7250 17556 7252
rect 17388 7198 17502 7250
rect 17554 7198 17556 7250
rect 17388 7196 17556 7198
rect 17500 7140 17556 7196
rect 17500 7074 17556 7084
rect 16940 6638 16942 6690
rect 16994 6638 16996 6690
rect 16940 6626 16996 6638
rect 16492 6066 16548 6076
rect 16716 6466 16772 6478
rect 16716 6414 16718 6466
rect 16770 6414 16772 6466
rect 16716 5908 16772 6414
rect 17500 6468 17556 6478
rect 17500 6374 17556 6412
rect 16828 6132 16884 6142
rect 16828 6038 16884 6076
rect 17500 6132 17556 6142
rect 17612 6132 17668 7420
rect 17836 6692 17892 10892
rect 18060 10722 18116 10734
rect 18060 10670 18062 10722
rect 18114 10670 18116 10722
rect 18060 10276 18116 10670
rect 18284 10610 18340 12348
rect 18396 12338 18452 12348
rect 18508 12850 18564 12862
rect 18508 12798 18510 12850
rect 18562 12798 18564 12850
rect 18508 12292 18564 12798
rect 18732 12850 18788 12862
rect 18732 12798 18734 12850
rect 18786 12798 18788 12850
rect 18732 12740 18788 12798
rect 18732 12674 18788 12684
rect 18508 12226 18564 12236
rect 18620 12290 18676 12302
rect 18620 12238 18622 12290
rect 18674 12238 18676 12290
rect 18620 11844 18676 12238
rect 18284 10558 18286 10610
rect 18338 10558 18340 10610
rect 18284 10500 18340 10558
rect 18284 10434 18340 10444
rect 18396 11788 18676 11844
rect 18732 12290 18788 12302
rect 18732 12238 18734 12290
rect 18786 12238 18788 12290
rect 18396 10276 18452 11788
rect 18620 11282 18676 11294
rect 18620 11230 18622 11282
rect 18674 11230 18676 11282
rect 18620 11060 18676 11230
rect 18620 10994 18676 11004
rect 18732 10612 18788 12238
rect 18060 10220 18452 10276
rect 18508 10556 18788 10612
rect 17948 9826 18004 9838
rect 17948 9774 17950 9826
rect 18002 9774 18004 9826
rect 17948 9268 18004 9774
rect 18060 9828 18116 10220
rect 18060 9762 18116 9772
rect 18172 9716 18228 9726
rect 18508 9716 18564 10556
rect 18620 10388 18676 10398
rect 18732 10388 18788 10398
rect 18620 10386 18732 10388
rect 18620 10334 18622 10386
rect 18674 10334 18732 10386
rect 18620 10332 18732 10334
rect 18620 10322 18676 10332
rect 18172 9714 18564 9716
rect 18172 9662 18174 9714
rect 18226 9662 18564 9714
rect 18172 9660 18564 9662
rect 18060 9268 18116 9278
rect 17948 9212 18060 9268
rect 17948 8372 18004 9212
rect 18060 9202 18116 9212
rect 18172 8482 18228 9660
rect 18732 8818 18788 10332
rect 18844 9380 18900 13020
rect 18956 13074 19908 13076
rect 18956 13022 18958 13074
rect 19010 13022 19854 13074
rect 19906 13022 19908 13074
rect 18956 13020 19908 13022
rect 18956 13010 19012 13020
rect 19852 13010 19908 13020
rect 19068 12852 19124 12862
rect 18956 12850 19124 12852
rect 18956 12798 19070 12850
rect 19122 12798 19124 12850
rect 18956 12796 19124 12798
rect 18956 12180 19012 12796
rect 19068 12786 19124 12796
rect 19516 12852 19572 12862
rect 19516 12758 19572 12796
rect 20412 12850 20468 13132
rect 20412 12798 20414 12850
rect 20466 12798 20468 12850
rect 20412 12786 20468 12798
rect 20188 12740 20244 12750
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19628 12292 19684 12302
rect 19516 12290 19684 12292
rect 19516 12238 19630 12290
rect 19682 12238 19684 12290
rect 19516 12236 19684 12238
rect 18956 11620 19012 12124
rect 19068 12178 19124 12190
rect 19068 12126 19070 12178
rect 19122 12126 19124 12178
rect 19068 11844 19124 12126
rect 19180 12068 19236 12078
rect 19516 12068 19572 12236
rect 19628 12226 19684 12236
rect 20188 12290 20244 12684
rect 20524 12740 20580 15260
rect 20860 15148 20916 17164
rect 21644 16996 21700 17006
rect 21532 16884 21588 16894
rect 21308 16100 21364 16110
rect 21308 16006 21364 16044
rect 21532 15652 21588 16828
rect 21644 15764 21700 16940
rect 21980 16882 22036 16894
rect 21980 16830 21982 16882
rect 22034 16830 22036 16882
rect 21868 16772 21924 16782
rect 21756 15988 21812 15998
rect 21868 15988 21924 16716
rect 21756 15986 21924 15988
rect 21756 15934 21758 15986
rect 21810 15934 21924 15986
rect 21756 15932 21924 15934
rect 21756 15922 21812 15932
rect 21868 15876 21924 15932
rect 21868 15810 21924 15820
rect 21980 16212 22036 16830
rect 22652 16324 22708 18396
rect 22764 18386 22820 18396
rect 22764 17554 22820 17566
rect 22764 17502 22766 17554
rect 22818 17502 22820 17554
rect 22764 16772 22820 17502
rect 22876 16996 22932 21534
rect 23324 21586 23380 21598
rect 23324 21534 23326 21586
rect 23378 21534 23380 21586
rect 23324 20244 23380 21534
rect 23436 21476 23492 21644
rect 23548 21698 23604 22988
rect 23884 21810 23940 23548
rect 23884 21758 23886 21810
rect 23938 21758 23940 21810
rect 23884 21746 23940 21758
rect 23548 21646 23550 21698
rect 23602 21646 23604 21698
rect 23548 21634 23604 21646
rect 23660 21700 23716 21710
rect 23660 21698 23828 21700
rect 23660 21646 23662 21698
rect 23714 21646 23828 21698
rect 23660 21644 23828 21646
rect 23660 21634 23716 21644
rect 23436 21410 23492 21420
rect 23772 21364 23828 21644
rect 23772 21298 23828 21308
rect 23324 20178 23380 20188
rect 23436 20356 23492 20366
rect 23436 19684 23492 20300
rect 23212 19628 23492 19684
rect 23212 19346 23268 19628
rect 23212 19294 23214 19346
rect 23266 19294 23268 19346
rect 23212 19282 23268 19294
rect 23772 19122 23828 19134
rect 23772 19070 23774 19122
rect 23826 19070 23828 19122
rect 23660 19012 23716 19022
rect 23324 18338 23380 18350
rect 23324 18286 23326 18338
rect 23378 18286 23380 18338
rect 23212 16996 23268 17006
rect 22876 16940 23212 16996
rect 22764 16706 22820 16716
rect 22764 16324 22820 16334
rect 22652 16268 22764 16324
rect 22764 16258 22820 16268
rect 21644 15708 21812 15764
rect 21532 15596 21700 15652
rect 21532 15426 21588 15438
rect 21532 15374 21534 15426
rect 21586 15374 21588 15426
rect 21420 15314 21476 15326
rect 21420 15262 21422 15314
rect 21474 15262 21476 15314
rect 20860 15092 21252 15148
rect 20636 14532 20692 14542
rect 20636 14306 20692 14476
rect 20636 14254 20638 14306
rect 20690 14254 20692 14306
rect 20636 13860 20692 14254
rect 20636 13794 20692 13804
rect 20636 12964 20692 12974
rect 21084 12964 21140 12974
rect 20636 12962 21084 12964
rect 20636 12910 20638 12962
rect 20690 12910 21084 12962
rect 20636 12908 21084 12910
rect 20636 12898 20692 12908
rect 20524 12674 20580 12684
rect 20188 12238 20190 12290
rect 20242 12238 20244 12290
rect 19180 12066 19572 12068
rect 19180 12014 19182 12066
rect 19234 12014 19572 12066
rect 19180 12012 19572 12014
rect 19740 12178 19796 12190
rect 19740 12126 19742 12178
rect 19794 12126 19796 12178
rect 19180 12002 19236 12012
rect 19628 11954 19684 11966
rect 19628 11902 19630 11954
rect 19682 11902 19684 11954
rect 19068 11788 19460 11844
rect 18956 11564 19124 11620
rect 19068 11394 19124 11564
rect 19068 11342 19070 11394
rect 19122 11342 19124 11394
rect 18956 11284 19012 11294
rect 18956 11190 19012 11228
rect 18956 10610 19012 10622
rect 18956 10558 18958 10610
rect 19010 10558 19012 10610
rect 18956 10052 19012 10558
rect 19068 10388 19124 11342
rect 19292 10500 19348 10510
rect 19180 10388 19236 10398
rect 19068 10386 19236 10388
rect 19068 10334 19182 10386
rect 19234 10334 19236 10386
rect 19068 10332 19236 10334
rect 19180 10322 19236 10332
rect 19292 10052 19348 10444
rect 18956 9986 19012 9996
rect 19180 9996 19348 10052
rect 19180 9938 19236 9996
rect 19180 9886 19182 9938
rect 19234 9886 19236 9938
rect 19180 9874 19236 9886
rect 19292 9828 19348 9838
rect 19404 9828 19460 11788
rect 19516 11396 19572 11406
rect 19516 11302 19572 11340
rect 19628 10836 19684 11902
rect 19740 11172 19796 12126
rect 20076 12180 20132 12190
rect 20076 12086 20132 12124
rect 20188 11396 20244 12238
rect 20300 12292 20356 12302
rect 20860 12292 20916 12302
rect 20356 12236 20468 12292
rect 20300 12226 20356 12236
rect 20188 11330 20244 11340
rect 20300 11394 20356 11406
rect 20300 11342 20302 11394
rect 20354 11342 20356 11394
rect 19740 11116 20244 11172
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 10836 20244 11116
rect 19628 10770 19684 10780
rect 20076 10780 20244 10836
rect 19516 10610 19572 10622
rect 19516 10558 19518 10610
rect 19570 10558 19572 10610
rect 19516 10388 19572 10558
rect 19516 10322 19572 10332
rect 19740 10276 19796 10286
rect 19628 10220 19740 10276
rect 19404 9772 19572 9828
rect 18844 9324 19236 9380
rect 18844 9156 18900 9166
rect 18844 8930 18900 9100
rect 18844 8878 18846 8930
rect 18898 8878 18900 8930
rect 18844 8866 18900 8878
rect 19068 9154 19124 9166
rect 19068 9102 19070 9154
rect 19122 9102 19124 9154
rect 19068 9044 19124 9102
rect 18732 8766 18734 8818
rect 18786 8766 18788 8818
rect 18732 8754 18788 8766
rect 18172 8430 18174 8482
rect 18226 8430 18228 8482
rect 18172 8418 18228 8430
rect 18620 8596 18676 8606
rect 17948 8306 18004 8316
rect 18620 8146 18676 8540
rect 18620 8094 18622 8146
rect 18674 8094 18676 8146
rect 18620 8082 18676 8094
rect 18732 7700 18788 7710
rect 18732 7588 18788 7644
rect 17836 6626 17892 6636
rect 18508 7586 18788 7588
rect 18508 7534 18734 7586
rect 18786 7534 18788 7586
rect 18508 7532 18788 7534
rect 18508 6580 18564 7532
rect 18732 7522 18788 7532
rect 18956 6692 19012 6702
rect 18508 6578 18900 6580
rect 18508 6526 18510 6578
rect 18562 6526 18900 6578
rect 18508 6524 18900 6526
rect 18508 6514 18564 6524
rect 17500 6130 17668 6132
rect 17500 6078 17502 6130
rect 17554 6078 17668 6130
rect 17500 6076 17668 6078
rect 18844 6130 18900 6524
rect 18844 6078 18846 6130
rect 18898 6078 18900 6130
rect 17500 6066 17556 6076
rect 18844 6066 18900 6078
rect 16716 5842 16772 5852
rect 16380 5796 16436 5806
rect 16156 5740 16380 5796
rect 16044 5182 16046 5234
rect 16098 5182 16100 5234
rect 16044 5170 16100 5182
rect 16380 5234 16436 5740
rect 16380 5182 16382 5234
rect 16434 5182 16436 5234
rect 16380 5170 16436 5182
rect 18844 5236 18900 5246
rect 18956 5236 19012 6636
rect 19068 5908 19124 8988
rect 19180 8036 19236 9324
rect 19292 8258 19348 9772
rect 19516 9044 19572 9772
rect 19628 9268 19684 10220
rect 19740 10210 19796 10220
rect 19740 10050 19796 10062
rect 19740 9998 19742 10050
rect 19794 9998 19796 10050
rect 19740 9604 19796 9998
rect 20076 9604 20132 10780
rect 20300 10052 20356 11342
rect 20412 10724 20468 12236
rect 20748 12180 20804 12190
rect 20748 12086 20804 12124
rect 20860 12066 20916 12236
rect 20860 12014 20862 12066
rect 20914 12014 20916 12066
rect 20860 12002 20916 12014
rect 21084 12178 21140 12908
rect 21084 12126 21086 12178
rect 21138 12126 21140 12178
rect 20524 11620 20580 11630
rect 20524 10836 20580 11564
rect 20748 11284 20804 11294
rect 20748 11282 21028 11284
rect 20748 11230 20750 11282
rect 20802 11230 21028 11282
rect 20748 11228 21028 11230
rect 20748 11218 20804 11228
rect 20636 11172 20692 11182
rect 20636 11078 20692 11116
rect 20524 10780 20692 10836
rect 20412 10668 20580 10724
rect 20300 9986 20356 9996
rect 20412 10498 20468 10510
rect 20412 10446 20414 10498
rect 20466 10446 20468 10498
rect 20412 9716 20468 10446
rect 20300 9604 20356 9614
rect 20076 9548 20244 9604
rect 19740 9538 19796 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9268 20244 9548
rect 19628 9212 19908 9268
rect 19740 9044 19796 9054
rect 19516 8988 19740 9044
rect 19740 8950 19796 8988
rect 19292 8206 19294 8258
rect 19346 8206 19348 8258
rect 19292 8194 19348 8206
rect 19852 8258 19908 9212
rect 20076 9212 20244 9268
rect 19852 8206 19854 8258
rect 19906 8206 19908 8258
rect 19852 8194 19908 8206
rect 19964 9044 20020 9054
rect 19964 8260 20020 8988
rect 20076 8428 20132 9212
rect 20300 8708 20356 9548
rect 20412 9156 20468 9660
rect 20412 9090 20468 9100
rect 20188 8652 20356 8708
rect 20188 8596 20244 8652
rect 20524 8596 20580 10668
rect 20636 9828 20692 10780
rect 20636 9044 20692 9772
rect 20636 8978 20692 8988
rect 20860 10610 20916 10622
rect 20860 10558 20862 10610
rect 20914 10558 20916 10610
rect 20860 9268 20916 10558
rect 20972 9268 21028 11228
rect 21084 10836 21140 12126
rect 21196 11060 21252 15092
rect 21308 14868 21364 14878
rect 21308 14530 21364 14812
rect 21308 14478 21310 14530
rect 21362 14478 21364 14530
rect 21308 14466 21364 14478
rect 21420 14532 21476 15262
rect 21420 14466 21476 14476
rect 21420 14308 21476 14318
rect 21420 14214 21476 14252
rect 21420 13748 21476 13758
rect 21308 13300 21364 13310
rect 21308 13074 21364 13244
rect 21308 13022 21310 13074
rect 21362 13022 21364 13074
rect 21308 13010 21364 13022
rect 21420 12962 21476 13692
rect 21532 13636 21588 15374
rect 21644 14530 21700 15596
rect 21644 14478 21646 14530
rect 21698 14478 21700 14530
rect 21644 14466 21700 14478
rect 21756 13970 21812 15708
rect 21868 15204 21924 15214
rect 21868 14642 21924 15148
rect 21868 14590 21870 14642
rect 21922 14590 21924 14642
rect 21868 14578 21924 14590
rect 21756 13918 21758 13970
rect 21810 13918 21812 13970
rect 21756 13906 21812 13918
rect 21980 13636 22036 16156
rect 23100 16100 23156 16110
rect 22428 16098 23156 16100
rect 22428 16046 23102 16098
rect 23154 16046 23156 16098
rect 22428 16044 23156 16046
rect 22092 15092 22148 15102
rect 22092 14530 22148 15036
rect 22092 14478 22094 14530
rect 22146 14478 22148 14530
rect 22092 13746 22148 14478
rect 22092 13694 22094 13746
rect 22146 13694 22148 13746
rect 22092 13682 22148 13694
rect 22204 15090 22260 15102
rect 22204 15038 22206 15090
rect 22258 15038 22260 15090
rect 22204 14980 22260 15038
rect 21532 13542 21588 13580
rect 21868 13580 22036 13636
rect 21756 13076 21812 13086
rect 21420 12910 21422 12962
rect 21474 12910 21476 12962
rect 21420 12898 21476 12910
rect 21644 12962 21700 12974
rect 21644 12910 21646 12962
rect 21698 12910 21700 12962
rect 21644 12852 21700 12910
rect 21644 12786 21700 12796
rect 21308 12740 21364 12750
rect 21308 12068 21364 12684
rect 21308 12012 21476 12068
rect 21420 11788 21476 12012
rect 21420 11732 21700 11788
rect 21196 10994 21252 11004
rect 21308 11170 21364 11182
rect 21308 11118 21310 11170
rect 21362 11118 21364 11170
rect 21196 10836 21252 10846
rect 21084 10834 21252 10836
rect 21084 10782 21198 10834
rect 21250 10782 21252 10834
rect 21084 10780 21252 10782
rect 21196 10770 21252 10780
rect 21308 10276 21364 11118
rect 21532 10836 21588 10846
rect 21644 10836 21700 11732
rect 21532 10834 21700 10836
rect 21532 10782 21534 10834
rect 21586 10782 21700 10834
rect 21532 10780 21700 10782
rect 21532 10770 21588 10780
rect 21308 10210 21364 10220
rect 21756 10050 21812 13020
rect 21868 12850 21924 13580
rect 22204 13524 22260 14924
rect 22428 14754 22484 16044
rect 23100 16034 23156 16044
rect 22540 15876 22596 15886
rect 23212 15876 23268 16940
rect 22540 15538 22596 15820
rect 22540 15486 22542 15538
rect 22594 15486 22596 15538
rect 22540 15474 22596 15486
rect 22988 15820 23268 15876
rect 22652 15204 22708 15214
rect 22988 15148 23044 15820
rect 23324 15652 23380 18286
rect 23660 17220 23716 18956
rect 23772 18340 23828 19070
rect 23996 18452 24052 25340
rect 24220 25394 24388 25396
rect 24220 25342 24334 25394
rect 24386 25342 24388 25394
rect 24220 25340 24388 25342
rect 24108 23938 24164 23950
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 24108 23716 24164 23886
rect 24108 23650 24164 23660
rect 24108 23380 24164 23390
rect 24108 21252 24164 23324
rect 24220 21700 24276 25340
rect 24332 25330 24388 25340
rect 24444 24722 24500 26012
rect 24556 26002 24612 26012
rect 24892 26180 24948 26190
rect 24668 25956 24724 25966
rect 24444 24670 24446 24722
rect 24498 24670 24500 24722
rect 24444 24658 24500 24670
rect 24556 25620 24612 25630
rect 24556 25284 24612 25564
rect 24332 24612 24388 24622
rect 24332 24052 24388 24556
rect 24332 23958 24388 23996
rect 24444 23940 24500 23950
rect 24444 23846 24500 23884
rect 24556 23492 24612 25228
rect 24668 24946 24724 25900
rect 24668 24894 24670 24946
rect 24722 24894 24724 24946
rect 24668 24882 24724 24894
rect 24780 25506 24836 25518
rect 24780 25454 24782 25506
rect 24834 25454 24836 25506
rect 24668 24164 24724 24174
rect 24780 24164 24836 25454
rect 24724 24108 24836 24164
rect 24668 23938 24724 24108
rect 24892 24052 24948 26124
rect 24668 23886 24670 23938
rect 24722 23886 24724 23938
rect 24668 23874 24724 23886
rect 24780 23996 24948 24052
rect 24220 21634 24276 21644
rect 24332 23436 24612 23492
rect 24220 21476 24276 21486
rect 24332 21476 24388 23436
rect 24780 23380 24836 23996
rect 24892 23828 24948 23838
rect 24892 23734 24948 23772
rect 24780 23314 24836 23324
rect 24556 23156 24612 23166
rect 24612 23100 24836 23156
rect 24556 23062 24612 23100
rect 24444 23042 24500 23054
rect 24444 22990 24446 23042
rect 24498 22990 24500 23042
rect 24444 22372 24500 22990
rect 24780 22594 24836 23100
rect 24780 22542 24782 22594
rect 24834 22542 24836 22594
rect 24780 22530 24836 22542
rect 24444 22306 24500 22316
rect 25004 22148 25060 26348
rect 25228 25844 25284 26908
rect 25340 27076 25396 27086
rect 25340 26852 25396 27020
rect 25564 26964 25620 28476
rect 25676 28466 25732 28476
rect 26012 27972 26068 27982
rect 25676 27858 25732 27870
rect 25676 27806 25678 27858
rect 25730 27806 25732 27858
rect 25676 27748 25732 27806
rect 25732 27692 25956 27748
rect 25676 27682 25732 27692
rect 25900 27074 25956 27692
rect 26012 27188 26068 27916
rect 26124 27412 26180 28588
rect 26236 28530 26292 28700
rect 26236 28478 26238 28530
rect 26290 28478 26292 28530
rect 26236 27972 26292 28478
rect 26236 27906 26292 27916
rect 26348 27970 26404 27982
rect 26348 27918 26350 27970
rect 26402 27918 26404 27970
rect 26348 27748 26404 27918
rect 26348 27682 26404 27692
rect 26572 27858 26628 27870
rect 26572 27806 26574 27858
rect 26626 27806 26628 27858
rect 26124 27346 26180 27356
rect 26572 27188 26628 27806
rect 26684 27860 26740 32398
rect 26908 31220 26964 36764
rect 27020 36596 27076 36988
rect 27020 36530 27076 36540
rect 27132 34914 27188 37548
rect 27356 36820 27412 38612
rect 27692 38388 27748 40462
rect 28140 41188 28196 41198
rect 27916 40292 27972 40302
rect 27972 40236 28084 40292
rect 27916 40198 27972 40236
rect 28028 38612 28084 40236
rect 28140 39730 28196 41132
rect 28252 40178 28308 40190
rect 28252 40126 28254 40178
rect 28306 40126 28308 40178
rect 28252 39956 28308 40126
rect 28252 39890 28308 39900
rect 28140 39678 28142 39730
rect 28194 39678 28196 39730
rect 28140 39666 28196 39678
rect 28252 39618 28308 39630
rect 28252 39566 28254 39618
rect 28306 39566 28308 39618
rect 28252 39508 28308 39566
rect 28252 39442 28308 39452
rect 28028 38556 28308 38612
rect 27692 37716 27748 38332
rect 28140 38388 28196 38398
rect 28140 38162 28196 38332
rect 28140 38110 28142 38162
rect 28194 38110 28196 38162
rect 28140 38098 28196 38110
rect 28252 38052 28308 38556
rect 27692 37650 27748 37660
rect 27804 37826 27860 37838
rect 27804 37774 27806 37826
rect 27858 37774 27860 37826
rect 27692 37266 27748 37278
rect 27692 37214 27694 37266
rect 27746 37214 27748 37266
rect 27692 37044 27748 37214
rect 27692 36978 27748 36988
rect 27804 37156 27860 37774
rect 28252 37716 28308 37996
rect 28364 37828 28420 41468
rect 28476 41188 28532 41198
rect 28476 41094 28532 41132
rect 28588 40852 28644 40862
rect 28588 40404 28644 40796
rect 28700 40740 28756 40750
rect 28700 40626 28756 40684
rect 28700 40574 28702 40626
rect 28754 40574 28756 40626
rect 28700 40562 28756 40574
rect 28588 40348 28756 40404
rect 28588 39956 28644 39966
rect 28476 39844 28532 39854
rect 28476 39750 28532 39788
rect 28588 38834 28644 39900
rect 28588 38782 28590 38834
rect 28642 38782 28644 38834
rect 28588 38770 28644 38782
rect 28700 38610 28756 40348
rect 28700 38558 28702 38610
rect 28754 38558 28756 38610
rect 28700 38546 28756 38558
rect 28476 38276 28532 38286
rect 28476 38050 28532 38220
rect 28476 37998 28478 38050
rect 28530 37998 28532 38050
rect 28476 37986 28532 37998
rect 28364 37772 28532 37828
rect 28252 37660 28420 37716
rect 27356 36764 27524 36820
rect 27132 34862 27134 34914
rect 27186 34862 27188 34914
rect 27132 34692 27188 34862
rect 27132 34626 27188 34636
rect 27356 34804 27412 34814
rect 27356 34356 27412 34748
rect 27132 34354 27412 34356
rect 27132 34302 27358 34354
rect 27410 34302 27412 34354
rect 27132 34300 27412 34302
rect 27020 33906 27076 33918
rect 27020 33854 27022 33906
rect 27074 33854 27076 33906
rect 27020 32562 27076 33854
rect 27132 33234 27188 34300
rect 27356 34290 27412 34300
rect 27132 33182 27134 33234
rect 27186 33182 27188 33234
rect 27132 33170 27188 33182
rect 27020 32510 27022 32562
rect 27074 32510 27076 32562
rect 27020 32498 27076 32510
rect 27468 32452 27524 36764
rect 27804 36370 27860 37100
rect 27916 37156 27972 37166
rect 27916 37154 28084 37156
rect 27916 37102 27918 37154
rect 27970 37102 28084 37154
rect 27916 37100 28084 37102
rect 27916 37090 27972 37100
rect 27916 36596 27972 36606
rect 27916 36502 27972 36540
rect 27804 36318 27806 36370
rect 27858 36318 27860 36370
rect 27804 36148 27860 36318
rect 27804 36082 27860 36092
rect 28028 36482 28084 37100
rect 28028 36430 28030 36482
rect 28082 36430 28084 36482
rect 28028 35252 28084 36430
rect 28252 36484 28308 36494
rect 28252 36390 28308 36428
rect 28364 36482 28420 37660
rect 28364 36430 28366 36482
rect 28418 36430 28420 36482
rect 28364 36418 28420 36430
rect 28140 35588 28196 35598
rect 28140 35494 28196 35532
rect 28476 35252 28532 37772
rect 28588 37268 28644 37278
rect 28588 37174 28644 37212
rect 28028 35186 28084 35196
rect 28252 35196 28532 35252
rect 28140 34914 28196 34926
rect 28140 34862 28142 34914
rect 28194 34862 28196 34914
rect 27580 34804 27636 34814
rect 27580 34710 27636 34748
rect 28140 34804 28196 34862
rect 28140 34738 28196 34748
rect 28252 34468 28308 35196
rect 28476 35028 28532 35038
rect 28476 34934 28532 34972
rect 28364 34914 28420 34926
rect 28364 34862 28366 34914
rect 28418 34862 28420 34914
rect 28364 34580 28420 34862
rect 28588 34916 28644 34926
rect 28588 34822 28644 34860
rect 28364 34524 28644 34580
rect 28252 34412 28420 34468
rect 28252 34242 28308 34254
rect 28252 34190 28254 34242
rect 28306 34190 28308 34242
rect 27692 34132 27748 34142
rect 27692 34130 27972 34132
rect 27692 34078 27694 34130
rect 27746 34078 27972 34130
rect 27692 34076 27972 34078
rect 27692 34066 27748 34076
rect 27804 33460 27860 33470
rect 27804 32676 27860 33404
rect 27916 33012 27972 34076
rect 28140 34020 28196 34030
rect 28140 33926 28196 33964
rect 28028 33908 28084 33918
rect 28028 33814 28084 33852
rect 28252 33684 28308 34190
rect 28140 33628 28308 33684
rect 27916 32956 28084 33012
rect 27916 32676 27972 32686
rect 27804 32620 27916 32676
rect 27916 32582 27972 32620
rect 27468 32396 27972 32452
rect 27692 31556 27748 31566
rect 27244 31220 27300 31230
rect 26908 31164 27244 31220
rect 27244 31154 27300 31164
rect 27692 31218 27748 31500
rect 27692 31166 27694 31218
rect 27746 31166 27748 31218
rect 27692 31154 27748 31166
rect 27356 30996 27412 31006
rect 27244 30940 27356 30996
rect 27020 30882 27076 30894
rect 27020 30830 27022 30882
rect 27074 30830 27076 30882
rect 26796 29426 26852 29438
rect 26796 29374 26798 29426
rect 26850 29374 26852 29426
rect 26796 29204 26852 29374
rect 27020 29316 27076 30830
rect 27244 29764 27300 30940
rect 27356 30902 27412 30940
rect 27804 30884 27860 30894
rect 27580 30882 27860 30884
rect 27580 30830 27806 30882
rect 27858 30830 27860 30882
rect 27580 30828 27860 30830
rect 27356 29988 27412 29998
rect 27580 29988 27636 30828
rect 27804 30818 27860 30828
rect 27356 29986 27636 29988
rect 27356 29934 27358 29986
rect 27410 29934 27636 29986
rect 27356 29932 27636 29934
rect 27692 30436 27748 30446
rect 27356 29922 27412 29932
rect 27244 29698 27300 29708
rect 27356 29316 27412 29326
rect 27020 29260 27356 29316
rect 27356 29250 27412 29260
rect 26796 29138 26852 29148
rect 27468 27972 27524 29932
rect 27580 29764 27636 29774
rect 27580 28082 27636 29708
rect 27580 28030 27582 28082
rect 27634 28030 27636 28082
rect 27580 28018 27636 28030
rect 27468 27906 27524 27916
rect 26684 27794 26740 27804
rect 26796 27858 26852 27870
rect 26796 27806 26798 27858
rect 26850 27806 26852 27858
rect 26012 27186 26516 27188
rect 26012 27134 26014 27186
rect 26066 27134 26516 27186
rect 26012 27132 26516 27134
rect 26012 27122 26068 27132
rect 25900 27022 25902 27074
rect 25954 27022 25956 27074
rect 25900 27010 25956 27022
rect 25676 26964 25732 26974
rect 25564 26962 25732 26964
rect 25564 26910 25678 26962
rect 25730 26910 25732 26962
rect 25564 26908 25732 26910
rect 25676 26898 25732 26908
rect 26348 26852 26404 26862
rect 25340 26796 25620 26852
rect 25228 25788 25508 25844
rect 25228 25506 25284 25518
rect 25228 25454 25230 25506
rect 25282 25454 25284 25506
rect 25228 24948 25284 25454
rect 25116 24892 25284 24948
rect 25452 24948 25508 25788
rect 25116 23828 25172 24892
rect 25452 24882 25508 24892
rect 25116 23762 25172 23772
rect 25228 24722 25284 24734
rect 25228 24670 25230 24722
rect 25282 24670 25284 24722
rect 25228 23378 25284 24670
rect 25564 24388 25620 26796
rect 26236 26516 26292 26526
rect 26236 26422 26292 26460
rect 26348 26514 26404 26796
rect 26348 26462 26350 26514
rect 26402 26462 26404 26514
rect 26348 26450 26404 26462
rect 25788 26402 25844 26414
rect 25788 26350 25790 26402
rect 25842 26350 25844 26402
rect 25788 25732 25844 26350
rect 26124 26402 26180 26414
rect 26124 26350 26126 26402
rect 26178 26350 26180 26402
rect 25900 26290 25956 26302
rect 25900 26238 25902 26290
rect 25954 26238 25956 26290
rect 25900 26068 25956 26238
rect 25900 26002 25956 26012
rect 26124 26292 26180 26350
rect 26124 25956 26180 26236
rect 26124 25890 26180 25900
rect 25788 25676 26180 25732
rect 25676 25618 25732 25630
rect 25676 25566 25678 25618
rect 25730 25566 25732 25618
rect 25676 24836 25732 25566
rect 26012 25506 26068 25518
rect 26012 25454 26014 25506
rect 26066 25454 26068 25506
rect 25676 24770 25732 24780
rect 25900 24948 25956 24958
rect 25900 24834 25956 24892
rect 25900 24782 25902 24834
rect 25954 24782 25956 24834
rect 25788 24722 25844 24734
rect 25788 24670 25790 24722
rect 25842 24670 25844 24722
rect 25676 24612 25732 24622
rect 25676 24518 25732 24556
rect 25788 24388 25844 24670
rect 25564 24332 25844 24388
rect 25900 24500 25956 24782
rect 25228 23326 25230 23378
rect 25282 23326 25284 23378
rect 25228 23156 25284 23326
rect 25228 23090 25284 23100
rect 25452 23828 25508 23838
rect 25564 23828 25620 24332
rect 25900 24276 25956 24444
rect 25676 24220 25956 24276
rect 25676 23938 25732 24220
rect 26012 24162 26068 25454
rect 26124 25284 26180 25676
rect 26460 25730 26516 27132
rect 26572 27122 26628 27132
rect 26684 27634 26740 27646
rect 26684 27582 26686 27634
rect 26738 27582 26740 27634
rect 26684 27074 26740 27582
rect 26684 27022 26686 27074
rect 26738 27022 26740 27074
rect 26684 27010 26740 27022
rect 26796 27076 26852 27806
rect 27580 27860 27636 27870
rect 27580 27300 27636 27804
rect 27692 27858 27748 30380
rect 27804 30100 27860 30110
rect 27804 28530 27860 30044
rect 27804 28478 27806 28530
rect 27858 28478 27860 28530
rect 27804 28466 27860 28478
rect 27916 28420 27972 32396
rect 28028 31890 28084 32956
rect 28140 32788 28196 33628
rect 28252 33460 28308 33470
rect 28252 33366 28308 33404
rect 28252 32788 28308 32798
rect 28140 32732 28252 32788
rect 28252 32694 28308 32732
rect 28364 32116 28420 34412
rect 28588 32788 28644 34524
rect 28812 34244 28868 42028
rect 29036 41970 29092 44044
rect 29148 42980 29204 44380
rect 29260 44434 29316 44494
rect 29260 44382 29262 44434
rect 29314 44382 29316 44434
rect 29260 43204 29316 44382
rect 29372 43540 29428 43550
rect 29372 43446 29428 43484
rect 29260 43148 29428 43204
rect 29260 42980 29316 42990
rect 29148 42978 29316 42980
rect 29148 42926 29262 42978
rect 29314 42926 29316 42978
rect 29148 42924 29316 42926
rect 29260 42914 29316 42924
rect 29036 41918 29038 41970
rect 29090 41918 29092 41970
rect 29036 40964 29092 41918
rect 29372 41412 29428 43148
rect 29484 42754 29540 45388
rect 30044 44994 30100 45006
rect 30044 44942 30046 44994
rect 30098 44942 30100 44994
rect 29708 44546 29764 44558
rect 29708 44494 29710 44546
rect 29762 44494 29764 44546
rect 29708 44434 29764 44494
rect 29708 44382 29710 44434
rect 29762 44382 29764 44434
rect 29708 44370 29764 44382
rect 29596 43762 29652 43774
rect 29596 43710 29598 43762
rect 29650 43710 29652 43762
rect 29596 43540 29652 43710
rect 29820 43764 29876 43774
rect 30044 43764 30100 44942
rect 30156 44996 30212 45006
rect 30156 44434 30212 44940
rect 30156 44382 30158 44434
rect 30210 44382 30212 44434
rect 30156 44100 30212 44382
rect 30156 44034 30212 44044
rect 30268 43876 30324 45500
rect 30380 45444 30436 45950
rect 30940 45780 30996 46956
rect 31276 46900 31332 46910
rect 31276 46002 31332 46844
rect 31388 46674 31444 48188
rect 31836 48132 31892 49196
rect 31612 48076 31892 48132
rect 31500 47460 31556 47470
rect 31500 47366 31556 47404
rect 31612 46786 31668 48076
rect 31948 47572 32004 49644
rect 32060 47684 32116 50764
rect 32284 49252 32340 51996
rect 32508 51716 32564 52110
rect 32620 51940 32676 52892
rect 32732 52274 32788 53676
rect 32844 53506 32900 53676
rect 32844 53454 32846 53506
rect 32898 53454 32900 53506
rect 32844 52612 32900 53454
rect 32844 52546 32900 52556
rect 33180 53508 33236 53518
rect 33292 53508 33348 55356
rect 33404 55186 33460 55918
rect 33404 55134 33406 55186
rect 33458 55134 33460 55186
rect 33404 55122 33460 55134
rect 33740 55188 33796 56702
rect 33852 56642 33908 56654
rect 33852 56590 33854 56642
rect 33906 56590 33908 56642
rect 33852 56082 33908 56590
rect 33852 56030 33854 56082
rect 33906 56030 33908 56082
rect 33852 56018 33908 56030
rect 33964 56642 34020 56654
rect 33964 56590 33966 56642
rect 34018 56590 34020 56642
rect 33964 56420 34020 56590
rect 33740 55122 33796 55132
rect 33964 55188 34020 56364
rect 33964 55122 34020 55132
rect 33852 54404 33908 54414
rect 33852 54310 33908 54348
rect 34076 54180 34132 59052
rect 34300 57650 34356 59276
rect 34300 57598 34302 57650
rect 34354 57598 34356 57650
rect 34300 57586 34356 57598
rect 34524 56644 34580 59724
rect 34636 59714 34692 59724
rect 34748 59332 34804 59342
rect 34748 59238 34804 59276
rect 35084 59218 35140 59230
rect 35084 59166 35086 59218
rect 35138 59166 35140 59218
rect 35084 58660 35140 59166
rect 35532 59108 35588 59118
rect 35532 59014 35588 59052
rect 36092 59106 36148 59118
rect 36092 59054 36094 59106
rect 36146 59054 36148 59106
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35084 58604 35588 58660
rect 35196 58210 35252 58222
rect 35196 58158 35198 58210
rect 35250 58158 35252 58210
rect 35196 57764 35252 58158
rect 35084 57762 35252 57764
rect 35084 57710 35198 57762
rect 35250 57710 35252 57762
rect 35084 57708 35252 57710
rect 34524 56578 34580 56588
rect 34636 57426 34692 57438
rect 34636 57374 34638 57426
rect 34690 57374 34692 57426
rect 34076 54114 34132 54124
rect 34188 56532 34244 56542
rect 33180 53506 33348 53508
rect 33180 53454 33182 53506
rect 33234 53454 33348 53506
rect 33180 53452 33348 53454
rect 32732 52222 32734 52274
rect 32786 52222 32788 52274
rect 32732 52210 32788 52222
rect 32844 52276 32900 52286
rect 32844 52162 32900 52220
rect 32844 52110 32846 52162
rect 32898 52110 32900 52162
rect 32844 52098 32900 52110
rect 33180 52052 33236 53452
rect 34188 53060 34244 56476
rect 34636 56420 34692 57374
rect 35084 56754 35140 57708
rect 35196 57698 35252 57708
rect 35532 57652 35588 58604
rect 36092 58212 36148 59054
rect 43708 58436 43764 58446
rect 36092 58146 36148 58156
rect 36428 58212 36484 58222
rect 36428 58210 36596 58212
rect 36428 58158 36430 58210
rect 36482 58158 36596 58210
rect 36428 58156 36596 58158
rect 36428 58146 36484 58156
rect 36428 57764 36484 57774
rect 36428 57670 36484 57708
rect 35532 57650 35812 57652
rect 35532 57598 35534 57650
rect 35586 57598 35812 57650
rect 35532 57596 35812 57598
rect 35532 57586 35588 57596
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 35084 56702 35086 56754
rect 35138 56702 35140 56754
rect 35084 56690 35140 56702
rect 34636 56194 34692 56364
rect 34636 56142 34638 56194
rect 34690 56142 34692 56194
rect 34636 56130 34692 56142
rect 35420 56084 35476 56094
rect 35420 55990 35476 56028
rect 34636 55970 34692 55982
rect 34636 55918 34638 55970
rect 34690 55918 34692 55970
rect 34636 54404 34692 55918
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35308 55524 35364 55534
rect 35308 55430 35364 55468
rect 35644 55412 35700 55422
rect 35644 55298 35700 55356
rect 35644 55246 35646 55298
rect 35698 55246 35700 55298
rect 35644 55234 35700 55246
rect 35756 54404 35812 57596
rect 36092 57540 36148 57550
rect 36092 57538 36484 57540
rect 36092 57486 36094 57538
rect 36146 57486 36484 57538
rect 36092 57484 36484 57486
rect 36092 57474 36148 57484
rect 36204 56644 36260 56654
rect 36204 56642 36372 56644
rect 36204 56590 36206 56642
rect 36258 56590 36372 56642
rect 36204 56588 36372 56590
rect 36204 56578 36260 56588
rect 36092 56084 36148 56094
rect 35868 55076 35924 55086
rect 35868 54628 35924 55020
rect 35868 54562 35924 54572
rect 35980 54404 36036 54414
rect 35756 54402 36036 54404
rect 35756 54350 35982 54402
rect 36034 54350 36036 54402
rect 35756 54348 36036 54350
rect 34636 54338 34692 54348
rect 35980 54338 36036 54348
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35084 53844 35140 53854
rect 34300 53620 34356 53630
rect 34300 53526 34356 53564
rect 34188 52994 34244 53004
rect 34524 53508 34580 53518
rect 33292 52946 33348 52958
rect 33292 52894 33294 52946
rect 33346 52894 33348 52946
rect 33292 52836 33348 52894
rect 33516 52946 33572 52958
rect 33516 52894 33518 52946
rect 33570 52894 33572 52946
rect 33292 52770 33348 52780
rect 33404 52834 33460 52846
rect 33404 52782 33406 52834
rect 33458 52782 33460 52834
rect 33180 51996 33348 52052
rect 32620 51884 32900 51940
rect 32508 51660 32676 51716
rect 32396 51604 32452 51642
rect 32396 51538 32452 51548
rect 32396 51380 32452 51390
rect 32396 49922 32452 51324
rect 32508 51378 32564 51390
rect 32508 51326 32510 51378
rect 32562 51326 32564 51378
rect 32508 50932 32564 51326
rect 32508 50866 32564 50876
rect 32620 50596 32676 51660
rect 32620 50530 32676 50540
rect 32732 50148 32788 50158
rect 32396 49870 32398 49922
rect 32450 49870 32452 49922
rect 32396 49858 32452 49870
rect 32620 50092 32732 50148
rect 32284 49196 32452 49252
rect 32060 47618 32116 47628
rect 32172 49028 32228 49038
rect 31836 47516 32004 47572
rect 31836 47012 31892 47516
rect 31948 47346 32004 47358
rect 31948 47294 31950 47346
rect 32002 47294 32004 47346
rect 31948 47236 32004 47294
rect 31948 47170 32004 47180
rect 32172 47236 32228 48972
rect 32284 49026 32340 49038
rect 32284 48974 32286 49026
rect 32338 48974 32340 49026
rect 32284 47460 32340 48974
rect 32284 47394 32340 47404
rect 31836 46956 32004 47012
rect 31612 46734 31614 46786
rect 31666 46734 31668 46786
rect 31612 46722 31668 46734
rect 31388 46622 31390 46674
rect 31442 46622 31444 46674
rect 31388 46610 31444 46622
rect 31276 45950 31278 46002
rect 31330 45950 31332 46002
rect 31276 45938 31332 45950
rect 30940 45686 30996 45724
rect 31164 45892 31220 45902
rect 30380 45378 30436 45388
rect 31164 44660 31220 45836
rect 31388 45666 31444 45678
rect 31388 45614 31390 45666
rect 31442 45614 31444 45666
rect 31388 45556 31444 45614
rect 31388 45490 31444 45500
rect 31164 44594 31220 44604
rect 31052 44212 31108 44222
rect 31052 44210 31556 44212
rect 31052 44158 31054 44210
rect 31106 44158 31556 44210
rect 31052 44156 31556 44158
rect 31052 44146 31108 44156
rect 30268 43810 30324 43820
rect 30380 43764 30436 43774
rect 30044 43708 30212 43764
rect 29596 43474 29652 43484
rect 29708 43538 29764 43550
rect 29708 43486 29710 43538
rect 29762 43486 29764 43538
rect 29708 42868 29764 43486
rect 29708 42802 29764 42812
rect 29820 42866 29876 43708
rect 29932 43538 29988 43550
rect 29932 43486 29934 43538
rect 29986 43486 29988 43538
rect 29932 43316 29988 43486
rect 29932 43250 29988 43260
rect 30044 43540 30100 43550
rect 30044 42978 30100 43484
rect 30044 42926 30046 42978
rect 30098 42926 30100 42978
rect 30044 42914 30100 42926
rect 29820 42814 29822 42866
rect 29874 42814 29876 42866
rect 29820 42802 29876 42814
rect 29484 42702 29486 42754
rect 29538 42702 29540 42754
rect 29484 41858 29540 42702
rect 29484 41806 29486 41858
rect 29538 41806 29540 41858
rect 29484 41794 29540 41806
rect 29708 42644 29764 42654
rect 29036 40898 29092 40908
rect 29260 41356 29428 41412
rect 28924 40402 28980 40414
rect 28924 40350 28926 40402
rect 28978 40350 28980 40402
rect 28924 39956 28980 40350
rect 29036 40404 29092 40414
rect 29036 40290 29092 40348
rect 29036 40238 29038 40290
rect 29090 40238 29092 40290
rect 29036 40226 29092 40238
rect 29148 40402 29204 40414
rect 29148 40350 29150 40402
rect 29202 40350 29204 40402
rect 29148 40068 29204 40350
rect 29148 40002 29204 40012
rect 28924 39890 28980 39900
rect 29260 39620 29316 41356
rect 29372 41186 29428 41198
rect 29372 41134 29374 41186
rect 29426 41134 29428 41186
rect 29372 40740 29428 41134
rect 29372 40674 29428 40684
rect 29484 40628 29540 40666
rect 29484 40562 29540 40572
rect 29148 39564 29316 39620
rect 29484 40402 29540 40414
rect 29484 40350 29486 40402
rect 29538 40350 29540 40402
rect 29148 39508 29204 39564
rect 29148 39442 29204 39452
rect 29260 39394 29316 39406
rect 29260 39342 29262 39394
rect 29314 39342 29316 39394
rect 29036 38834 29092 38846
rect 29036 38782 29038 38834
rect 29090 38782 29092 38834
rect 28924 38500 28980 38510
rect 28924 38164 28980 38444
rect 28924 37154 28980 38108
rect 28924 37102 28926 37154
rect 28978 37102 28980 37154
rect 28924 37090 28980 37102
rect 29036 37268 29092 38782
rect 29260 38834 29316 39342
rect 29484 38948 29540 40350
rect 29596 39620 29652 39630
rect 29596 39526 29652 39564
rect 29484 38882 29540 38892
rect 29260 38782 29262 38834
rect 29314 38782 29316 38834
rect 29260 38668 29316 38782
rect 29260 38612 29428 38668
rect 29148 37940 29204 37950
rect 29148 37846 29204 37884
rect 29036 35364 29092 37212
rect 29148 37716 29204 37726
rect 29148 36370 29204 37660
rect 29372 37266 29428 38612
rect 29372 37214 29374 37266
rect 29426 37214 29428 37266
rect 29372 37202 29428 37214
rect 29484 37938 29540 37950
rect 29484 37886 29486 37938
rect 29538 37886 29540 37938
rect 29148 36318 29150 36370
rect 29202 36318 29204 36370
rect 29148 35922 29204 36318
rect 29148 35870 29150 35922
rect 29202 35870 29204 35922
rect 29148 35858 29204 35870
rect 29372 36484 29428 36494
rect 29484 36484 29540 37886
rect 29372 36482 29540 36484
rect 29372 36430 29374 36482
rect 29426 36430 29540 36482
rect 29372 36428 29540 36430
rect 29372 35588 29428 36428
rect 29372 35522 29428 35532
rect 29036 35308 29540 35364
rect 28700 34188 28868 34244
rect 29148 34802 29204 34814
rect 29148 34750 29150 34802
rect 29202 34750 29204 34802
rect 28700 33012 28756 34188
rect 29148 34132 29204 34750
rect 29260 34690 29316 34702
rect 29260 34638 29262 34690
rect 29314 34638 29316 34690
rect 29260 34356 29316 34638
rect 29372 34692 29428 34702
rect 29372 34598 29428 34636
rect 29260 34290 29316 34300
rect 28812 34076 29204 34132
rect 28812 34018 28868 34076
rect 28812 33966 28814 34018
rect 28866 33966 28868 34018
rect 28812 33236 28868 33966
rect 29260 33908 29316 33918
rect 29484 33908 29540 35308
rect 29596 35028 29652 35038
rect 29596 34130 29652 34972
rect 29596 34078 29598 34130
rect 29650 34078 29652 34130
rect 29596 34066 29652 34078
rect 29260 33906 29540 33908
rect 29260 33854 29262 33906
rect 29314 33854 29540 33906
rect 29260 33852 29540 33854
rect 29260 33842 29316 33852
rect 29372 33460 29428 33470
rect 29260 33404 29372 33460
rect 29260 33346 29316 33404
rect 29372 33394 29428 33404
rect 29260 33294 29262 33346
rect 29314 33294 29316 33346
rect 29260 33282 29316 33294
rect 28812 33170 28868 33180
rect 28700 32956 29092 33012
rect 28812 32788 28868 32798
rect 28588 32732 28812 32788
rect 28812 32694 28868 32732
rect 28028 31838 28030 31890
rect 28082 31838 28084 31890
rect 28028 31826 28084 31838
rect 28252 32060 28420 32116
rect 28476 32676 28532 32686
rect 28252 31444 28308 32060
rect 28364 31892 28420 31902
rect 28364 31798 28420 31836
rect 28476 31778 28532 32620
rect 28924 32564 28980 32574
rect 28924 32470 28980 32508
rect 28476 31726 28478 31778
rect 28530 31726 28532 31778
rect 28476 31714 28532 31726
rect 28700 31892 28756 31902
rect 28252 31388 28420 31444
rect 28252 31220 28308 31230
rect 28028 28420 28084 28430
rect 27916 28418 28084 28420
rect 27916 28366 28030 28418
rect 28082 28366 28084 28418
rect 27916 28364 28084 28366
rect 28028 28354 28084 28364
rect 27692 27806 27694 27858
rect 27746 27806 27748 27858
rect 27692 27794 27748 27806
rect 27692 27300 27748 27310
rect 27580 27298 27748 27300
rect 27580 27246 27694 27298
rect 27746 27246 27748 27298
rect 27580 27244 27748 27246
rect 26796 27010 26852 27020
rect 26908 27188 26964 27198
rect 26684 26852 26740 26862
rect 26908 26852 26964 27132
rect 27356 26852 27412 26862
rect 26684 26292 26740 26796
rect 26796 26796 26964 26852
rect 27132 26850 27412 26852
rect 27132 26798 27358 26850
rect 27410 26798 27412 26850
rect 27132 26796 27412 26798
rect 26796 26514 26852 26796
rect 26796 26462 26798 26514
rect 26850 26462 26852 26514
rect 26796 26450 26852 26462
rect 26684 26236 26852 26292
rect 26460 25678 26462 25730
rect 26514 25678 26516 25730
rect 26460 25666 26516 25678
rect 26236 25508 26292 25518
rect 26236 25414 26292 25452
rect 26124 25228 26292 25284
rect 26012 24110 26014 24162
rect 26066 24110 26068 24162
rect 26012 24098 26068 24110
rect 25676 23886 25678 23938
rect 25730 23886 25732 23938
rect 25676 23874 25732 23886
rect 26124 23938 26180 23950
rect 26124 23886 26126 23938
rect 26178 23886 26180 23938
rect 25452 23826 25620 23828
rect 25452 23774 25454 23826
rect 25506 23774 25620 23826
rect 25452 23772 25620 23774
rect 25788 23828 25844 23838
rect 25900 23828 25956 23838
rect 25844 23826 25956 23828
rect 25844 23774 25902 23826
rect 25954 23774 25956 23826
rect 25844 23772 25956 23774
rect 25452 22596 25508 23772
rect 25788 23154 25844 23772
rect 25900 23762 25956 23772
rect 26124 23604 26180 23886
rect 26236 23828 26292 25228
rect 26684 25172 26740 25182
rect 26348 24164 26404 24174
rect 26348 24070 26404 24108
rect 26236 23762 26292 23772
rect 26124 23538 26180 23548
rect 25788 23102 25790 23154
rect 25842 23102 25844 23154
rect 25788 23090 25844 23102
rect 26460 23268 26516 23278
rect 25676 22596 25732 22606
rect 25452 22594 25732 22596
rect 25452 22542 25678 22594
rect 25730 22542 25732 22594
rect 25452 22540 25732 22542
rect 25676 22530 25732 22540
rect 25228 22484 25284 22494
rect 25228 22370 25284 22428
rect 25228 22318 25230 22370
rect 25282 22318 25284 22370
rect 25228 22306 25284 22318
rect 26460 22372 26516 23212
rect 26460 22278 26516 22316
rect 25004 22082 25060 22092
rect 24668 21812 24724 21822
rect 24556 21588 24612 21598
rect 24556 21494 24612 21532
rect 24220 21474 24388 21476
rect 24220 21422 24222 21474
rect 24274 21422 24388 21474
rect 24220 21420 24388 21422
rect 24220 21410 24276 21420
rect 24108 20132 24164 21196
rect 24668 20914 24724 21756
rect 25116 21700 25172 21710
rect 25004 21252 25060 21262
rect 24668 20862 24670 20914
rect 24722 20862 24724 20914
rect 24668 20850 24724 20862
rect 24892 21028 24948 21038
rect 24892 20802 24948 20972
rect 24892 20750 24894 20802
rect 24946 20750 24948 20802
rect 24892 20738 24948 20750
rect 25004 20468 25060 21196
rect 25116 20690 25172 21644
rect 26460 21700 26516 21710
rect 26460 21606 26516 21644
rect 25340 21588 25396 21598
rect 25340 21494 25396 21532
rect 25116 20638 25118 20690
rect 25170 20638 25172 20690
rect 25116 20626 25172 20638
rect 25228 21140 25284 21150
rect 25228 20690 25284 21084
rect 25228 20638 25230 20690
rect 25282 20638 25284 20690
rect 24892 20412 25060 20468
rect 24332 20244 24388 20254
rect 24388 20188 24500 20244
rect 24332 20178 24388 20188
rect 24108 20066 24164 20076
rect 24108 19908 24164 19918
rect 24108 18674 24164 19852
rect 24220 19906 24276 19918
rect 24220 19854 24222 19906
rect 24274 19854 24276 19906
rect 24220 19796 24276 19854
rect 24220 19730 24276 19740
rect 24220 19234 24276 19246
rect 24220 19182 24222 19234
rect 24274 19182 24276 19234
rect 24220 19012 24276 19182
rect 24220 18946 24276 18956
rect 24332 19124 24388 19134
rect 24108 18622 24110 18674
rect 24162 18622 24164 18674
rect 24108 18610 24164 18622
rect 24332 18674 24388 19068
rect 24332 18622 24334 18674
rect 24386 18622 24388 18674
rect 24332 18610 24388 18622
rect 24220 18452 24276 18462
rect 23996 18450 24276 18452
rect 23996 18398 24222 18450
rect 24274 18398 24276 18450
rect 23996 18396 24276 18398
rect 24220 18386 24276 18396
rect 23772 18274 23828 18284
rect 23884 18338 23940 18350
rect 23884 18286 23886 18338
rect 23938 18286 23940 18338
rect 23884 18116 23940 18286
rect 23884 18050 23940 18060
rect 23772 17220 23828 17230
rect 23660 17164 23772 17220
rect 23772 17154 23828 17164
rect 24332 17108 24388 17118
rect 24444 17108 24500 20188
rect 24668 20132 24724 20142
rect 24724 20076 24836 20132
rect 24668 20066 24724 20076
rect 24780 20018 24836 20076
rect 24780 19966 24782 20018
rect 24834 19966 24836 20018
rect 24780 19954 24836 19966
rect 24892 19572 24948 20412
rect 25228 19684 25284 20638
rect 25676 20802 25732 20814
rect 25676 20750 25678 20802
rect 25730 20750 25732 20802
rect 25452 20020 25508 20030
rect 25452 19926 25508 19964
rect 25228 19618 25284 19628
rect 25564 19906 25620 19918
rect 25564 19854 25566 19906
rect 25618 19854 25620 19906
rect 25564 19572 25620 19854
rect 24892 19516 25060 19572
rect 24556 19122 24612 19134
rect 24556 19070 24558 19122
rect 24610 19070 24612 19122
rect 24556 18900 24612 19070
rect 24668 19124 24724 19134
rect 24668 19030 24724 19068
rect 24556 18834 24612 18844
rect 24780 19010 24836 19022
rect 24780 18958 24782 19010
rect 24834 18958 24836 19010
rect 24668 18676 24724 18686
rect 24668 18450 24724 18620
rect 24668 18398 24670 18450
rect 24722 18398 24724 18450
rect 24668 18386 24724 18398
rect 24668 17444 24724 17454
rect 24332 17106 24500 17108
rect 24332 17054 24334 17106
rect 24386 17054 24500 17106
rect 24332 17052 24500 17054
rect 24556 17108 24612 17118
rect 24332 17042 24388 17052
rect 24556 17014 24612 17052
rect 23884 16996 23940 17006
rect 23884 16902 23940 16940
rect 24668 16994 24724 17388
rect 24668 16942 24670 16994
rect 24722 16942 24724 16994
rect 24668 16930 24724 16942
rect 23548 16884 23604 16894
rect 23548 16790 23604 16828
rect 24108 16884 24164 16894
rect 24108 16882 24276 16884
rect 24108 16830 24110 16882
rect 24162 16830 24276 16882
rect 24108 16828 24276 16830
rect 24108 16818 24164 16828
rect 23996 16772 24052 16782
rect 23996 16678 24052 16716
rect 23436 15988 23492 15998
rect 23436 15894 23492 15932
rect 24108 15876 24164 15886
rect 24108 15782 24164 15820
rect 22652 14756 22708 15148
rect 22428 14702 22430 14754
rect 22482 14702 22484 14754
rect 22428 14690 22484 14702
rect 22540 14754 22708 14756
rect 22540 14702 22654 14754
rect 22706 14702 22708 14754
rect 22540 14700 22708 14702
rect 22316 13860 22372 13870
rect 22540 13860 22596 14700
rect 22652 14690 22708 14700
rect 22764 15092 23044 15148
rect 23212 15204 23268 15242
rect 23212 15138 23268 15148
rect 22316 13858 22596 13860
rect 22316 13806 22318 13858
rect 22370 13806 22596 13858
rect 22316 13804 22596 13806
rect 22316 13794 22372 13804
rect 22204 13458 22260 13468
rect 21868 12798 21870 12850
rect 21922 12798 21924 12850
rect 21868 11620 21924 12798
rect 21980 13412 22036 13422
rect 21980 12292 22036 13356
rect 22652 13300 22708 13310
rect 22652 12962 22708 13244
rect 22652 12910 22654 12962
rect 22706 12910 22708 12962
rect 22652 12898 22708 12910
rect 22092 12740 22148 12778
rect 22092 12674 22148 12684
rect 22764 12628 22820 15092
rect 22876 14420 22932 14430
rect 22876 13746 22932 14364
rect 22876 13694 22878 13746
rect 22930 13694 22932 13746
rect 22876 13188 22932 13694
rect 23100 13858 23156 13870
rect 23100 13806 23102 13858
rect 23154 13806 23156 13858
rect 23100 13524 23156 13806
rect 23324 13524 23380 15596
rect 23436 15316 23492 15326
rect 23436 15222 23492 15260
rect 23772 15202 23828 15214
rect 23772 15150 23774 15202
rect 23826 15150 23828 15202
rect 23772 14532 23828 15150
rect 24108 15204 24164 15242
rect 24108 15138 24164 15148
rect 24220 15148 24276 16828
rect 24556 16100 24612 16110
rect 24332 15876 24388 15886
rect 24332 15316 24388 15820
rect 24388 15260 24500 15316
rect 24332 15250 24388 15260
rect 24220 15092 24388 15148
rect 23772 14466 23828 14476
rect 23996 14420 24052 14430
rect 23996 13970 24052 14364
rect 23996 13918 23998 13970
rect 24050 13918 24052 13970
rect 23996 13906 24052 13918
rect 24332 13970 24388 15092
rect 24444 14980 24500 15260
rect 24444 14914 24500 14924
rect 24332 13918 24334 13970
rect 24386 13918 24388 13970
rect 24332 13906 24388 13918
rect 24444 14418 24500 14430
rect 24444 14366 24446 14418
rect 24498 14366 24500 14418
rect 23660 13636 23716 13646
rect 23660 13542 23716 13580
rect 23324 13468 23604 13524
rect 23100 13458 23156 13468
rect 22876 13122 22932 13132
rect 22988 13300 23044 13310
rect 22876 12964 22932 12974
rect 22876 12870 22932 12908
rect 22764 12572 22932 12628
rect 21980 12226 22036 12236
rect 22092 12516 22148 12526
rect 22092 12290 22148 12460
rect 22428 12404 22484 12414
rect 22092 12238 22094 12290
rect 22146 12238 22148 12290
rect 22092 12226 22148 12238
rect 22316 12292 22372 12302
rect 22316 12198 22372 12236
rect 22316 11956 22372 11966
rect 22428 11956 22484 12348
rect 22764 12404 22820 12414
rect 22764 12178 22820 12348
rect 22764 12126 22766 12178
rect 22818 12126 22820 12178
rect 22764 12114 22820 12126
rect 22372 11900 22484 11956
rect 22540 12066 22596 12078
rect 22540 12014 22542 12066
rect 22594 12014 22596 12066
rect 21868 11564 22260 11620
rect 21868 11396 21924 11406
rect 21868 11302 21924 11340
rect 21868 10836 21924 10846
rect 21868 10742 21924 10780
rect 22092 10836 22148 10846
rect 22092 10742 22148 10780
rect 21980 10500 22036 10510
rect 21980 10498 22148 10500
rect 21980 10446 21982 10498
rect 22034 10446 22148 10498
rect 21980 10444 22148 10446
rect 21980 10434 22036 10444
rect 21756 9998 21758 10050
rect 21810 9998 21812 10050
rect 21420 9716 21476 9726
rect 21420 9622 21476 9660
rect 21644 9716 21700 9726
rect 20972 9212 21252 9268
rect 20188 8530 20244 8540
rect 20300 8540 20580 8596
rect 20748 8932 20804 8942
rect 20076 8372 20244 8428
rect 20076 8260 20132 8270
rect 19964 8258 20132 8260
rect 19964 8206 20078 8258
rect 20130 8206 20132 8258
rect 19964 8204 20132 8206
rect 20076 8194 20132 8204
rect 19180 7980 19460 8036
rect 19068 5842 19124 5852
rect 18844 5234 19012 5236
rect 18844 5182 18846 5234
rect 18898 5182 19012 5234
rect 18844 5180 19012 5182
rect 19404 5234 19460 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20076 7586 20132 7598
rect 20076 7534 20078 7586
rect 20130 7534 20132 7586
rect 20076 6804 20132 7534
rect 20188 7364 20244 8372
rect 20300 8370 20356 8540
rect 20636 8484 20692 8494
rect 20524 8428 20636 8484
rect 20300 8318 20302 8370
rect 20354 8318 20356 8370
rect 20300 8306 20356 8318
rect 20412 8372 20468 8382
rect 20412 8258 20468 8316
rect 20412 8206 20414 8258
rect 20466 8206 20468 8258
rect 20412 8194 20468 8206
rect 20412 7700 20468 7710
rect 20524 7700 20580 8428
rect 20636 8418 20692 8428
rect 20412 7698 20580 7700
rect 20412 7646 20414 7698
rect 20466 7646 20580 7698
rect 20412 7644 20580 7646
rect 20412 7634 20468 7644
rect 20300 7588 20356 7598
rect 20300 7494 20356 7532
rect 20300 7364 20356 7374
rect 20188 7362 20356 7364
rect 20188 7310 20302 7362
rect 20354 7310 20356 7362
rect 20188 7308 20356 7310
rect 20300 7298 20356 7308
rect 20076 6738 20132 6748
rect 20188 7140 20244 7150
rect 20188 6690 20244 7084
rect 20524 6802 20580 7644
rect 20636 7700 20692 7710
rect 20748 7700 20804 8876
rect 20636 7698 20804 7700
rect 20636 7646 20638 7698
rect 20690 7646 20804 7698
rect 20636 7644 20804 7646
rect 20636 7634 20692 7644
rect 20524 6750 20526 6802
rect 20578 6750 20580 6802
rect 20524 6738 20580 6750
rect 20860 6804 20916 9212
rect 20972 9042 21028 9054
rect 20972 8990 20974 9042
rect 21026 8990 21028 9042
rect 20972 7588 21028 8990
rect 21084 9044 21140 9054
rect 21084 8950 21140 8988
rect 21196 7700 21252 9212
rect 21644 9042 21700 9660
rect 21644 8990 21646 9042
rect 21698 8990 21700 9042
rect 21084 7588 21140 7598
rect 20972 7532 21084 7588
rect 21196 7588 21252 7644
rect 21420 8596 21476 8606
rect 21420 8258 21476 8540
rect 21420 8206 21422 8258
rect 21474 8206 21476 8258
rect 21196 7532 21364 7588
rect 21084 7250 21140 7532
rect 21084 7198 21086 7250
rect 21138 7198 21140 7250
rect 21084 7186 21140 7198
rect 20860 6738 20916 6748
rect 20188 6638 20190 6690
rect 20242 6638 20244 6690
rect 20188 6626 20244 6638
rect 19628 6580 19684 6590
rect 19628 6486 19684 6524
rect 20412 6580 20468 6590
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20412 6130 20468 6524
rect 21308 6578 21364 7532
rect 21308 6526 21310 6578
rect 21362 6526 21364 6578
rect 21308 6514 21364 6526
rect 20412 6078 20414 6130
rect 20466 6078 20468 6130
rect 20412 6066 20468 6078
rect 20860 6356 20916 6366
rect 19852 5908 19908 5918
rect 19852 5814 19908 5852
rect 20860 5908 20916 6300
rect 21084 6356 21140 6366
rect 21420 6356 21476 8206
rect 21644 8484 21700 8990
rect 21756 8932 21812 9998
rect 21980 9716 22036 9726
rect 21980 9622 22036 9660
rect 21756 8838 21812 8876
rect 21644 7474 21700 8428
rect 22092 8370 22148 10444
rect 22092 8318 22094 8370
rect 22146 8318 22148 8370
rect 22092 8306 22148 8318
rect 21644 7422 21646 7474
rect 21698 7422 21700 7474
rect 21644 7410 21700 7422
rect 22204 7028 22260 11564
rect 22316 11396 22372 11900
rect 22316 11394 22484 11396
rect 22316 11342 22318 11394
rect 22370 11342 22484 11394
rect 22316 11340 22484 11342
rect 22316 11330 22372 11340
rect 22092 6972 22260 7028
rect 22316 10722 22372 10734
rect 22316 10670 22318 10722
rect 22370 10670 22372 10722
rect 21644 6692 21700 6702
rect 21644 6598 21700 6636
rect 21980 6580 22036 6590
rect 21980 6486 22036 6524
rect 20972 6132 21028 6142
rect 20972 6038 21028 6076
rect 20300 5348 20356 5358
rect 19404 5182 19406 5234
rect 19458 5182 19460 5234
rect 18844 5170 18900 5180
rect 19404 5170 19460 5182
rect 19964 5236 20020 5246
rect 19964 5142 20020 5180
rect 20300 5234 20356 5292
rect 20300 5182 20302 5234
rect 20354 5182 20356 5234
rect 20300 5170 20356 5182
rect 20860 5234 20916 5852
rect 20860 5182 20862 5234
rect 20914 5182 20916 5234
rect 20860 5170 20916 5182
rect 21084 5348 21140 6300
rect 15484 5124 15540 5134
rect 15148 5068 15484 5124
rect 15484 5030 15540 5068
rect 16940 5124 16996 5134
rect 16940 4340 16996 5068
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 21084 4562 21140 5292
rect 21084 4510 21086 4562
rect 21138 4510 21140 4562
rect 21084 4498 21140 4510
rect 21308 6300 21476 6356
rect 22092 6356 22148 6972
rect 22204 6804 22260 6814
rect 22204 6710 22260 6748
rect 22316 6580 22372 10670
rect 22428 8596 22484 11340
rect 22540 10612 22596 12014
rect 22540 10546 22596 10556
rect 22652 11732 22708 11742
rect 22652 11060 22708 11676
rect 22540 9714 22596 9726
rect 22540 9662 22542 9714
rect 22594 9662 22596 9714
rect 22540 8932 22596 9662
rect 22540 8866 22596 8876
rect 22428 8530 22484 8540
rect 22428 7476 22484 7486
rect 22428 7382 22484 7420
rect 22316 6514 22372 6524
rect 21308 4564 21364 6300
rect 22092 6290 22148 6300
rect 22204 6468 22260 6478
rect 21868 6244 21924 6254
rect 21420 6132 21476 6142
rect 21420 6038 21476 6076
rect 21644 6132 21700 6142
rect 21644 5236 21700 6076
rect 21532 4900 21588 4910
rect 21644 4900 21700 5180
rect 21868 5234 21924 6188
rect 21980 6132 22036 6142
rect 21980 6038 22036 6076
rect 22204 6132 22260 6412
rect 22652 6132 22708 11004
rect 22764 11396 22820 11406
rect 22764 9604 22820 11340
rect 22876 10836 22932 12572
rect 22988 12290 23044 13244
rect 23212 13188 23268 13198
rect 23436 13188 23492 13198
rect 23212 13186 23380 13188
rect 23212 13134 23214 13186
rect 23266 13134 23380 13186
rect 23212 13132 23380 13134
rect 23212 13122 23268 13132
rect 23212 12964 23268 12974
rect 22988 12238 22990 12290
rect 23042 12238 23044 12290
rect 22988 12226 23044 12238
rect 23100 12738 23156 12750
rect 23100 12686 23102 12738
rect 23154 12686 23156 12738
rect 23100 11508 23156 12686
rect 23212 12290 23268 12908
rect 23212 12238 23214 12290
rect 23266 12238 23268 12290
rect 23212 12226 23268 12238
rect 23324 12180 23380 13132
rect 23436 12962 23492 13132
rect 23436 12910 23438 12962
rect 23490 12910 23492 12962
rect 23436 12628 23492 12910
rect 23436 12562 23492 12572
rect 23436 12180 23492 12190
rect 23324 12124 23436 12180
rect 23436 12086 23492 12124
rect 23548 11956 23604 13468
rect 23996 13412 24052 13422
rect 23996 12962 24052 13356
rect 24332 13188 24388 13198
rect 24332 12964 24388 13132
rect 23996 12910 23998 12962
rect 24050 12910 24052 12962
rect 23996 12898 24052 12910
rect 24108 12962 24388 12964
rect 24108 12910 24334 12962
rect 24386 12910 24388 12962
rect 24108 12908 24388 12910
rect 23772 12852 23828 12862
rect 23100 11442 23156 11452
rect 23212 11900 23604 11956
rect 23660 12850 23828 12852
rect 23660 12798 23774 12850
rect 23826 12798 23828 12850
rect 23660 12796 23828 12798
rect 23660 12178 23716 12796
rect 23772 12786 23828 12796
rect 23660 12126 23662 12178
rect 23714 12126 23716 12178
rect 23660 11956 23716 12126
rect 22988 11284 23044 11294
rect 22988 11282 23156 11284
rect 22988 11230 22990 11282
rect 23042 11230 23156 11282
rect 22988 11228 23156 11230
rect 22988 11218 23044 11228
rect 22876 10770 22932 10780
rect 22988 10386 23044 10398
rect 22988 10334 22990 10386
rect 23042 10334 23044 10386
rect 22876 10052 22932 10062
rect 22876 9958 22932 9996
rect 22988 9828 23044 10334
rect 23100 10386 23156 11228
rect 23212 10724 23268 11900
rect 23660 11890 23716 11900
rect 23772 12402 23828 12414
rect 24108 12404 24164 12908
rect 24332 12898 24388 12908
rect 23772 12350 23774 12402
rect 23826 12350 23828 12402
rect 23548 11732 23604 11742
rect 23548 11172 23604 11676
rect 23548 11106 23604 11116
rect 23660 11620 23716 11630
rect 23212 10722 23380 10724
rect 23212 10670 23214 10722
rect 23266 10670 23380 10722
rect 23212 10668 23380 10670
rect 23212 10658 23268 10668
rect 23100 10334 23102 10386
rect 23154 10334 23156 10386
rect 23100 10322 23156 10334
rect 23212 9828 23268 9838
rect 22988 9772 23156 9828
rect 22988 9604 23044 9614
rect 22764 9602 23044 9604
rect 22764 9550 22990 9602
rect 23042 9550 23044 9602
rect 22764 9548 23044 9550
rect 22988 9538 23044 9548
rect 22988 8372 23044 8382
rect 22876 7588 22932 7598
rect 22876 7474 22932 7532
rect 22876 7422 22878 7474
rect 22930 7422 22932 7474
rect 22876 7410 22932 7422
rect 22988 6692 23044 8316
rect 23100 6914 23156 9772
rect 23212 9734 23268 9772
rect 23324 9492 23380 10668
rect 23548 10612 23604 10622
rect 23548 10518 23604 10556
rect 23548 10276 23604 10286
rect 23436 9716 23492 9726
rect 23436 9622 23492 9660
rect 23324 9426 23380 9436
rect 23212 9042 23268 9054
rect 23212 8990 23214 9042
rect 23266 8990 23268 9042
rect 23212 7364 23268 8990
rect 23436 9042 23492 9054
rect 23436 8990 23438 9042
rect 23490 8990 23492 9042
rect 23324 8932 23380 8942
rect 23324 8838 23380 8876
rect 23436 7588 23492 8990
rect 23436 7522 23492 7532
rect 23212 7362 23380 7364
rect 23212 7310 23214 7362
rect 23266 7310 23380 7362
rect 23212 7308 23380 7310
rect 23212 7298 23268 7308
rect 23100 6862 23102 6914
rect 23154 6862 23156 6914
rect 23100 6850 23156 6862
rect 22988 6580 23044 6636
rect 23100 6580 23156 6590
rect 22988 6578 23156 6580
rect 22988 6526 23102 6578
rect 23154 6526 23156 6578
rect 22988 6524 23156 6526
rect 23100 6514 23156 6524
rect 23212 6578 23268 6590
rect 23212 6526 23214 6578
rect 23266 6526 23268 6578
rect 23212 6468 23268 6526
rect 23212 6402 23268 6412
rect 22988 6132 23044 6142
rect 22652 6130 23044 6132
rect 22652 6078 22990 6130
rect 23042 6078 23044 6130
rect 22652 6076 23044 6078
rect 22204 6066 22260 6076
rect 22988 6066 23044 6076
rect 22428 5908 22484 5946
rect 22428 5842 22484 5852
rect 21868 5182 21870 5234
rect 21922 5182 21924 5234
rect 21868 5170 21924 5182
rect 22428 5682 22484 5694
rect 22428 5630 22430 5682
rect 22482 5630 22484 5682
rect 22428 5234 22484 5630
rect 23324 5684 23380 7308
rect 23548 6692 23604 10220
rect 23660 9380 23716 11564
rect 23772 10610 23828 12350
rect 23772 10558 23774 10610
rect 23826 10558 23828 10610
rect 23772 10546 23828 10558
rect 23884 12348 24108 12404
rect 23660 9324 23828 9380
rect 23660 9154 23716 9166
rect 23660 9102 23662 9154
rect 23714 9102 23716 9154
rect 23660 7476 23716 9102
rect 23660 7410 23716 7420
rect 23772 6692 23828 9324
rect 23548 6626 23604 6636
rect 23660 6636 23828 6692
rect 23548 6468 23604 6478
rect 23324 5590 23380 5628
rect 23436 6356 23492 6366
rect 23436 6130 23492 6300
rect 23436 6078 23438 6130
rect 23490 6078 23492 6130
rect 22428 5182 22430 5234
rect 22482 5182 22484 5234
rect 22428 5170 22484 5182
rect 22988 5236 23044 5246
rect 22988 5142 23044 5180
rect 23212 5012 23268 5022
rect 21532 4898 21700 4900
rect 21532 4846 21534 4898
rect 21586 4846 21700 4898
rect 21532 4844 21700 4846
rect 21980 4900 22036 4910
rect 21532 4834 21588 4844
rect 21532 4564 21588 4574
rect 21980 4564 22036 4844
rect 21308 4562 22036 4564
rect 21308 4510 21534 4562
rect 21586 4510 21982 4562
rect 22034 4510 22036 4562
rect 21308 4508 22036 4510
rect 21532 4498 21588 4508
rect 21980 4498 22036 4508
rect 22764 4788 22820 4798
rect 22764 4562 22820 4732
rect 22764 4510 22766 4562
rect 22818 4510 22820 4562
rect 22764 4498 22820 4510
rect 23212 4562 23268 4956
rect 23212 4510 23214 4562
rect 23266 4510 23268 4562
rect 23212 4498 23268 4510
rect 16940 4274 16996 4284
rect 23436 3388 23492 6078
rect 23548 3666 23604 6412
rect 23660 6132 23716 6636
rect 23772 6466 23828 6478
rect 23772 6414 23774 6466
rect 23826 6414 23828 6466
rect 23772 6356 23828 6414
rect 23772 6290 23828 6300
rect 23660 6066 23716 6076
rect 23660 5908 23716 5918
rect 23660 5234 23716 5852
rect 23660 5182 23662 5234
rect 23714 5182 23716 5234
rect 23660 4788 23716 5182
rect 23660 4722 23716 4732
rect 23772 5572 23828 5582
rect 23660 4564 23716 4574
rect 23772 4564 23828 5516
rect 23884 5236 23940 12348
rect 24108 12338 24164 12348
rect 24220 12738 24276 12750
rect 24220 12686 24222 12738
rect 24274 12686 24276 12738
rect 24108 12178 24164 12190
rect 24108 12126 24110 12178
rect 24162 12126 24164 12178
rect 23996 12068 24052 12078
rect 23996 11620 24052 12012
rect 23996 11554 24052 11564
rect 23996 11284 24052 11294
rect 23996 10836 24052 11228
rect 24108 10948 24164 12126
rect 24220 11732 24276 12686
rect 24332 12404 24388 12414
rect 24332 12290 24388 12348
rect 24332 12238 24334 12290
rect 24386 12238 24388 12290
rect 24332 12226 24388 12238
rect 24444 11844 24500 14366
rect 24556 13970 24612 16044
rect 24668 15876 24724 15886
rect 24668 15538 24724 15820
rect 24668 15486 24670 15538
rect 24722 15486 24724 15538
rect 24668 15474 24724 15486
rect 24556 13918 24558 13970
rect 24610 13918 24612 13970
rect 24556 13906 24612 13918
rect 24668 13860 24724 13870
rect 24780 13860 24836 18958
rect 24892 19012 24948 19022
rect 24892 18918 24948 18956
rect 24892 18452 24948 18462
rect 24892 17778 24948 18396
rect 24892 17726 24894 17778
rect 24946 17726 24948 17778
rect 24892 17556 24948 17726
rect 24892 17490 24948 17500
rect 25004 17108 25060 19516
rect 25564 19506 25620 19516
rect 25564 19234 25620 19246
rect 25564 19182 25566 19234
rect 25618 19182 25620 19234
rect 25564 18228 25620 19182
rect 25004 17042 25060 17052
rect 25116 17444 25172 17454
rect 25564 17444 25620 18172
rect 25676 17892 25732 20750
rect 26124 20690 26180 20702
rect 26124 20638 26126 20690
rect 26178 20638 26180 20690
rect 25900 20578 25956 20590
rect 25900 20526 25902 20578
rect 25954 20526 25956 20578
rect 25900 20130 25956 20526
rect 25900 20078 25902 20130
rect 25954 20078 25956 20130
rect 25900 18676 25956 20078
rect 26124 20132 26180 20638
rect 26572 20690 26628 20702
rect 26572 20638 26574 20690
rect 26626 20638 26628 20690
rect 26124 20076 26404 20132
rect 26348 20018 26404 20076
rect 26348 19966 26350 20018
rect 26402 19966 26404 20018
rect 26236 19908 26292 19918
rect 26236 19124 26292 19852
rect 26348 19796 26404 19966
rect 26348 19236 26404 19740
rect 26572 19460 26628 20638
rect 26684 20132 26740 25116
rect 26796 24722 26852 26236
rect 26796 24670 26798 24722
rect 26850 24670 26852 24722
rect 26796 24658 26852 24670
rect 27020 25508 27076 25518
rect 27132 25508 27188 26796
rect 27356 26786 27412 26796
rect 27580 26852 27636 27244
rect 27692 27234 27748 27244
rect 27804 26964 27860 26974
rect 27580 26786 27636 26796
rect 27692 26908 27804 26964
rect 27020 25506 27188 25508
rect 27020 25454 27022 25506
rect 27074 25454 27188 25506
rect 27020 25452 27188 25454
rect 27580 25730 27636 25742
rect 27580 25678 27582 25730
rect 27634 25678 27636 25730
rect 26684 20066 26740 20076
rect 26796 24052 26852 24062
rect 26684 19460 26740 19470
rect 26572 19404 26684 19460
rect 26684 19366 26740 19404
rect 26348 19170 26404 19180
rect 26684 19234 26740 19246
rect 26684 19182 26686 19234
rect 26738 19182 26740 19234
rect 26236 19058 26292 19068
rect 26684 18900 26740 19182
rect 26684 18834 26740 18844
rect 25900 18610 25956 18620
rect 25788 18564 25844 18574
rect 25788 18470 25844 18508
rect 26796 18116 26852 23996
rect 27020 23938 27076 25452
rect 27132 24500 27188 24510
rect 27132 24406 27188 24444
rect 27580 24164 27636 25678
rect 27020 23886 27022 23938
rect 27074 23886 27076 23938
rect 27020 23874 27076 23886
rect 27132 24162 27636 24164
rect 27132 24110 27582 24162
rect 27634 24110 27636 24162
rect 27132 24108 27636 24110
rect 27132 21026 27188 24108
rect 27580 24098 27636 24108
rect 27356 23828 27412 23838
rect 27356 22370 27412 23772
rect 27692 23548 27748 26908
rect 27804 26898 27860 26908
rect 27916 26962 27972 26974
rect 27916 26910 27918 26962
rect 27970 26910 27972 26962
rect 27916 26292 27972 26910
rect 27916 24722 27972 26236
rect 28028 26402 28084 26414
rect 28028 26350 28030 26402
rect 28082 26350 28084 26402
rect 28028 25060 28084 26350
rect 28140 25394 28196 25406
rect 28140 25342 28142 25394
rect 28194 25342 28196 25394
rect 28140 25284 28196 25342
rect 28140 25218 28196 25228
rect 28140 25060 28196 25070
rect 28028 25004 28140 25060
rect 28140 24994 28196 25004
rect 27916 24670 27918 24722
rect 27970 24670 27972 24722
rect 27916 24658 27972 24670
rect 28252 23940 28308 31164
rect 28364 29652 28420 31388
rect 28700 30882 28756 31836
rect 28924 30996 28980 31006
rect 29036 30996 29092 32956
rect 29372 32564 29428 32574
rect 29372 32470 29428 32508
rect 29708 31892 29764 42588
rect 30156 42530 30212 43708
rect 30380 43670 30436 43708
rect 31500 43762 31556 44156
rect 31500 43710 31502 43762
rect 31554 43710 31556 43762
rect 31500 43698 31556 43710
rect 30604 43652 30660 43662
rect 30268 43538 30324 43550
rect 30268 43486 30270 43538
rect 30322 43486 30324 43538
rect 30268 42980 30324 43486
rect 30604 43540 30660 43596
rect 31612 43650 31668 43662
rect 31612 43598 31614 43650
rect 31666 43598 31668 43650
rect 31052 43540 31108 43550
rect 30604 43538 30772 43540
rect 30604 43486 30606 43538
rect 30658 43486 30772 43538
rect 30604 43484 30772 43486
rect 30604 43474 30660 43484
rect 30604 43092 30660 43102
rect 30492 42980 30548 42990
rect 30268 42924 30492 42980
rect 30492 42754 30548 42924
rect 30492 42702 30494 42754
rect 30546 42702 30548 42754
rect 30492 42690 30548 42702
rect 30156 42478 30158 42530
rect 30210 42478 30212 42530
rect 30156 42466 30212 42478
rect 30604 42308 30660 43036
rect 30380 42252 30660 42308
rect 30716 42754 30772 43484
rect 31052 43446 31108 43484
rect 31500 43428 31556 43438
rect 30716 42702 30718 42754
rect 30770 42702 30772 42754
rect 30716 42532 30772 42702
rect 30828 43314 30884 43326
rect 30828 43262 30830 43314
rect 30882 43262 30884 43314
rect 30828 42756 30884 43262
rect 31164 43316 31220 43326
rect 31388 43316 31444 43326
rect 30940 42756 30996 42766
rect 30828 42754 30996 42756
rect 30828 42702 30942 42754
rect 30994 42702 30996 42754
rect 30828 42700 30996 42702
rect 30044 41970 30100 41982
rect 30044 41918 30046 41970
rect 30098 41918 30100 41970
rect 29820 41188 29876 41198
rect 29876 41132 29988 41188
rect 29820 41094 29876 41132
rect 29820 40178 29876 40190
rect 29820 40126 29822 40178
rect 29874 40126 29876 40178
rect 29820 39844 29876 40126
rect 29820 38050 29876 39788
rect 29932 39506 29988 41132
rect 30044 40852 30100 41918
rect 30268 41970 30324 41982
rect 30268 41918 30270 41970
rect 30322 41918 30324 41970
rect 30156 41860 30212 41870
rect 30156 41766 30212 41804
rect 30044 40786 30100 40796
rect 30268 40740 30324 41918
rect 30156 40684 30324 40740
rect 29932 39454 29934 39506
rect 29986 39454 29988 39506
rect 29932 39442 29988 39454
rect 30044 40404 30100 40414
rect 30156 40404 30212 40684
rect 30268 40516 30324 40526
rect 30380 40516 30436 42252
rect 30716 42196 30772 42476
rect 30492 42140 30772 42196
rect 30492 41188 30548 42140
rect 30604 41970 30660 41982
rect 30604 41918 30606 41970
rect 30658 41918 30660 41970
rect 30604 41412 30660 41918
rect 30940 41748 30996 42700
rect 31164 42754 31220 43260
rect 31164 42702 31166 42754
rect 31218 42702 31220 42754
rect 31164 42644 31220 42702
rect 31164 42578 31220 42588
rect 31276 43314 31444 43316
rect 31276 43262 31390 43314
rect 31442 43262 31444 43314
rect 31276 43260 31444 43262
rect 31052 42532 31108 42542
rect 31052 41970 31108 42476
rect 31276 42530 31332 43260
rect 31388 43250 31444 43260
rect 31276 42478 31278 42530
rect 31330 42478 31332 42530
rect 31276 42466 31332 42478
rect 31388 42980 31444 42990
rect 31276 42084 31332 42094
rect 31388 42084 31444 42924
rect 31500 42754 31556 43372
rect 31612 42868 31668 43598
rect 31724 42868 31780 42878
rect 31612 42866 31780 42868
rect 31612 42814 31726 42866
rect 31778 42814 31780 42866
rect 31612 42812 31780 42814
rect 31724 42802 31780 42812
rect 31836 42868 31892 42878
rect 31500 42702 31502 42754
rect 31554 42702 31556 42754
rect 31500 42690 31556 42702
rect 31836 42754 31892 42812
rect 31836 42702 31838 42754
rect 31890 42702 31892 42754
rect 31836 42084 31892 42702
rect 31948 42532 32004 46956
rect 32172 46786 32228 47180
rect 32172 46734 32174 46786
rect 32226 46734 32228 46786
rect 32172 46722 32228 46734
rect 32396 45892 32452 49196
rect 32620 49138 32676 50092
rect 32732 50082 32788 50092
rect 32844 49924 32900 51884
rect 33068 49924 33124 49934
rect 32844 49922 33124 49924
rect 32844 49870 33070 49922
rect 33122 49870 33124 49922
rect 32844 49868 33124 49870
rect 33068 49858 33124 49868
rect 33180 49924 33236 49934
rect 33180 49830 33236 49868
rect 33292 49812 33348 51996
rect 33404 51380 33460 52782
rect 33516 52388 33572 52894
rect 33516 52322 33572 52332
rect 33964 52946 34020 52958
rect 33964 52894 33966 52946
rect 34018 52894 34020 52946
rect 33404 51314 33460 51324
rect 33516 52164 33572 52174
rect 33516 51378 33572 52108
rect 33516 51326 33518 51378
rect 33570 51326 33572 51378
rect 33516 51314 33572 51326
rect 33628 52052 33684 52062
rect 33628 51154 33684 51996
rect 33964 51492 34020 52894
rect 34524 52946 34580 53452
rect 34524 52894 34526 52946
rect 34578 52894 34580 52946
rect 34524 52882 34580 52894
rect 35084 52948 35140 53788
rect 36092 53730 36148 56028
rect 36204 56082 36260 56094
rect 36204 56030 36206 56082
rect 36258 56030 36260 56082
rect 36204 54740 36260 56030
rect 36316 55300 36372 56588
rect 36316 55234 36372 55244
rect 36316 55076 36372 55086
rect 36428 55076 36484 57484
rect 36316 55074 36484 55076
rect 36316 55022 36318 55074
rect 36370 55022 36484 55074
rect 36316 55020 36484 55022
rect 36316 55010 36372 55020
rect 36428 54964 36484 55020
rect 36428 54898 36484 54908
rect 36316 54740 36372 54750
rect 36204 54738 36372 54740
rect 36204 54686 36318 54738
rect 36370 54686 36372 54738
rect 36204 54684 36372 54686
rect 36316 54674 36372 54684
rect 36540 54740 36596 58156
rect 37100 58210 37156 58222
rect 37100 58158 37102 58210
rect 37154 58158 37156 58210
rect 37100 57988 37156 58158
rect 37100 57922 37156 57932
rect 40012 58212 40068 58222
rect 39564 57876 39620 57886
rect 36876 57540 36932 57550
rect 37324 57540 37380 57550
rect 36876 57538 37044 57540
rect 36876 57486 36878 57538
rect 36930 57486 37044 57538
rect 36876 57484 37044 57486
rect 36876 57474 36932 57484
rect 36988 55860 37044 57484
rect 37324 57446 37380 57484
rect 37772 57538 37828 57550
rect 37772 57486 37774 57538
rect 37826 57486 37828 57538
rect 37212 57090 37268 57102
rect 37212 57038 37214 57090
rect 37266 57038 37268 57090
rect 37100 56756 37156 56766
rect 37100 56662 37156 56700
rect 37100 56084 37156 56094
rect 37100 55990 37156 56028
rect 36988 55804 37156 55860
rect 36876 55524 36932 55534
rect 36540 54674 36596 54684
rect 36652 55300 36708 55310
rect 36652 54516 36708 55244
rect 36092 53678 36094 53730
rect 36146 53678 36148 53730
rect 36092 53666 36148 53678
rect 36204 54514 36708 54516
rect 36204 54462 36654 54514
rect 36706 54462 36708 54514
rect 36204 54460 36708 54462
rect 36204 53730 36260 54460
rect 36652 54450 36708 54460
rect 36764 54964 36820 54974
rect 36204 53678 36206 53730
rect 36258 53678 36260 53730
rect 36204 53666 36260 53678
rect 35420 53508 35476 53518
rect 35420 53414 35476 53452
rect 36204 53508 36260 53518
rect 35084 52854 35140 52892
rect 34748 52836 34804 52846
rect 34748 52834 35028 52836
rect 34748 52782 34750 52834
rect 34802 52782 35028 52834
rect 34748 52780 35028 52782
rect 34748 52770 34804 52780
rect 33964 51398 34020 51436
rect 34188 52722 34244 52734
rect 34188 52670 34190 52722
rect 34242 52670 34244 52722
rect 33628 51102 33630 51154
rect 33682 51102 33684 51154
rect 33628 51090 33684 51102
rect 33516 50708 33572 50718
rect 33516 50614 33572 50652
rect 33404 50594 33460 50606
rect 33404 50542 33406 50594
rect 33458 50542 33460 50594
rect 33404 50034 33460 50542
rect 33404 49982 33406 50034
rect 33458 49982 33460 50034
rect 33404 49970 33460 49982
rect 33740 49922 33796 49934
rect 33740 49870 33742 49922
rect 33794 49870 33796 49922
rect 33292 49756 33460 49812
rect 32620 49086 32622 49138
rect 32674 49086 32676 49138
rect 32620 49074 32676 49086
rect 33180 48692 33236 48702
rect 33068 48356 33124 48366
rect 33068 48242 33124 48300
rect 33180 48354 33236 48636
rect 33180 48302 33182 48354
rect 33234 48302 33236 48354
rect 33180 48290 33236 48302
rect 33068 48190 33070 48242
rect 33122 48190 33124 48242
rect 32620 48130 32676 48142
rect 32620 48078 32622 48130
rect 32674 48078 32676 48130
rect 32620 47348 32676 48078
rect 33068 47796 33124 48190
rect 33068 47730 33124 47740
rect 33068 47572 33124 47582
rect 33068 47348 33124 47516
rect 32620 47346 33124 47348
rect 32620 47294 33070 47346
rect 33122 47294 33124 47346
rect 32620 47292 33124 47294
rect 32508 46788 32564 46798
rect 32508 46694 32564 46732
rect 32284 45836 32452 45892
rect 32172 45780 32228 45790
rect 32172 44994 32228 45724
rect 32172 44942 32174 44994
rect 32226 44942 32228 44994
rect 32172 44930 32228 44942
rect 32172 43650 32228 43662
rect 32172 43598 32174 43650
rect 32226 43598 32228 43650
rect 32060 43540 32116 43550
rect 32060 42868 32116 43484
rect 32060 42754 32116 42812
rect 32060 42702 32062 42754
rect 32114 42702 32116 42754
rect 32060 42690 32116 42702
rect 32172 42644 32228 43598
rect 32172 42578 32228 42588
rect 31948 42466 32004 42476
rect 31276 42082 31444 42084
rect 31276 42030 31278 42082
rect 31330 42030 31444 42082
rect 31276 42028 31444 42030
rect 31724 42028 31892 42084
rect 31276 42018 31332 42028
rect 31052 41918 31054 41970
rect 31106 41918 31108 41970
rect 31052 41906 31108 41918
rect 30940 41692 31108 41748
rect 30604 41356 30996 41412
rect 30940 41298 30996 41356
rect 30940 41246 30942 41298
rect 30994 41246 30996 41298
rect 30604 41188 30660 41198
rect 30492 41186 30660 41188
rect 30492 41134 30606 41186
rect 30658 41134 30660 41186
rect 30492 41132 30660 41134
rect 30604 41122 30660 41132
rect 30268 40514 30436 40516
rect 30268 40462 30270 40514
rect 30322 40462 30436 40514
rect 30268 40460 30436 40462
rect 30268 40450 30324 40460
rect 30044 40402 30212 40404
rect 30044 40350 30046 40402
rect 30098 40350 30212 40402
rect 30044 40348 30212 40350
rect 30044 40292 30100 40348
rect 29932 38388 29988 38398
rect 30044 38388 30100 40236
rect 30380 39508 30436 40460
rect 30828 40964 30884 40974
rect 30492 40404 30548 40414
rect 30492 40310 30548 40348
rect 29988 38332 30100 38388
rect 30268 39506 30436 39508
rect 30268 39454 30382 39506
rect 30434 39454 30436 39506
rect 30268 39452 30436 39454
rect 29932 38322 29988 38332
rect 29820 37998 29822 38050
rect 29874 37998 29876 38050
rect 29820 37986 29876 37998
rect 29932 38052 29988 38062
rect 30156 38052 30212 38062
rect 29988 38050 30212 38052
rect 29988 37998 30158 38050
rect 30210 37998 30212 38050
rect 29988 37996 30212 37998
rect 29932 37986 29988 37996
rect 30156 37986 30212 37996
rect 30268 38052 30324 39452
rect 30380 39442 30436 39452
rect 30716 39060 30772 39070
rect 30268 37986 30324 37996
rect 30380 38948 30436 38958
rect 30380 36482 30436 38892
rect 30716 38946 30772 39004
rect 30716 38894 30718 38946
rect 30770 38894 30772 38946
rect 30716 38882 30772 38894
rect 30828 38668 30884 40908
rect 30940 39842 30996 41246
rect 31052 41074 31108 41692
rect 31724 41636 31780 42028
rect 32284 41972 32340 45836
rect 32396 45668 32452 45678
rect 32396 45574 32452 45612
rect 32844 45556 32900 45566
rect 32956 45556 33012 47292
rect 33068 47282 33124 47292
rect 33292 47458 33348 47470
rect 33292 47406 33294 47458
rect 33346 47406 33348 47458
rect 33292 45892 33348 47406
rect 33404 47068 33460 49756
rect 33740 49476 33796 49870
rect 34188 49810 34244 52670
rect 34636 52724 34692 52734
rect 34188 49758 34190 49810
rect 34242 49758 34244 49810
rect 34188 49746 34244 49758
rect 34300 52276 34356 52286
rect 33740 49410 33796 49420
rect 34188 49476 34244 49486
rect 33628 48916 33684 48926
rect 33628 47682 33684 48860
rect 33740 48692 33796 48702
rect 33740 48354 33796 48636
rect 33740 48302 33742 48354
rect 33794 48302 33796 48354
rect 33740 48290 33796 48302
rect 33852 48132 33908 48142
rect 33852 48038 33908 48076
rect 33628 47630 33630 47682
rect 33682 47630 33684 47682
rect 33628 47618 33684 47630
rect 34076 47346 34132 47358
rect 34076 47294 34078 47346
rect 34130 47294 34132 47346
rect 33404 47012 33572 47068
rect 33292 45826 33348 45836
rect 33404 46786 33460 46798
rect 33404 46734 33406 46786
rect 33458 46734 33460 46786
rect 33068 45780 33124 45790
rect 33124 45724 33236 45780
rect 33068 45714 33124 45724
rect 32900 45500 33012 45556
rect 32844 45490 32900 45500
rect 32844 45108 32900 45118
rect 32844 44546 32900 45052
rect 32844 44494 32846 44546
rect 32898 44494 32900 44546
rect 32844 44482 32900 44494
rect 33068 43652 33124 43662
rect 33068 43558 33124 43596
rect 31948 41916 32340 41972
rect 32396 43538 32452 43550
rect 32396 43486 32398 43538
rect 32450 43486 32452 43538
rect 32396 41972 32452 43486
rect 32508 42868 32564 42878
rect 32508 42774 32564 42812
rect 33180 42754 33236 45724
rect 33404 45332 33460 46734
rect 33516 46116 33572 47012
rect 34076 47012 34132 47294
rect 34076 46946 34132 46956
rect 33852 46786 33908 46798
rect 33852 46734 33854 46786
rect 33906 46734 33908 46786
rect 33516 46050 33572 46060
rect 33628 46674 33684 46686
rect 33628 46622 33630 46674
rect 33682 46622 33684 46674
rect 33404 45266 33460 45276
rect 33516 45666 33572 45678
rect 33516 45614 33518 45666
rect 33570 45614 33572 45666
rect 33404 45108 33460 45118
rect 33516 45108 33572 45614
rect 33404 45106 33572 45108
rect 33404 45054 33406 45106
rect 33458 45054 33572 45106
rect 33404 45052 33572 45054
rect 33404 44996 33460 45052
rect 33292 44882 33348 44894
rect 33292 44830 33294 44882
rect 33346 44830 33348 44882
rect 33292 44324 33348 44830
rect 33292 44258 33348 44268
rect 33404 43762 33460 44940
rect 33628 44324 33684 46622
rect 33852 46676 33908 46734
rect 33852 46620 34132 46676
rect 33740 46562 33796 46574
rect 33740 46510 33742 46562
rect 33794 46510 33796 46562
rect 33740 46116 33796 46510
rect 33740 46050 33796 46060
rect 33964 45780 34020 45790
rect 33964 45686 34020 45724
rect 33740 45108 33796 45118
rect 34076 45108 34132 46620
rect 34188 46674 34244 49420
rect 34300 49026 34356 52220
rect 34636 52052 34692 52668
rect 34972 52388 35028 52780
rect 35868 52834 35924 52846
rect 35868 52782 35870 52834
rect 35922 52782 35924 52834
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 34972 52332 35364 52388
rect 34860 52164 34916 52202
rect 34860 52098 34916 52108
rect 35084 52162 35140 52174
rect 35084 52110 35086 52162
rect 35138 52110 35140 52162
rect 34300 48974 34302 49026
rect 34354 48974 34356 49026
rect 34300 48242 34356 48974
rect 34300 48190 34302 48242
rect 34354 48190 34356 48242
rect 34300 47684 34356 48190
rect 34412 52050 34692 52052
rect 34412 51998 34638 52050
rect 34690 51998 34692 52050
rect 34412 51996 34692 51998
rect 34412 48914 34468 51996
rect 34636 51986 34692 51996
rect 34748 52052 34804 52062
rect 34636 51604 34692 51614
rect 34524 51044 34580 51054
rect 34524 50818 34580 50988
rect 34524 50766 34526 50818
rect 34578 50766 34580 50818
rect 34524 50754 34580 50766
rect 34412 48862 34414 48914
rect 34466 48862 34468 48914
rect 34412 48132 34468 48862
rect 34412 48066 34468 48076
rect 34524 50596 34580 50606
rect 34300 47618 34356 47628
rect 34300 47460 34356 47470
rect 34300 47366 34356 47404
rect 34188 46622 34190 46674
rect 34242 46622 34244 46674
rect 34188 46610 34244 46622
rect 34300 45668 34356 45678
rect 34300 45574 34356 45612
rect 34076 45052 34468 45108
rect 33740 45014 33796 45052
rect 33964 44996 34020 45006
rect 33964 44902 34020 44940
rect 34300 44884 34356 44894
rect 33628 44258 33684 44268
rect 34188 44882 34356 44884
rect 34188 44830 34302 44882
rect 34354 44830 34356 44882
rect 34188 44828 34356 44830
rect 33404 43710 33406 43762
rect 33458 43710 33460 43762
rect 33404 43698 33460 43710
rect 34076 43650 34132 43662
rect 34076 43598 34078 43650
rect 34130 43598 34132 43650
rect 34076 43092 34132 43598
rect 34188 43538 34244 44828
rect 34300 44818 34356 44828
rect 34412 44436 34468 45052
rect 34412 44342 34468 44380
rect 34300 44324 34356 44334
rect 34300 43764 34356 44268
rect 34412 43764 34468 43774
rect 34300 43708 34412 43764
rect 34412 43698 34468 43708
rect 34188 43486 34190 43538
rect 34242 43486 34244 43538
rect 34188 43474 34244 43486
rect 34300 43540 34356 43550
rect 34076 43026 34132 43036
rect 34300 42756 34356 43484
rect 33180 42702 33182 42754
rect 33234 42702 33236 42754
rect 33180 42690 33236 42702
rect 34076 42754 34356 42756
rect 34076 42702 34302 42754
rect 34354 42702 34356 42754
rect 34076 42700 34356 42702
rect 32620 42644 32676 42654
rect 32620 42550 32676 42588
rect 33404 42532 33460 42542
rect 33404 42530 33572 42532
rect 33404 42478 33406 42530
rect 33458 42478 33572 42530
rect 33404 42476 33572 42478
rect 33404 42466 33460 42476
rect 31836 41860 31892 41870
rect 31836 41766 31892 41804
rect 31724 41580 31892 41636
rect 31052 41022 31054 41074
rect 31106 41022 31108 41074
rect 31052 41010 31108 41022
rect 31388 41186 31444 41198
rect 31388 41134 31390 41186
rect 31442 41134 31444 41186
rect 31164 40852 31220 40862
rect 31388 40852 31444 41134
rect 31220 40796 31444 40852
rect 31724 41074 31780 41086
rect 31724 41022 31726 41074
rect 31778 41022 31780 41074
rect 31164 40290 31220 40796
rect 31500 40740 31556 40750
rect 31164 40238 31166 40290
rect 31218 40238 31220 40290
rect 31164 40226 31220 40238
rect 31276 40402 31332 40414
rect 31276 40350 31278 40402
rect 31330 40350 31332 40402
rect 31276 40292 31332 40350
rect 31276 40226 31332 40236
rect 31164 40068 31220 40078
rect 30940 39790 30942 39842
rect 30994 39790 30996 39842
rect 30940 39778 30996 39790
rect 31052 39956 31108 39966
rect 31052 39618 31108 39900
rect 31164 39732 31220 40012
rect 31164 39730 31332 39732
rect 31164 39678 31166 39730
rect 31218 39678 31332 39730
rect 31164 39676 31332 39678
rect 31164 39666 31220 39676
rect 31052 39566 31054 39618
rect 31106 39566 31108 39618
rect 31052 38836 31108 39566
rect 31052 38834 31220 38836
rect 31052 38782 31054 38834
rect 31106 38782 31220 38834
rect 31052 38780 31220 38782
rect 31052 38770 31108 38780
rect 30380 36430 30382 36482
rect 30434 36430 30436 36482
rect 30380 36418 30436 36430
rect 30604 38612 30660 38622
rect 30604 37044 30660 38556
rect 30380 36148 30436 36158
rect 29820 35252 29876 35262
rect 29820 34242 29876 35196
rect 29820 34190 29822 34242
rect 29874 34190 29876 34242
rect 29820 34178 29876 34190
rect 29932 34916 29988 34926
rect 30156 34916 30212 34926
rect 29988 34914 30212 34916
rect 29988 34862 30158 34914
rect 30210 34862 30212 34914
rect 29988 34860 30212 34862
rect 29932 33908 29988 34860
rect 30156 34850 30212 34860
rect 30268 34802 30324 34814
rect 30268 34750 30270 34802
rect 30322 34750 30324 34802
rect 29932 33852 30100 33908
rect 30044 33458 30100 33852
rect 30044 33406 30046 33458
rect 30098 33406 30100 33458
rect 29932 33348 29988 33358
rect 29932 32788 29988 33292
rect 29932 32722 29988 32732
rect 29708 31826 29764 31836
rect 29708 31666 29764 31678
rect 29708 31614 29710 31666
rect 29762 31614 29764 31666
rect 28924 30994 29092 30996
rect 28924 30942 28926 30994
rect 28978 30942 29092 30994
rect 28924 30940 29092 30942
rect 28924 30930 28980 30940
rect 28700 30830 28702 30882
rect 28754 30830 28756 30882
rect 28700 30660 28756 30830
rect 28756 30604 28980 30660
rect 28700 30594 28756 30604
rect 28476 30436 28532 30446
rect 28476 30210 28532 30380
rect 28476 30158 28478 30210
rect 28530 30158 28532 30210
rect 28476 30146 28532 30158
rect 28364 29596 28868 29652
rect 28812 29538 28868 29596
rect 28812 29486 28814 29538
rect 28866 29486 28868 29538
rect 28700 29426 28756 29438
rect 28700 29374 28702 29426
rect 28754 29374 28756 29426
rect 28700 29316 28756 29374
rect 28700 29250 28756 29260
rect 28476 29204 28532 29214
rect 28364 28756 28420 28766
rect 28364 28530 28420 28700
rect 28476 28642 28532 29148
rect 28476 28590 28478 28642
rect 28530 28590 28532 28642
rect 28476 28578 28532 28590
rect 28364 28478 28366 28530
rect 28418 28478 28420 28530
rect 28364 28466 28420 28478
rect 28812 28420 28868 29486
rect 28812 28354 28868 28364
rect 28588 27972 28644 27982
rect 28588 27878 28644 27916
rect 28476 26962 28532 26974
rect 28476 26910 28478 26962
rect 28530 26910 28532 26962
rect 28364 26404 28420 26414
rect 28364 24836 28420 26348
rect 28476 25732 28532 26910
rect 28924 26908 28980 30604
rect 29036 30212 29092 30940
rect 29148 31554 29204 31566
rect 29148 31502 29150 31554
rect 29202 31502 29204 31554
rect 29148 30436 29204 31502
rect 29596 30996 29652 31006
rect 29596 30902 29652 30940
rect 29148 30370 29204 30380
rect 29484 30770 29540 30782
rect 29484 30718 29486 30770
rect 29538 30718 29540 30770
rect 29036 30156 29204 30212
rect 29036 29428 29092 29438
rect 29036 29334 29092 29372
rect 29148 28756 29204 30156
rect 29484 28868 29540 30718
rect 29708 30210 29764 31614
rect 30044 31220 30100 33406
rect 30156 33348 30212 33358
rect 30268 33348 30324 34750
rect 30380 34242 30436 36092
rect 30604 35922 30660 36988
rect 30604 35870 30606 35922
rect 30658 35870 30660 35922
rect 30604 35858 30660 35870
rect 30716 38612 30884 38668
rect 30380 34190 30382 34242
rect 30434 34190 30436 34242
rect 30380 34178 30436 34190
rect 30380 33572 30436 33582
rect 30380 33570 30660 33572
rect 30380 33518 30382 33570
rect 30434 33518 30660 33570
rect 30380 33516 30660 33518
rect 30380 33506 30436 33516
rect 30212 33292 30324 33348
rect 30156 33282 30212 33292
rect 30492 33012 30548 33022
rect 30492 32786 30548 32956
rect 30492 32734 30494 32786
rect 30546 32734 30548 32786
rect 30492 32722 30548 32734
rect 30380 32564 30436 32574
rect 30268 31556 30324 31566
rect 30268 31462 30324 31500
rect 30044 31154 30100 31164
rect 30380 31218 30436 32508
rect 30380 31166 30382 31218
rect 30434 31166 30436 31218
rect 30380 31154 30436 31166
rect 29708 30158 29710 30210
rect 29762 30158 29764 30210
rect 29708 29092 29764 30158
rect 29708 29026 29764 29036
rect 29932 31106 29988 31118
rect 29932 31054 29934 31106
rect 29986 31054 29988 31106
rect 29932 30098 29988 31054
rect 29932 30046 29934 30098
rect 29986 30046 29988 30098
rect 29148 28662 29204 28700
rect 29372 28812 29540 28868
rect 29932 28868 29988 30046
rect 30492 30324 30548 30334
rect 30492 29426 30548 30268
rect 30492 29374 30494 29426
rect 30546 29374 30548 29426
rect 30492 29362 30548 29374
rect 30156 29316 30212 29326
rect 30156 29222 30212 29260
rect 28476 25666 28532 25676
rect 28700 26852 28980 26908
rect 29148 26962 29204 26974
rect 29148 26910 29150 26962
rect 29202 26910 29204 26962
rect 28700 25618 28756 26852
rect 29036 26628 29092 26638
rect 29036 26290 29092 26572
rect 29148 26516 29204 26910
rect 29148 26450 29204 26460
rect 29260 26962 29316 26974
rect 29260 26910 29262 26962
rect 29314 26910 29316 26962
rect 29036 26238 29038 26290
rect 29090 26238 29092 26290
rect 29036 26226 29092 26238
rect 28700 25566 28702 25618
rect 28754 25566 28756 25618
rect 28700 25554 28756 25566
rect 29148 26068 29204 26078
rect 28364 24780 28532 24836
rect 28476 24276 28532 24780
rect 29148 24834 29204 26012
rect 29148 24782 29150 24834
rect 29202 24782 29204 24834
rect 29148 24770 29204 24782
rect 28364 23940 28420 23950
rect 28140 23938 28420 23940
rect 28140 23886 28366 23938
rect 28418 23886 28420 23938
rect 28140 23884 28420 23886
rect 27916 23828 27972 23838
rect 27916 23734 27972 23772
rect 27692 23492 27860 23548
rect 27804 23380 27860 23492
rect 27692 23324 27860 23380
rect 27580 23268 27636 23278
rect 27580 23154 27636 23212
rect 27580 23102 27582 23154
rect 27634 23102 27636 23154
rect 27580 23090 27636 23102
rect 27356 22318 27358 22370
rect 27410 22318 27412 22370
rect 27356 21364 27412 22318
rect 27356 21298 27412 21308
rect 27468 22484 27524 22494
rect 27132 20974 27134 21026
rect 27186 20974 27188 21026
rect 27132 20962 27188 20974
rect 27468 21026 27524 22428
rect 27468 20974 27470 21026
rect 27522 20974 27524 21026
rect 27468 20962 27524 20974
rect 27692 20804 27748 23324
rect 27916 23268 27972 23278
rect 27804 23156 27860 23166
rect 27804 23062 27860 23100
rect 27468 20748 27748 20804
rect 27916 20802 27972 23212
rect 28028 22932 28084 22942
rect 28028 22258 28084 22876
rect 28028 22206 28030 22258
rect 28082 22206 28084 22258
rect 28028 22194 28084 22206
rect 28028 21698 28084 21710
rect 28028 21646 28030 21698
rect 28082 21646 28084 21698
rect 28028 21252 28084 21646
rect 28028 21186 28084 21196
rect 27916 20750 27918 20802
rect 27970 20750 27972 20802
rect 27244 20132 27300 20142
rect 27132 20020 27188 20030
rect 27020 19234 27076 19246
rect 27020 19182 27022 19234
rect 27074 19182 27076 19234
rect 27020 19012 27076 19182
rect 27132 19234 27188 19964
rect 27132 19182 27134 19234
rect 27186 19182 27188 19234
rect 27132 19170 27188 19182
rect 27244 19906 27300 20076
rect 27244 19854 27246 19906
rect 27298 19854 27300 19906
rect 27020 18946 27076 18956
rect 27244 18564 27300 19854
rect 27244 18498 27300 18508
rect 27356 19794 27412 19806
rect 27356 19742 27358 19794
rect 27410 19742 27412 19794
rect 27020 18340 27076 18350
rect 27020 18246 27076 18284
rect 26796 18050 26852 18060
rect 25676 17798 25732 17836
rect 26460 18004 26516 18014
rect 25116 15652 25172 17388
rect 25452 17388 25620 17444
rect 25900 17780 25956 17790
rect 25452 16994 25508 17388
rect 25452 16942 25454 16994
rect 25506 16942 25508 16994
rect 25452 16930 25508 16942
rect 25788 16996 25844 17006
rect 25788 16902 25844 16940
rect 25564 16882 25620 16894
rect 25564 16830 25566 16882
rect 25618 16830 25620 16882
rect 25564 16772 25620 16830
rect 25564 16706 25620 16716
rect 25676 16770 25732 16782
rect 25676 16718 25678 16770
rect 25730 16718 25732 16770
rect 25564 16324 25620 16334
rect 25228 15876 25284 15886
rect 25228 15874 25508 15876
rect 25228 15822 25230 15874
rect 25282 15822 25508 15874
rect 25228 15820 25508 15822
rect 25228 15810 25284 15820
rect 25116 15540 25172 15596
rect 25228 15540 25284 15550
rect 25116 15538 25284 15540
rect 25116 15486 25230 15538
rect 25282 15486 25284 15538
rect 25116 15484 25284 15486
rect 25228 15474 25284 15484
rect 24668 13858 24836 13860
rect 24668 13806 24670 13858
rect 24722 13806 24836 13858
rect 24668 13804 24836 13806
rect 24892 15204 24948 15214
rect 24668 13794 24724 13804
rect 24668 13524 24724 13534
rect 24668 12850 24724 13468
rect 24668 12798 24670 12850
rect 24722 12798 24724 12850
rect 24668 12786 24724 12798
rect 24780 12178 24836 12190
rect 24780 12126 24782 12178
rect 24834 12126 24836 12178
rect 24556 12068 24612 12078
rect 24556 11974 24612 12012
rect 24444 11788 24724 11844
rect 24220 11676 24612 11732
rect 24332 11508 24388 11518
rect 24108 10882 24164 10892
rect 24220 11172 24276 11182
rect 23996 9938 24052 10780
rect 23996 9886 23998 9938
rect 24050 9886 24052 9938
rect 23996 7812 24052 9886
rect 24220 10276 24276 11116
rect 24332 10722 24388 11452
rect 24556 10834 24612 11676
rect 24556 10782 24558 10834
rect 24610 10782 24612 10834
rect 24556 10770 24612 10782
rect 24332 10670 24334 10722
rect 24386 10670 24388 10722
rect 24332 10658 24388 10670
rect 24668 10498 24724 11788
rect 24780 10724 24836 12126
rect 24780 10658 24836 10668
rect 24668 10446 24670 10498
rect 24722 10446 24724 10498
rect 24668 10434 24724 10446
rect 24220 9826 24276 10220
rect 24892 9828 24948 15148
rect 25228 14532 25284 14542
rect 25228 14438 25284 14476
rect 25340 14306 25396 14318
rect 25340 14254 25342 14306
rect 25394 14254 25396 14306
rect 25340 14196 25396 14254
rect 25340 14130 25396 14140
rect 25452 14308 25508 15820
rect 25564 15538 25620 16268
rect 25676 16100 25732 16718
rect 25676 16034 25732 16044
rect 25564 15486 25566 15538
rect 25618 15486 25620 15538
rect 25564 15474 25620 15486
rect 25452 13970 25508 14252
rect 25452 13918 25454 13970
rect 25506 13918 25508 13970
rect 25452 13906 25508 13918
rect 25788 14532 25844 14542
rect 25564 13748 25620 13758
rect 25452 13524 25508 13534
rect 25004 12964 25060 12974
rect 25060 12908 25172 12964
rect 25004 12870 25060 12908
rect 25116 11506 25172 12908
rect 25340 12404 25396 12414
rect 25452 12404 25508 13468
rect 25340 12402 25508 12404
rect 25340 12350 25342 12402
rect 25394 12350 25508 12402
rect 25340 12348 25508 12350
rect 25340 12338 25396 12348
rect 25116 11454 25118 11506
rect 25170 11454 25172 11506
rect 25116 11442 25172 11454
rect 25340 12180 25396 12190
rect 25228 11396 25284 11406
rect 25228 11060 25284 11340
rect 25116 11004 25284 11060
rect 24220 9774 24222 9826
rect 24274 9774 24276 9826
rect 24220 9762 24276 9774
rect 24780 9772 24948 9828
rect 25004 9938 25060 9950
rect 25004 9886 25006 9938
rect 25058 9886 25060 9938
rect 24332 9492 24388 9502
rect 24108 9268 24164 9278
rect 24108 9174 24164 9212
rect 24220 8372 24276 8382
rect 24220 8278 24276 8316
rect 23996 7756 24276 7812
rect 24108 7588 24164 7598
rect 23884 5170 23940 5180
rect 23996 7532 24108 7588
rect 23660 4562 23828 4564
rect 23660 4510 23662 4562
rect 23714 4510 23828 4562
rect 23660 4508 23828 4510
rect 23660 4498 23716 4508
rect 23548 3614 23550 3666
rect 23602 3614 23604 3666
rect 23548 3602 23604 3614
rect 23996 3668 24052 7532
rect 24108 7522 24164 7532
rect 24220 7028 24276 7756
rect 24108 6972 24276 7028
rect 24108 5682 24164 6972
rect 24332 6916 24388 9436
rect 24668 8930 24724 8942
rect 24668 8878 24670 8930
rect 24722 8878 24724 8930
rect 24444 8818 24500 8830
rect 24444 8766 24446 8818
rect 24498 8766 24500 8818
rect 24444 8260 24500 8766
rect 24444 8194 24500 8204
rect 24668 8148 24724 8878
rect 24780 8428 24836 9772
rect 25004 9156 25060 9886
rect 25004 9090 25060 9100
rect 25116 9826 25172 11004
rect 25228 10836 25284 10846
rect 25228 10742 25284 10780
rect 25116 9774 25118 9826
rect 25170 9774 25172 9826
rect 24780 8372 24948 8428
rect 24780 8260 24836 8270
rect 24780 8166 24836 8204
rect 24668 8082 24724 8092
rect 24108 5630 24110 5682
rect 24162 5630 24164 5682
rect 24108 5572 24164 5630
rect 24108 5506 24164 5516
rect 24220 6860 24388 6916
rect 24556 7476 24612 7486
rect 24108 5346 24164 5358
rect 24108 5294 24110 5346
rect 24162 5294 24164 5346
rect 24108 5234 24164 5294
rect 24108 5182 24110 5234
rect 24162 5182 24164 5234
rect 24108 5012 24164 5182
rect 24108 4946 24164 4956
rect 24108 4564 24164 4574
rect 24220 4564 24276 6860
rect 24332 6692 24388 6702
rect 24332 6598 24388 6636
rect 24332 6132 24388 6142
rect 24332 6038 24388 6076
rect 24108 4562 24220 4564
rect 24108 4510 24110 4562
rect 24162 4510 24220 4562
rect 24108 4508 24220 4510
rect 24556 4564 24612 7420
rect 24668 7028 24724 7038
rect 24668 6690 24724 6972
rect 24668 6638 24670 6690
rect 24722 6638 24724 6690
rect 24668 6468 24724 6638
rect 24668 6402 24724 6412
rect 24892 6468 24948 8372
rect 25116 8260 25172 9774
rect 25228 10052 25284 10062
rect 25228 9154 25284 9996
rect 25340 9266 25396 12124
rect 25452 11172 25508 11182
rect 25452 10834 25508 11116
rect 25452 10782 25454 10834
rect 25506 10782 25508 10834
rect 25452 10770 25508 10782
rect 25452 10498 25508 10510
rect 25452 10446 25454 10498
rect 25506 10446 25508 10498
rect 25452 10388 25508 10446
rect 25452 10322 25508 10332
rect 25564 10164 25620 13692
rect 25676 13746 25732 13758
rect 25676 13694 25678 13746
rect 25730 13694 25732 13746
rect 25676 12964 25732 13694
rect 25788 13524 25844 14476
rect 25788 13458 25844 13468
rect 25900 13300 25956 17724
rect 26348 17666 26404 17678
rect 26348 17614 26350 17666
rect 26402 17614 26404 17666
rect 26348 17220 26404 17614
rect 26348 17154 26404 17164
rect 26012 17108 26068 17118
rect 26012 17014 26068 17052
rect 26124 16098 26180 16110
rect 26124 16046 26126 16098
rect 26178 16046 26180 16098
rect 26124 15876 26180 16046
rect 26012 15820 26124 15876
rect 26012 15428 26068 15820
rect 26124 15810 26180 15820
rect 26012 15362 26068 15372
rect 26012 15204 26068 15214
rect 26012 14868 26068 15148
rect 26460 15204 26516 17948
rect 26684 17668 26740 17678
rect 26684 17666 26852 17668
rect 26684 17614 26686 17666
rect 26738 17614 26852 17666
rect 26684 17612 26852 17614
rect 26684 17602 26740 17612
rect 26684 16994 26740 17006
rect 26684 16942 26686 16994
rect 26738 16942 26740 16994
rect 26684 16210 26740 16942
rect 26796 16772 26852 17612
rect 27132 17666 27188 17678
rect 27132 17614 27134 17666
rect 27186 17614 27188 17666
rect 27020 16996 27076 17006
rect 27132 16996 27188 17614
rect 27020 16994 27188 16996
rect 27020 16942 27022 16994
rect 27074 16942 27188 16994
rect 27020 16940 27188 16942
rect 27244 17668 27300 17678
rect 27244 17108 27300 17612
rect 27356 17444 27412 19742
rect 27356 17378 27412 17388
rect 27020 16884 27076 16940
rect 27020 16818 27076 16828
rect 27244 16882 27300 17052
rect 27244 16830 27246 16882
rect 27298 16830 27300 16882
rect 27244 16818 27300 16830
rect 26796 16324 26852 16716
rect 27468 16660 27524 20748
rect 27916 20738 27972 20750
rect 27692 19908 27748 19918
rect 27692 19814 27748 19852
rect 28140 17220 28196 23884
rect 28364 23874 28420 23884
rect 28476 23826 28532 24220
rect 29260 24050 29316 26910
rect 29260 23998 29262 24050
rect 29314 23998 29316 24050
rect 29260 23986 29316 23998
rect 29372 23940 29428 28812
rect 29932 28802 29988 28812
rect 30380 28756 30436 28766
rect 29708 28644 29764 28654
rect 29708 28550 29764 28588
rect 30380 28642 30436 28700
rect 30380 28590 30382 28642
rect 30434 28590 30436 28642
rect 30380 27858 30436 28590
rect 30492 28754 30548 28766
rect 30492 28702 30494 28754
rect 30546 28702 30548 28754
rect 30492 28644 30548 28702
rect 30492 28578 30548 28588
rect 30380 27806 30382 27858
rect 30434 27806 30436 27858
rect 30380 27794 30436 27806
rect 29932 27074 29988 27086
rect 29932 27022 29934 27074
rect 29986 27022 29988 27074
rect 29484 26850 29540 26862
rect 29484 26798 29486 26850
rect 29538 26798 29540 26850
rect 29484 25396 29540 26798
rect 29484 25330 29540 25340
rect 29372 23874 29428 23884
rect 29820 25284 29876 25294
rect 29820 24722 29876 25228
rect 29820 24670 29822 24722
rect 29874 24670 29876 24722
rect 29820 23938 29876 24670
rect 29820 23886 29822 23938
rect 29874 23886 29876 23938
rect 29820 23874 29876 23886
rect 28476 23774 28478 23826
rect 28530 23774 28532 23826
rect 28476 23762 28532 23774
rect 29484 23826 29540 23838
rect 29484 23774 29486 23826
rect 29538 23774 29540 23826
rect 28588 23716 28644 23726
rect 28476 23156 28532 23166
rect 28588 23156 28644 23660
rect 28700 23716 28756 23726
rect 28700 23714 28980 23716
rect 28700 23662 28702 23714
rect 28754 23662 28980 23714
rect 28700 23660 28980 23662
rect 28700 23650 28756 23660
rect 28476 23154 28644 23156
rect 28476 23102 28478 23154
rect 28530 23102 28644 23154
rect 28476 23100 28644 23102
rect 28476 23090 28532 23100
rect 28476 22372 28532 22382
rect 28364 22316 28476 22372
rect 28252 22148 28308 22158
rect 28252 20690 28308 22092
rect 28252 20638 28254 20690
rect 28306 20638 28308 20690
rect 28252 20626 28308 20638
rect 28252 20020 28308 20030
rect 28252 19926 28308 19964
rect 28364 18676 28420 22316
rect 28476 22306 28532 22316
rect 28700 19794 28756 19806
rect 28700 19742 28702 19794
rect 28754 19742 28756 19794
rect 28364 18620 28532 18676
rect 28028 17164 28196 17220
rect 28252 18450 28308 18462
rect 28252 18398 28254 18450
rect 28306 18398 28308 18450
rect 27244 16604 27524 16660
rect 27580 16882 27636 16894
rect 27580 16830 27582 16882
rect 27634 16830 27636 16882
rect 27580 16660 27636 16830
rect 26796 16268 26964 16324
rect 26684 16158 26686 16210
rect 26738 16158 26740 16210
rect 26684 16146 26740 16158
rect 26460 15138 26516 15148
rect 26572 15874 26628 15886
rect 26572 15822 26574 15874
rect 26626 15822 26628 15874
rect 26012 14802 26068 14812
rect 26124 15092 26180 15102
rect 26124 14530 26180 15036
rect 26124 14478 26126 14530
rect 26178 14478 26180 14530
rect 26124 14420 26180 14478
rect 26124 14354 26180 14364
rect 26236 14980 26292 14990
rect 26236 13746 26292 14924
rect 26572 14530 26628 15822
rect 26796 15874 26852 15886
rect 26796 15822 26798 15874
rect 26850 15822 26852 15874
rect 26796 15092 26852 15822
rect 26796 15026 26852 15036
rect 26908 15090 26964 16268
rect 26908 15038 26910 15090
rect 26962 15038 26964 15090
rect 26908 15026 26964 15038
rect 26572 14478 26574 14530
rect 26626 14478 26628 14530
rect 26572 14420 26628 14478
rect 26460 13860 26516 13870
rect 26572 13860 26628 14364
rect 27244 13972 27300 16604
rect 27580 16594 27636 16604
rect 28028 16436 28084 17164
rect 28140 16996 28196 17006
rect 28140 16902 28196 16940
rect 28252 16660 28308 18398
rect 28364 18450 28420 18462
rect 28364 18398 28366 18450
rect 28418 18398 28420 18450
rect 28364 18228 28420 18398
rect 28364 18162 28420 18172
rect 28476 17668 28532 18620
rect 28700 18340 28756 19742
rect 28924 18452 28980 23660
rect 29148 23714 29204 23726
rect 29148 23662 29150 23714
rect 29202 23662 29204 23714
rect 29148 22484 29204 23662
rect 29372 23714 29428 23726
rect 29372 23662 29374 23714
rect 29426 23662 29428 23714
rect 29372 23268 29428 23662
rect 29372 23202 29428 23212
rect 29260 22932 29316 22942
rect 29484 22932 29540 23774
rect 29932 23716 29988 27022
rect 30492 26962 30548 26974
rect 30492 26910 30494 26962
rect 30546 26910 30548 26962
rect 30492 26852 30548 26910
rect 30604 26908 30660 33516
rect 30716 32788 30772 38612
rect 31164 38164 31220 38780
rect 31276 38724 31332 39676
rect 31276 38658 31332 38668
rect 31500 39618 31556 40684
rect 31724 40292 31780 41022
rect 31724 40226 31780 40236
rect 31500 39566 31502 39618
rect 31554 39566 31556 39618
rect 31500 38276 31556 39566
rect 31612 40178 31668 40190
rect 31612 40126 31614 40178
rect 31666 40126 31668 40178
rect 31612 39396 31668 40126
rect 31612 39330 31668 39340
rect 31836 38948 31892 41580
rect 31948 40964 32004 41916
rect 32396 41906 32452 41916
rect 33404 42082 33460 42094
rect 33404 42030 33406 42082
rect 33458 42030 33460 42082
rect 32172 41748 32228 41758
rect 32172 41746 32564 41748
rect 32172 41694 32174 41746
rect 32226 41694 32564 41746
rect 32172 41692 32564 41694
rect 32172 41682 32228 41692
rect 32172 41524 32228 41534
rect 32172 41186 32228 41468
rect 32172 41134 32174 41186
rect 32226 41134 32228 41186
rect 32172 41122 32228 41134
rect 32508 41186 32564 41692
rect 32508 41134 32510 41186
rect 32562 41134 32564 41186
rect 32508 41122 32564 41134
rect 32732 41636 32788 41646
rect 32732 41074 32788 41580
rect 32844 41300 32900 41310
rect 33404 41300 33460 42030
rect 32844 41298 33460 41300
rect 32844 41246 32846 41298
rect 32898 41246 33460 41298
rect 32844 41244 33460 41246
rect 33516 41412 33572 42476
rect 33740 42530 33796 42542
rect 33740 42478 33742 42530
rect 33794 42478 33796 42530
rect 33740 41748 33796 42478
rect 33740 41682 33796 41692
rect 32844 41234 32900 41244
rect 32732 41022 32734 41074
rect 32786 41022 32788 41074
rect 31948 40908 32340 40964
rect 31948 38948 32004 38958
rect 31836 38892 31948 38948
rect 31948 38882 32004 38892
rect 32172 38834 32228 38846
rect 32172 38782 32174 38834
rect 32226 38782 32228 38834
rect 32060 38724 32116 38734
rect 32060 38388 32116 38668
rect 32172 38612 32228 38782
rect 32172 38546 32228 38556
rect 32060 38332 32228 38388
rect 31500 38210 31556 38220
rect 31164 38098 31220 38108
rect 32060 38164 32116 38174
rect 32060 38070 32116 38108
rect 31948 38052 32004 38062
rect 31948 37958 32004 37996
rect 31164 37940 31220 37950
rect 31164 37266 31220 37884
rect 31164 37214 31166 37266
rect 31218 37214 31220 37266
rect 31164 37202 31220 37214
rect 31500 37268 31556 37278
rect 31500 37174 31556 37212
rect 32172 37156 32228 38332
rect 32172 36594 32228 37100
rect 32172 36542 32174 36594
rect 32226 36542 32228 36594
rect 32172 36530 32228 36542
rect 31612 36484 31668 36494
rect 31052 36260 31108 36270
rect 31052 34130 31108 36204
rect 31388 35028 31444 35038
rect 31612 35028 31668 36428
rect 31948 36482 32004 36494
rect 31948 36430 31950 36482
rect 32002 36430 32004 36482
rect 31948 36148 32004 36430
rect 31948 36082 32004 36092
rect 31388 35026 31668 35028
rect 31388 34974 31390 35026
rect 31442 34974 31668 35026
rect 31388 34972 31668 34974
rect 31948 35588 32004 35598
rect 32284 35588 32340 40908
rect 32732 40852 32788 41022
rect 33404 41076 33460 41086
rect 33404 40982 33460 41020
rect 32732 40786 32788 40796
rect 32956 40962 33012 40974
rect 32956 40910 32958 40962
rect 33010 40910 33012 40962
rect 32620 40290 32676 40302
rect 32620 40238 32622 40290
rect 32674 40238 32676 40290
rect 32620 39844 32676 40238
rect 32676 39788 32900 39844
rect 32620 39778 32676 39788
rect 32844 39618 32900 39788
rect 32956 39730 33012 40910
rect 33516 40516 33572 41356
rect 34076 41412 34132 42700
rect 34300 42690 34356 42700
rect 34076 41410 34244 41412
rect 34076 41358 34078 41410
rect 34130 41358 34244 41410
rect 34076 41356 34244 41358
rect 34076 41346 34132 41356
rect 33740 40964 33796 40974
rect 33740 40962 33908 40964
rect 33740 40910 33742 40962
rect 33794 40910 33908 40962
rect 33740 40908 33908 40910
rect 33740 40898 33796 40908
rect 33628 40516 33684 40526
rect 33516 40514 33684 40516
rect 33516 40462 33630 40514
rect 33682 40462 33684 40514
rect 33516 40460 33684 40462
rect 33628 40450 33684 40460
rect 32956 39678 32958 39730
rect 33010 39678 33012 39730
rect 32956 39666 33012 39678
rect 33516 40292 33572 40302
rect 32844 39566 32846 39618
rect 32898 39566 32900 39618
rect 32844 39554 32900 39566
rect 33516 39618 33572 40236
rect 33516 39566 33518 39618
rect 33570 39566 33572 39618
rect 33516 39554 33572 39566
rect 33852 39618 33908 40908
rect 34188 40404 34244 41356
rect 34300 41188 34356 41198
rect 34300 41094 34356 41132
rect 34524 40964 34580 50540
rect 34636 50594 34692 51548
rect 34748 50706 34804 51996
rect 34972 51940 35028 51950
rect 34748 50654 34750 50706
rect 34802 50654 34804 50706
rect 34748 50642 34804 50654
rect 34860 51828 34916 51838
rect 34636 50542 34638 50594
rect 34690 50542 34692 50594
rect 34636 46228 34692 50542
rect 34860 50428 34916 51772
rect 34972 51380 35028 51884
rect 34972 51286 35028 51324
rect 35084 50932 35140 52110
rect 35308 51268 35364 52332
rect 35420 52276 35476 52286
rect 35420 52162 35476 52220
rect 35420 52110 35422 52162
rect 35474 52110 35476 52162
rect 35420 52098 35476 52110
rect 35532 52164 35588 52174
rect 35756 52164 35812 52174
rect 35588 52162 35812 52164
rect 35588 52110 35758 52162
rect 35810 52110 35812 52162
rect 35588 52108 35812 52110
rect 35532 52098 35588 52108
rect 35756 52098 35812 52108
rect 35868 52164 35924 52782
rect 36204 52164 36260 53452
rect 36428 52500 36484 52510
rect 35868 52098 35924 52108
rect 36092 52108 36204 52164
rect 35420 51940 35476 51950
rect 35420 51846 35476 51884
rect 35756 51492 35812 51502
rect 35420 51380 35476 51390
rect 35476 51324 35588 51380
rect 35420 51314 35476 51324
rect 35308 51202 35364 51212
rect 34748 50372 34916 50428
rect 34972 50876 35140 50932
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 34972 50428 35028 50876
rect 35084 50596 35140 50634
rect 35084 50530 35140 50540
rect 35308 50594 35364 50606
rect 35308 50542 35310 50594
rect 35362 50542 35364 50594
rect 34972 50372 35140 50428
rect 34748 49810 34804 50372
rect 34748 49758 34750 49810
rect 34802 49758 34804 49810
rect 34748 49746 34804 49758
rect 34972 49252 35028 49262
rect 34972 49158 35028 49196
rect 35084 48692 35140 50372
rect 35308 49588 35364 50542
rect 35532 49810 35588 51324
rect 35756 50370 35812 51436
rect 36092 50818 36148 52108
rect 36204 52070 36260 52108
rect 36316 52276 36372 52286
rect 36316 51492 36372 52220
rect 36092 50766 36094 50818
rect 36146 50766 36148 50818
rect 36092 50754 36148 50766
rect 36204 51436 36372 51492
rect 36428 51828 36484 52444
rect 36540 51940 36596 51950
rect 36596 51884 36708 51940
rect 36540 51874 36596 51884
rect 35756 50318 35758 50370
rect 35810 50318 35812 50370
rect 35756 50306 35812 50318
rect 35868 50596 35924 50606
rect 35532 49758 35534 49810
rect 35586 49758 35588 49810
rect 35532 49746 35588 49758
rect 35756 49588 35812 49598
rect 35308 49532 35588 49588
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35308 48804 35364 48814
rect 35308 48710 35364 48748
rect 35084 48626 35140 48636
rect 35308 48468 35364 48478
rect 35308 48354 35364 48412
rect 35308 48302 35310 48354
rect 35362 48302 35364 48354
rect 35308 48290 35364 48302
rect 34860 48244 34916 48254
rect 34860 48150 34916 48188
rect 35084 48132 35140 48142
rect 35084 47458 35140 48076
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35084 47406 35086 47458
rect 35138 47406 35140 47458
rect 35084 47394 35140 47406
rect 35308 47684 35364 47694
rect 35532 47684 35588 49532
rect 35644 49026 35700 49038
rect 35644 48974 35646 49026
rect 35698 48974 35700 49026
rect 35644 48916 35700 48974
rect 35644 48850 35700 48860
rect 35308 47458 35364 47628
rect 35308 47406 35310 47458
rect 35362 47406 35364 47458
rect 35308 47394 35364 47406
rect 35420 47628 35588 47684
rect 35644 48692 35700 48702
rect 35644 47682 35700 48636
rect 35756 48354 35812 49532
rect 35868 49138 35924 50540
rect 35868 49086 35870 49138
rect 35922 49086 35924 49138
rect 35868 49074 35924 49086
rect 35980 49364 36036 49374
rect 35756 48302 35758 48354
rect 35810 48302 35812 48354
rect 35756 48290 35812 48302
rect 35644 47630 35646 47682
rect 35698 47630 35700 47682
rect 35420 47234 35476 47628
rect 35644 47618 35700 47630
rect 35868 47460 35924 47470
rect 35980 47460 36036 49308
rect 36204 49026 36260 51436
rect 36428 51378 36484 51772
rect 36652 51492 36708 51884
rect 36764 51716 36820 54908
rect 36876 54628 36932 55468
rect 36988 55300 37044 55310
rect 36988 55206 37044 55244
rect 36876 54514 36932 54572
rect 36876 54462 36878 54514
rect 36930 54462 36932 54514
rect 36876 54450 36932 54462
rect 36988 53732 37044 53742
rect 37100 53732 37156 55804
rect 37212 55412 37268 57038
rect 37660 56644 37716 56654
rect 37212 55346 37268 55356
rect 37548 56642 37716 56644
rect 37548 56590 37662 56642
rect 37714 56590 37716 56642
rect 37548 56588 37716 56590
rect 37324 55188 37380 55198
rect 37212 54628 37268 54638
rect 37212 54534 37268 54572
rect 37324 54516 37380 55132
rect 37436 54516 37492 54526
rect 37324 54514 37492 54516
rect 37324 54462 37438 54514
rect 37490 54462 37492 54514
rect 37324 54460 37492 54462
rect 37436 54450 37492 54460
rect 37044 53676 37156 53732
rect 36988 53666 37044 53676
rect 37212 53508 37268 53518
rect 37100 52388 37156 52398
rect 37100 52294 37156 52332
rect 36988 52164 37044 52174
rect 36988 52070 37044 52108
rect 36764 51660 36932 51716
rect 36764 51492 36820 51502
rect 36652 51490 36820 51492
rect 36652 51438 36766 51490
rect 36818 51438 36820 51490
rect 36652 51436 36820 51438
rect 36764 51426 36820 51436
rect 36428 51326 36430 51378
rect 36482 51326 36484 51378
rect 36428 51314 36484 51326
rect 36316 51268 36372 51278
rect 36316 50820 36372 51212
rect 36316 50706 36372 50764
rect 36316 50654 36318 50706
rect 36370 50654 36372 50706
rect 36316 50642 36372 50654
rect 36204 48974 36206 49026
rect 36258 48974 36260 49026
rect 36204 48962 36260 48974
rect 36316 50484 36372 50494
rect 36876 50428 36932 51660
rect 37212 51604 37268 53452
rect 37212 51538 37268 51548
rect 37436 52836 37492 52846
rect 37100 51380 37156 51390
rect 36092 48916 36148 48926
rect 36092 48822 36148 48860
rect 36092 48244 36148 48254
rect 36316 48244 36372 50428
rect 36652 50372 36932 50428
rect 36988 51378 37156 51380
rect 36988 51326 37102 51378
rect 37154 51326 37156 51378
rect 36988 51324 37156 51326
rect 36988 50428 37044 51324
rect 37100 51314 37156 51324
rect 37100 51156 37156 51166
rect 37100 51154 37380 51156
rect 37100 51102 37102 51154
rect 37154 51102 37380 51154
rect 37100 51100 37380 51102
rect 37100 51090 37156 51100
rect 37324 50482 37380 51100
rect 37436 50708 37492 52780
rect 37436 50642 37492 50652
rect 37324 50430 37326 50482
rect 37378 50430 37380 50482
rect 36988 50372 37156 50428
rect 37324 50418 37380 50430
rect 36652 50148 36708 50372
rect 36652 50082 36708 50092
rect 36652 49924 36708 49934
rect 36540 49922 36708 49924
rect 36540 49870 36654 49922
rect 36706 49870 36708 49922
rect 36540 49868 36708 49870
rect 36540 48466 36596 49868
rect 36652 49858 36708 49868
rect 37100 49138 37156 50372
rect 37548 49924 37604 56588
rect 37660 56578 37716 56588
rect 37772 56532 37828 57486
rect 37772 56466 37828 56476
rect 37996 57540 38052 57550
rect 37996 56642 38052 57484
rect 37996 56590 37998 56642
rect 38050 56590 38052 56642
rect 37884 56084 37940 56094
rect 37772 56082 37940 56084
rect 37772 56030 37886 56082
rect 37938 56030 37940 56082
rect 37772 56028 37940 56030
rect 37660 55972 37716 55982
rect 37660 55878 37716 55916
rect 37772 55300 37828 56028
rect 37884 56018 37940 56028
rect 37772 54738 37828 55244
rect 37996 55076 38052 56590
rect 38444 57204 38500 57214
rect 38444 56306 38500 57148
rect 38556 57090 38612 57102
rect 38556 57038 38558 57090
rect 38610 57038 38612 57090
rect 38556 56978 38612 57038
rect 38556 56926 38558 56978
rect 38610 56926 38612 56978
rect 38556 56914 38612 56926
rect 39564 56980 39620 57820
rect 40012 57874 40068 58156
rect 40684 58212 40740 58222
rect 40012 57822 40014 57874
rect 40066 57822 40068 57874
rect 40012 57810 40068 57822
rect 40236 58100 40292 58110
rect 39564 56886 39620 56924
rect 39340 56756 39396 56766
rect 38892 56642 38948 56654
rect 38892 56590 38894 56642
rect 38946 56590 38948 56642
rect 38444 56254 38446 56306
rect 38498 56254 38500 56306
rect 38444 56242 38500 56254
rect 38556 56420 38612 56430
rect 38556 56306 38612 56364
rect 38556 56254 38558 56306
rect 38610 56254 38612 56306
rect 38332 56082 38388 56094
rect 38332 56030 38334 56082
rect 38386 56030 38388 56082
rect 38332 55972 38388 56030
rect 38332 55906 38388 55916
rect 38556 55468 38612 56254
rect 38892 55636 38948 56590
rect 39004 56644 39060 56654
rect 39004 55972 39060 56588
rect 39004 55906 39060 55916
rect 38892 55570 38948 55580
rect 39004 55748 39060 55758
rect 38556 55412 38836 55468
rect 38892 55412 38948 55422
rect 38780 55410 38948 55412
rect 38780 55358 38894 55410
rect 38946 55358 38948 55410
rect 38780 55356 38948 55358
rect 38892 55346 38948 55356
rect 39004 55298 39060 55692
rect 39004 55246 39006 55298
rect 39058 55246 39060 55298
rect 39004 55234 39060 55246
rect 37996 55010 38052 55020
rect 37772 54686 37774 54738
rect 37826 54686 37828 54738
rect 37772 54674 37828 54686
rect 38892 54964 38948 54974
rect 38444 54628 38500 54638
rect 38108 54516 38164 54526
rect 37996 54514 38164 54516
rect 37996 54462 38110 54514
rect 38162 54462 38164 54514
rect 37996 54460 38164 54462
rect 37660 53620 37716 53630
rect 37660 53526 37716 53564
rect 37996 52834 38052 54460
rect 38108 54450 38164 54460
rect 38444 53396 38500 54572
rect 38892 54402 38948 54908
rect 38892 54350 38894 54402
rect 38946 54350 38948 54402
rect 38780 54292 38836 54302
rect 38668 54290 38836 54292
rect 38668 54238 38782 54290
rect 38834 54238 38836 54290
rect 38668 54236 38836 54238
rect 38668 53956 38724 54236
rect 38780 54226 38836 54236
rect 38892 54180 38948 54350
rect 39340 54738 39396 56700
rect 40236 56756 40292 58044
rect 40572 57876 40628 57886
rect 40236 56690 40292 56700
rect 40460 56756 40516 56766
rect 40124 56642 40180 56654
rect 40124 56590 40126 56642
rect 40178 56590 40180 56642
rect 39452 55972 39508 55982
rect 39452 55878 39508 55916
rect 40124 55970 40180 56590
rect 40460 56196 40516 56700
rect 40460 56130 40516 56140
rect 40124 55918 40126 55970
rect 40178 55918 40180 55970
rect 39676 55300 39732 55310
rect 39676 55206 39732 55244
rect 39340 54686 39342 54738
rect 39394 54686 39396 54738
rect 39340 54290 39396 54686
rect 40124 54628 40180 55918
rect 40124 54562 40180 54572
rect 40460 55972 40516 55982
rect 39788 54404 39844 54414
rect 39340 54238 39342 54290
rect 39394 54238 39396 54290
rect 39340 54226 39396 54238
rect 39564 54402 39844 54404
rect 39564 54350 39790 54402
rect 39842 54350 39844 54402
rect 39564 54348 39844 54350
rect 38892 54114 38948 54124
rect 37996 52782 37998 52834
rect 38050 52782 38052 52834
rect 37996 52770 38052 52782
rect 38332 53340 38444 53396
rect 38108 52724 38164 52734
rect 38108 51490 38164 52668
rect 38332 52276 38388 53340
rect 38444 53330 38500 53340
rect 38556 53900 38724 53956
rect 38556 52836 38612 53900
rect 38556 52770 38612 52780
rect 38668 53732 38724 53742
rect 39452 53732 39508 53742
rect 38668 53060 38724 53676
rect 39116 53730 39508 53732
rect 39116 53678 39454 53730
rect 39506 53678 39508 53730
rect 39116 53676 39508 53678
rect 38780 53508 38836 53518
rect 39116 53508 39172 53676
rect 39452 53666 39508 53676
rect 38780 53506 39172 53508
rect 38780 53454 38782 53506
rect 38834 53454 39172 53506
rect 38780 53452 39172 53454
rect 39228 53506 39284 53518
rect 39228 53454 39230 53506
rect 39282 53454 39284 53506
rect 38780 53442 38836 53452
rect 38444 52722 38500 52734
rect 38444 52670 38446 52722
rect 38498 52670 38500 52722
rect 38444 52500 38500 52670
rect 38444 52434 38500 52444
rect 38556 52612 38612 52622
rect 38332 52220 38500 52276
rect 38108 51438 38110 51490
rect 38162 51438 38164 51490
rect 38108 50428 38164 51438
rect 38332 52052 38388 52062
rect 38332 51490 38388 51996
rect 38444 52050 38500 52220
rect 38444 51998 38446 52050
rect 38498 51998 38500 52050
rect 38444 51986 38500 51998
rect 38332 51438 38334 51490
rect 38386 51438 38388 51490
rect 38332 51426 38388 51438
rect 38108 50372 38388 50428
rect 38332 50036 38388 50372
rect 38444 50036 38500 50046
rect 38332 50034 38500 50036
rect 38332 49982 38446 50034
rect 38498 49982 38500 50034
rect 38332 49980 38500 49982
rect 38444 49970 38500 49980
rect 37100 49086 37102 49138
rect 37154 49086 37156 49138
rect 37100 49074 37156 49086
rect 37436 49364 37492 49374
rect 36876 49028 36932 49038
rect 36876 48934 36932 48972
rect 37212 49028 37268 49038
rect 37212 48916 37268 48972
rect 37436 49026 37492 49308
rect 37436 48974 37438 49026
rect 37490 48974 37492 49026
rect 37436 48962 37492 48974
rect 37100 48860 37268 48916
rect 37324 48914 37380 48926
rect 37324 48862 37326 48914
rect 37378 48862 37380 48914
rect 36652 48804 36708 48814
rect 36708 48748 36820 48804
rect 36652 48738 36708 48748
rect 36540 48414 36542 48466
rect 36594 48414 36596 48466
rect 36540 48402 36596 48414
rect 36652 48354 36708 48366
rect 36652 48302 36654 48354
rect 36706 48302 36708 48354
rect 36092 48242 36372 48244
rect 36092 48190 36094 48242
rect 36146 48190 36372 48242
rect 36092 48188 36372 48190
rect 36428 48242 36484 48254
rect 36428 48190 36430 48242
rect 36482 48190 36484 48242
rect 36092 48178 36148 48188
rect 35868 47458 36036 47460
rect 35868 47406 35870 47458
rect 35922 47406 36036 47458
rect 35868 47404 36036 47406
rect 35868 47394 35924 47404
rect 35420 47182 35422 47234
rect 35474 47182 35476 47234
rect 35420 47170 35476 47182
rect 36316 47234 36372 47246
rect 36316 47182 36318 47234
rect 36370 47182 36372 47234
rect 36316 47012 36372 47182
rect 34972 46564 35028 46574
rect 34972 46470 35028 46508
rect 35756 46452 35812 46462
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34636 45556 34692 46172
rect 35196 45892 35252 45902
rect 34860 45778 34916 45790
rect 34860 45726 34862 45778
rect 34914 45726 34916 45778
rect 34860 45668 34916 45726
rect 35196 45778 35252 45836
rect 35196 45726 35198 45778
rect 35250 45726 35252 45778
rect 35196 45714 35252 45726
rect 35532 45890 35588 45902
rect 35532 45838 35534 45890
rect 35586 45838 35588 45890
rect 34860 45602 34916 45612
rect 34636 45490 34692 45500
rect 35532 45444 35588 45838
rect 35532 45378 35588 45388
rect 35196 45332 35252 45342
rect 34972 45276 35196 45332
rect 34636 45108 34692 45118
rect 34636 44994 34692 45052
rect 34636 44942 34638 44994
rect 34690 44942 34692 44994
rect 34636 42756 34692 44942
rect 34860 44996 34916 45006
rect 34860 44902 34916 44940
rect 34860 44436 34916 44446
rect 34860 43538 34916 44380
rect 34972 44322 35028 45276
rect 35196 45238 35252 45276
rect 35420 45332 35476 45342
rect 35420 45108 35476 45276
rect 35644 45220 35700 45230
rect 35644 45126 35700 45164
rect 35420 45042 35476 45052
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34972 44270 34974 44322
rect 35026 44270 35028 44322
rect 34972 44258 35028 44270
rect 34860 43486 34862 43538
rect 34914 43486 34916 43538
rect 34748 42980 34804 42990
rect 34860 42980 34916 43486
rect 35308 43764 35364 43774
rect 35308 43538 35364 43708
rect 35308 43486 35310 43538
rect 35362 43486 35364 43538
rect 35308 43474 35364 43486
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34748 42978 34916 42980
rect 34748 42926 34750 42978
rect 34802 42926 34916 42978
rect 34748 42924 34916 42926
rect 34748 42914 34804 42924
rect 34636 42700 34916 42756
rect 34748 41860 34804 41870
rect 34748 41186 34804 41804
rect 34748 41134 34750 41186
rect 34802 41134 34804 41186
rect 34748 41122 34804 41134
rect 34860 41188 34916 42700
rect 35084 42754 35140 42766
rect 35084 42702 35086 42754
rect 35138 42702 35140 42754
rect 35084 42196 35140 42702
rect 35308 42644 35364 42654
rect 35644 42644 35700 42654
rect 35308 42550 35364 42588
rect 35532 42642 35700 42644
rect 35532 42590 35646 42642
rect 35698 42590 35700 42642
rect 35532 42588 35700 42590
rect 35196 42196 35252 42206
rect 34860 41122 34916 41132
rect 34972 42194 35252 42196
rect 34972 42142 35198 42194
rect 35250 42142 35252 42194
rect 34972 42140 35252 42142
rect 34972 41074 35028 42140
rect 35196 42130 35252 42140
rect 35532 41972 35588 42588
rect 35644 42578 35700 42588
rect 34972 41022 34974 41074
rect 35026 41022 35028 41074
rect 34972 41010 35028 41022
rect 35084 41748 35140 41758
rect 35084 41076 35140 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35532 41412 35588 41916
rect 35644 41860 35700 41870
rect 35644 41766 35700 41804
rect 35532 41318 35588 41356
rect 34524 40898 34580 40908
rect 34972 40852 35028 40862
rect 34188 40338 34244 40348
rect 34860 40404 34916 40414
rect 34860 40310 34916 40348
rect 34636 40292 34692 40302
rect 33852 39566 33854 39618
rect 33906 39566 33908 39618
rect 33852 39554 33908 39566
rect 34524 39844 34580 39854
rect 33964 39508 34020 39518
rect 33964 39414 34020 39452
rect 32508 39396 32564 39406
rect 33068 39396 33124 39406
rect 32508 39394 32676 39396
rect 32508 39342 32510 39394
rect 32562 39342 32676 39394
rect 32508 39340 32676 39342
rect 32508 39330 32564 39340
rect 32508 38836 32564 38874
rect 32620 38836 32676 39340
rect 33068 39394 33236 39396
rect 33068 39342 33070 39394
rect 33122 39342 33236 39394
rect 33068 39340 33236 39342
rect 33068 39330 33124 39340
rect 33180 38948 33236 39340
rect 34188 38948 34244 38958
rect 33180 38892 33348 38948
rect 32956 38836 33012 38846
rect 32620 38834 33012 38836
rect 32620 38782 32958 38834
rect 33010 38782 33012 38834
rect 32620 38780 33012 38782
rect 32508 38770 32564 38780
rect 32956 38500 33012 38780
rect 33180 38722 33236 38734
rect 33180 38670 33182 38722
rect 33234 38670 33236 38722
rect 33180 38668 33236 38670
rect 32956 38434 33012 38444
rect 33068 38612 33236 38668
rect 32956 38276 33012 38286
rect 32956 37938 33012 38220
rect 32956 37886 32958 37938
rect 33010 37886 33012 37938
rect 32956 37874 33012 37886
rect 32508 37492 32564 37502
rect 32508 35924 32564 37436
rect 32956 36370 33012 36382
rect 32956 36318 32958 36370
rect 33010 36318 33012 36370
rect 32508 35922 32900 35924
rect 32508 35870 32510 35922
rect 32562 35870 32900 35922
rect 32508 35868 32900 35870
rect 32508 35858 32564 35868
rect 31948 35586 32340 35588
rect 31948 35534 31950 35586
rect 32002 35534 32340 35586
rect 31948 35532 32340 35534
rect 31388 34962 31444 34972
rect 31836 34914 31892 34926
rect 31836 34862 31838 34914
rect 31890 34862 31892 34914
rect 31836 34804 31892 34862
rect 31724 34132 31780 34142
rect 31052 34078 31054 34130
rect 31106 34078 31108 34130
rect 31052 34066 31108 34078
rect 31388 34130 31780 34132
rect 31388 34078 31726 34130
rect 31778 34078 31780 34130
rect 31388 34076 31780 34078
rect 30828 34018 30884 34030
rect 30828 33966 30830 34018
rect 30882 33966 30884 34018
rect 30828 33348 30884 33966
rect 31388 34018 31444 34076
rect 31724 34066 31780 34076
rect 31388 33966 31390 34018
rect 31442 33966 31444 34018
rect 31388 33954 31444 33966
rect 31836 33908 31892 34748
rect 30828 33282 30884 33292
rect 31500 33852 31892 33908
rect 31164 33012 31220 33022
rect 30716 32732 30884 32788
rect 30716 31668 30772 31678
rect 30716 31218 30772 31612
rect 30716 31166 30718 31218
rect 30770 31166 30772 31218
rect 30716 31154 30772 31166
rect 30604 26852 30772 26908
rect 30492 26786 30548 26796
rect 30492 26290 30548 26302
rect 30492 26238 30494 26290
rect 30546 26238 30548 26290
rect 30492 26068 30548 26238
rect 30380 26012 30492 26068
rect 30044 25284 30100 25294
rect 30044 25190 30100 25228
rect 30380 24946 30436 26012
rect 30492 26002 30548 26012
rect 30380 24894 30382 24946
rect 30434 24894 30436 24946
rect 30380 24276 30436 24894
rect 30492 25732 30548 25742
rect 30492 24946 30548 25676
rect 30492 24894 30494 24946
rect 30546 24894 30548 24946
rect 30492 24882 30548 24894
rect 30604 24948 30660 24958
rect 30604 24854 30660 24892
rect 30380 24210 30436 24220
rect 30716 23940 30772 26852
rect 30828 26852 30884 32732
rect 30940 31892 30996 31902
rect 30940 30324 30996 31836
rect 31164 31668 31220 32956
rect 31500 32786 31556 33852
rect 31724 33460 31780 33470
rect 31724 33346 31780 33404
rect 31724 33294 31726 33346
rect 31778 33294 31780 33346
rect 31724 33282 31780 33294
rect 31836 33348 31892 33358
rect 31500 32734 31502 32786
rect 31554 32734 31556 32786
rect 31500 32722 31556 32734
rect 31836 32564 31892 33292
rect 31836 32470 31892 32508
rect 31948 32004 32004 35532
rect 32396 34356 32452 34366
rect 32396 34262 32452 34300
rect 32172 34242 32228 34254
rect 32172 34190 32174 34242
rect 32226 34190 32228 34242
rect 32060 33236 32116 33246
rect 32060 32562 32116 33180
rect 32172 33124 32228 34190
rect 32172 33058 32228 33068
rect 32284 34242 32340 34254
rect 32284 34190 32286 34242
rect 32338 34190 32340 34242
rect 32284 33012 32340 34190
rect 32508 34130 32564 34142
rect 32508 34078 32510 34130
rect 32562 34078 32564 34130
rect 32508 33684 32564 34078
rect 32508 33618 32564 33628
rect 32732 33460 32788 33470
rect 32732 33366 32788 33404
rect 32284 32956 32452 33012
rect 32060 32510 32062 32562
rect 32114 32510 32116 32562
rect 32060 32498 32116 32510
rect 32172 32900 32228 32910
rect 31948 31938 32004 31948
rect 31164 31666 31556 31668
rect 31164 31614 31166 31666
rect 31218 31614 31556 31666
rect 31164 31612 31556 31614
rect 31164 31602 31220 31612
rect 31164 31220 31220 31230
rect 31164 31126 31220 31164
rect 31500 30994 31556 31612
rect 31500 30942 31502 30994
rect 31554 30942 31556 30994
rect 31500 30930 31556 30942
rect 31948 31444 32004 31454
rect 30940 30230 30996 30268
rect 31836 30324 31892 30334
rect 31164 30210 31220 30222
rect 31164 30158 31166 30210
rect 31218 30158 31220 30210
rect 31164 29426 31220 30158
rect 31836 29652 31892 30268
rect 31948 29988 32004 31388
rect 32172 31106 32228 32844
rect 32396 31668 32452 32956
rect 32508 32452 32564 32462
rect 32508 31668 32564 32396
rect 32732 31668 32788 31678
rect 32508 31666 32788 31668
rect 32508 31614 32734 31666
rect 32786 31614 32788 31666
rect 32508 31612 32788 31614
rect 32396 31602 32452 31612
rect 32172 31054 32174 31106
rect 32226 31054 32228 31106
rect 32172 31042 32228 31054
rect 32284 31554 32340 31566
rect 32284 31502 32286 31554
rect 32338 31502 32340 31554
rect 32284 31220 32340 31502
rect 32732 31556 32788 31612
rect 32732 31490 32788 31500
rect 32844 31444 32900 35868
rect 32956 35252 33012 36318
rect 33068 36260 33124 38612
rect 33292 38052 33348 38892
rect 33404 38836 33460 38846
rect 33404 38742 33460 38780
rect 33516 38834 33572 38846
rect 33516 38782 33518 38834
rect 33570 38782 33572 38834
rect 33292 37986 33348 37996
rect 33404 38164 33460 38174
rect 33404 37266 33460 38108
rect 33404 37214 33406 37266
rect 33458 37214 33460 37266
rect 33404 37202 33460 37214
rect 33068 36194 33124 36204
rect 33180 37044 33236 37054
rect 33516 37044 33572 38782
rect 34188 38274 34244 38892
rect 34188 38222 34190 38274
rect 34242 38222 34244 38274
rect 34188 38210 34244 38222
rect 34300 38500 34356 38510
rect 34524 38500 34580 39788
rect 34636 38668 34692 40236
rect 34972 39396 35028 40796
rect 35084 39620 35140 41020
rect 35756 40740 35812 46396
rect 36316 45892 36372 46956
rect 36428 46900 36484 48190
rect 36652 48244 36708 48302
rect 36764 48354 36820 48748
rect 36764 48302 36766 48354
rect 36818 48302 36820 48354
rect 36764 48290 36820 48302
rect 36652 47460 36708 48188
rect 36652 47394 36708 47404
rect 36428 46834 36484 46844
rect 36988 47348 37044 47358
rect 36316 45826 36372 45836
rect 35868 45666 35924 45678
rect 36540 45668 36596 45678
rect 35868 45614 35870 45666
rect 35922 45614 35924 45666
rect 35868 45220 35924 45614
rect 35868 45154 35924 45164
rect 36428 45666 36596 45668
rect 36428 45614 36542 45666
rect 36594 45614 36596 45666
rect 36428 45612 36596 45614
rect 36316 45108 36372 45118
rect 36428 45108 36484 45612
rect 36540 45602 36596 45612
rect 36372 45052 36484 45108
rect 36540 45218 36596 45230
rect 36540 45166 36542 45218
rect 36594 45166 36596 45218
rect 36316 45042 36372 45052
rect 36316 44548 36372 44558
rect 36540 44548 36596 45166
rect 36316 44546 36540 44548
rect 36316 44494 36318 44546
rect 36370 44494 36540 44546
rect 36316 44492 36540 44494
rect 36316 44482 36372 44492
rect 36540 44454 36596 44492
rect 36876 45108 36932 45118
rect 36204 44324 36260 44334
rect 36204 44230 36260 44268
rect 36876 43652 36932 45052
rect 36988 44212 37044 47292
rect 37100 46562 37156 48860
rect 37324 48804 37380 48862
rect 37324 48738 37380 48748
rect 37436 48468 37492 48478
rect 37548 48468 37604 49868
rect 37884 49812 37940 49822
rect 38556 49812 38612 52556
rect 38668 51378 38724 53004
rect 39004 53058 39060 53452
rect 39004 53006 39006 53058
rect 39058 53006 39060 53058
rect 39004 52994 39060 53006
rect 38780 52724 38836 52734
rect 38780 52630 38836 52668
rect 38668 51326 38670 51378
rect 38722 51326 38724 51378
rect 38668 51314 38724 51326
rect 38892 52164 38948 52174
rect 38892 49922 38948 52108
rect 39228 52164 39284 53454
rect 39340 53060 39396 53070
rect 39340 52966 39396 53004
rect 39228 52098 39284 52108
rect 39564 51828 39620 54348
rect 39788 54338 39844 54348
rect 40236 54402 40292 54414
rect 40236 54350 40238 54402
rect 40290 54350 40292 54402
rect 40012 53732 40068 53742
rect 40012 53638 40068 53676
rect 39788 53004 40180 53060
rect 39788 51940 39844 53004
rect 40124 52946 40180 53004
rect 40124 52894 40126 52946
rect 40178 52894 40180 52946
rect 40124 52882 40180 52894
rect 40012 52836 40068 52846
rect 39228 51772 39620 51828
rect 39676 51938 39844 51940
rect 39676 51886 39790 51938
rect 39842 51886 39844 51938
rect 39676 51884 39844 51886
rect 39004 51154 39060 51166
rect 39004 51102 39006 51154
rect 39058 51102 39060 51154
rect 39004 50596 39060 51102
rect 39004 50530 39060 50540
rect 39116 50820 39172 50830
rect 39116 50370 39172 50764
rect 39116 50318 39118 50370
rect 39170 50318 39172 50370
rect 39116 50306 39172 50318
rect 39228 50708 39284 51772
rect 38892 49870 38894 49922
rect 38946 49870 38948 49922
rect 38892 49858 38948 49870
rect 37492 48412 37604 48468
rect 37660 49252 37716 49262
rect 37660 48466 37716 49196
rect 37884 49252 37940 49756
rect 37884 49186 37940 49196
rect 38444 49756 38612 49812
rect 38108 49028 38164 49038
rect 38108 48934 38164 48972
rect 37884 48804 37940 48814
rect 37884 48802 38276 48804
rect 37884 48750 37886 48802
rect 37938 48750 38276 48802
rect 37884 48748 38276 48750
rect 37884 48738 37940 48748
rect 37660 48414 37662 48466
rect 37714 48414 37716 48466
rect 37212 48244 37268 48254
rect 37212 48150 37268 48188
rect 37436 48242 37492 48412
rect 37660 48402 37716 48414
rect 37772 48580 37828 48590
rect 37436 48190 37438 48242
rect 37490 48190 37492 48242
rect 37436 48178 37492 48190
rect 37772 48242 37828 48524
rect 37772 48190 37774 48242
rect 37826 48190 37828 48242
rect 37772 48178 37828 48190
rect 38108 48580 38164 48590
rect 38108 48242 38164 48524
rect 38108 48190 38110 48242
rect 38162 48190 38164 48242
rect 38108 48020 38164 48190
rect 38108 47954 38164 47964
rect 37884 47908 37940 47918
rect 37660 47852 37884 47908
rect 37212 47684 37268 47694
rect 37212 47348 37268 47628
rect 37660 47460 37716 47852
rect 37884 47842 37940 47852
rect 37996 47572 38052 47582
rect 37212 47254 37268 47292
rect 37324 47458 37716 47460
rect 37324 47406 37662 47458
rect 37714 47406 37716 47458
rect 37324 47404 37716 47406
rect 37100 46510 37102 46562
rect 37154 46510 37156 46562
rect 37100 46498 37156 46510
rect 37324 46340 37380 47404
rect 37660 47394 37716 47404
rect 37772 47570 38052 47572
rect 37772 47518 37998 47570
rect 38050 47518 38052 47570
rect 37772 47516 38052 47518
rect 37100 46284 37380 46340
rect 37100 46114 37156 46284
rect 37100 46062 37102 46114
rect 37154 46062 37156 46114
rect 37100 46050 37156 46062
rect 37548 45556 37604 45566
rect 37212 45108 37268 45118
rect 37100 44996 37156 45006
rect 37100 44322 37156 44940
rect 37100 44270 37102 44322
rect 37154 44270 37156 44322
rect 37100 44258 37156 44270
rect 36988 44146 37044 44156
rect 36876 43586 36932 43596
rect 36988 43650 37044 43662
rect 36988 43598 36990 43650
rect 37042 43598 37044 43650
rect 36652 43540 36708 43550
rect 36652 43446 36708 43484
rect 36540 42532 36596 42542
rect 36428 42530 36596 42532
rect 36428 42478 36542 42530
rect 36594 42478 36596 42530
rect 36428 42476 36596 42478
rect 35756 40674 35812 40684
rect 35868 40964 35924 40974
rect 35644 40402 35700 40414
rect 35644 40350 35646 40402
rect 35698 40350 35700 40402
rect 35420 40292 35476 40302
rect 35420 40198 35476 40236
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35644 39732 35700 40350
rect 35644 39676 35812 39732
rect 35084 39618 35588 39620
rect 35084 39566 35086 39618
rect 35138 39566 35588 39618
rect 35084 39564 35588 39566
rect 35084 39554 35140 39564
rect 34972 39340 35140 39396
rect 34636 38612 34916 38668
rect 34524 38444 34692 38500
rect 34076 38052 34132 38062
rect 34076 37958 34132 37996
rect 34076 37716 34132 37726
rect 33180 37042 33572 37044
rect 33180 36990 33182 37042
rect 33234 36990 33572 37042
rect 33180 36988 33572 36990
rect 33628 37266 33684 37278
rect 33628 37214 33630 37266
rect 33682 37214 33684 37266
rect 33628 37044 33684 37214
rect 33852 37156 33908 37166
rect 33852 37062 33908 37100
rect 33684 36988 33796 37044
rect 33180 35698 33236 36988
rect 33628 36978 33684 36988
rect 33740 36708 33796 36988
rect 33740 36652 34020 36708
rect 33852 35812 33908 35822
rect 33628 35810 33908 35812
rect 33628 35758 33854 35810
rect 33906 35758 33908 35810
rect 33628 35756 33908 35758
rect 33180 35646 33182 35698
rect 33234 35646 33236 35698
rect 33180 35634 33236 35646
rect 33516 35698 33572 35710
rect 33516 35646 33518 35698
rect 33570 35646 33572 35698
rect 33012 35196 33124 35252
rect 32956 35186 33012 35196
rect 33068 34914 33124 35196
rect 33068 34862 33070 34914
rect 33122 34862 33124 34914
rect 33068 34850 33124 34862
rect 33180 34356 33236 34366
rect 33236 34300 33460 34356
rect 33180 34290 33236 34300
rect 33404 34242 33460 34300
rect 33404 34190 33406 34242
rect 33458 34190 33460 34242
rect 33404 34178 33460 34190
rect 33068 33348 33124 33358
rect 33068 33254 33124 33292
rect 33292 33236 33348 33246
rect 33292 33142 33348 33180
rect 33516 33012 33572 35646
rect 33404 32956 33572 33012
rect 33068 32562 33124 32574
rect 33292 32564 33348 32574
rect 33404 32564 33460 32956
rect 33516 32788 33572 32798
rect 33516 32694 33572 32732
rect 33068 32510 33070 32562
rect 33122 32510 33124 32562
rect 33068 32452 33124 32510
rect 33068 32386 33124 32396
rect 33180 32562 33460 32564
rect 33180 32510 33294 32562
rect 33346 32510 33460 32562
rect 33180 32508 33460 32510
rect 32956 31668 33012 31678
rect 33180 31668 33236 32508
rect 33292 32498 33348 32508
rect 33628 32340 33684 35756
rect 33852 35746 33908 35756
rect 33964 34914 34020 36652
rect 34076 35140 34132 37660
rect 34188 37268 34244 37278
rect 34188 35812 34244 37212
rect 34300 36820 34356 38444
rect 34412 38164 34468 38174
rect 34636 38164 34692 38444
rect 34412 38162 34692 38164
rect 34412 38110 34414 38162
rect 34466 38110 34692 38162
rect 34412 38108 34692 38110
rect 34412 37044 34468 38108
rect 34860 38050 34916 38612
rect 34860 37998 34862 38050
rect 34914 37998 34916 38050
rect 34860 37986 34916 37998
rect 35084 38050 35140 39340
rect 35532 38834 35588 39564
rect 35532 38782 35534 38834
rect 35586 38782 35588 38834
rect 35532 38770 35588 38782
rect 35756 38668 35812 39676
rect 35868 39508 35924 40908
rect 36092 40516 36148 40526
rect 35980 39508 36036 39518
rect 35868 39506 36036 39508
rect 35868 39454 35982 39506
rect 36034 39454 36036 39506
rect 35868 39452 36036 39454
rect 35980 38834 36036 39452
rect 35980 38782 35982 38834
rect 36034 38782 36036 38834
rect 35980 38770 36036 38782
rect 35532 38612 35812 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35084 37998 35086 38050
rect 35138 37998 35140 38050
rect 35084 37986 35140 37998
rect 34636 37940 34692 37950
rect 34412 36978 34468 36988
rect 34524 37492 34580 37502
rect 34300 36764 34468 36820
rect 34188 35810 34356 35812
rect 34188 35758 34190 35810
rect 34242 35758 34356 35810
rect 34188 35756 34356 35758
rect 34188 35746 34244 35756
rect 34132 35084 34244 35140
rect 34076 35074 34132 35084
rect 33964 34862 33966 34914
rect 34018 34862 34020 34914
rect 33964 34850 34020 34862
rect 33292 32338 33684 32340
rect 33292 32286 33630 32338
rect 33682 32286 33684 32338
rect 33292 32284 33684 32286
rect 33292 32002 33348 32284
rect 33628 32274 33684 32284
rect 33740 33348 33796 33358
rect 33740 33234 33796 33292
rect 33740 33182 33742 33234
rect 33794 33182 33796 33234
rect 33292 31950 33294 32002
rect 33346 31950 33348 32002
rect 33292 31938 33348 31950
rect 33012 31612 33236 31668
rect 33404 31780 33460 31790
rect 33740 31780 33796 33182
rect 33852 33122 33908 33134
rect 33852 33070 33854 33122
rect 33906 33070 33908 33122
rect 33852 32564 33908 33070
rect 33852 32470 33908 32508
rect 34188 32004 34244 35084
rect 34300 35028 34356 35756
rect 34412 35700 34468 36764
rect 34524 36370 34580 37436
rect 34524 36318 34526 36370
rect 34578 36318 34580 36370
rect 34524 36306 34580 36318
rect 34412 35606 34468 35644
rect 34412 35028 34468 35038
rect 34300 35026 34468 35028
rect 34300 34974 34414 35026
rect 34466 34974 34468 35026
rect 34300 34972 34468 34974
rect 34412 34962 34468 34972
rect 34412 33348 34468 33358
rect 34412 33254 34468 33292
rect 34300 33234 34356 33246
rect 34300 33182 34302 33234
rect 34354 33182 34356 33234
rect 34300 33012 34356 33182
rect 34524 33236 34580 33246
rect 34412 33012 34468 33022
rect 34300 32956 34412 33012
rect 34412 32946 34468 32956
rect 34524 32786 34580 33180
rect 34524 32734 34526 32786
rect 34578 32734 34580 32786
rect 34188 31910 34244 31948
rect 34300 32452 34356 32462
rect 33404 31778 33740 31780
rect 33404 31726 33406 31778
rect 33458 31726 33740 31778
rect 33404 31724 33740 31726
rect 32956 31574 33012 31612
rect 32844 31378 32900 31388
rect 33068 31220 33124 31230
rect 32284 31218 33124 31220
rect 32284 31166 33070 31218
rect 33122 31166 33124 31218
rect 32284 31164 33124 31166
rect 32284 30994 32340 31164
rect 33068 31154 33124 31164
rect 33404 31218 33460 31724
rect 33740 31686 33796 31724
rect 34300 31778 34356 32396
rect 34524 32452 34580 32734
rect 34524 32386 34580 32396
rect 34300 31726 34302 31778
rect 34354 31726 34356 31778
rect 34300 31714 34356 31726
rect 34524 31668 34580 31678
rect 34524 31574 34580 31612
rect 33404 31166 33406 31218
rect 33458 31166 33460 31218
rect 33404 31154 33460 31166
rect 33516 31554 33572 31566
rect 33516 31502 33518 31554
rect 33570 31502 33572 31554
rect 32284 30942 32286 30994
rect 32338 30942 32340 30994
rect 32284 30930 32340 30942
rect 32060 30434 32116 30446
rect 32060 30382 32062 30434
rect 32114 30382 32116 30434
rect 32060 30100 32116 30382
rect 33516 30212 33572 31502
rect 33852 31556 33908 31566
rect 33852 31218 33908 31500
rect 33852 31166 33854 31218
rect 33906 31166 33908 31218
rect 33852 31154 33908 31166
rect 34636 31108 34692 37884
rect 35084 37828 35140 37838
rect 35084 36708 35140 37772
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35084 36652 35252 36708
rect 34972 36484 35028 36494
rect 34860 36372 34916 36382
rect 34860 36278 34916 36316
rect 34972 35812 35028 36428
rect 35084 36482 35140 36494
rect 35084 36430 35086 36482
rect 35138 36430 35140 36482
rect 35084 36148 35140 36430
rect 35084 36082 35140 36092
rect 35196 35922 35252 36652
rect 35420 36260 35476 36270
rect 35420 36166 35476 36204
rect 35196 35870 35198 35922
rect 35250 35870 35252 35922
rect 35196 35858 35252 35870
rect 35420 35924 35476 35934
rect 35420 35830 35476 35868
rect 35084 35812 35140 35822
rect 34972 35810 35140 35812
rect 34972 35758 35086 35810
rect 35138 35758 35140 35810
rect 34972 35756 35140 35758
rect 35084 35746 35140 35756
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35308 35028 35364 35038
rect 35532 35028 35588 38612
rect 36092 38052 36148 40460
rect 36428 39844 36484 42476
rect 36540 42466 36596 42476
rect 36764 42082 36820 42094
rect 36764 42030 36766 42082
rect 36818 42030 36820 42082
rect 36764 41972 36820 42030
rect 36764 41906 36820 41916
rect 36988 41412 37044 43598
rect 37212 43540 37268 45052
rect 37436 44548 37492 44558
rect 37324 44324 37380 44334
rect 37324 44210 37380 44268
rect 37324 44158 37326 44210
rect 37378 44158 37380 44210
rect 37324 44146 37380 44158
rect 37436 44210 37492 44492
rect 37436 44158 37438 44210
rect 37490 44158 37492 44210
rect 37436 44146 37492 44158
rect 37548 44100 37604 45500
rect 37772 44324 37828 47516
rect 37996 47506 38052 47516
rect 38220 46898 38276 48748
rect 38444 48356 38500 49756
rect 38780 49588 38836 49598
rect 38780 49494 38836 49532
rect 38556 49028 38612 49038
rect 38556 48934 38612 48972
rect 38892 48802 38948 48814
rect 38892 48750 38894 48802
rect 38946 48750 38948 48802
rect 38444 48300 38612 48356
rect 38444 48130 38500 48142
rect 38444 48078 38446 48130
rect 38498 48078 38500 48130
rect 38444 47908 38500 48078
rect 38444 47842 38500 47852
rect 38220 46846 38222 46898
rect 38274 46846 38276 46898
rect 38220 45780 38276 46846
rect 38220 45686 38276 45724
rect 38556 45332 38612 48300
rect 38220 45276 38612 45332
rect 38780 48130 38836 48142
rect 38780 48078 38782 48130
rect 38834 48078 38836 48130
rect 38780 46788 38836 48078
rect 38892 47348 38948 48750
rect 39228 48468 39284 50652
rect 39452 51490 39508 51502
rect 39452 51438 39454 51490
rect 39506 51438 39508 51490
rect 39452 50428 39508 51438
rect 39564 50484 39620 50494
rect 39452 50372 39620 50428
rect 39340 49586 39396 49598
rect 39340 49534 39342 49586
rect 39394 49534 39396 49586
rect 39340 49026 39396 49534
rect 39340 48974 39342 49026
rect 39394 48974 39396 49026
rect 39340 48962 39396 48974
rect 39452 48916 39508 48926
rect 39452 48822 39508 48860
rect 39228 48402 39284 48412
rect 39564 48244 39620 50372
rect 39676 50484 39732 51884
rect 39788 51874 39844 51884
rect 39900 52834 40068 52836
rect 39900 52782 40014 52834
rect 40066 52782 40068 52834
rect 39900 52780 40068 52782
rect 39788 51604 39844 51614
rect 39900 51604 39956 52780
rect 40012 52770 40068 52780
rect 39788 51602 39900 51604
rect 39788 51550 39790 51602
rect 39842 51550 39900 51602
rect 39788 51548 39900 51550
rect 39788 51538 39844 51548
rect 39900 51510 39956 51548
rect 40236 51602 40292 54350
rect 40460 53956 40516 55916
rect 40572 55298 40628 57820
rect 40684 56866 40740 58156
rect 40796 58210 40852 58222
rect 40796 58158 40798 58210
rect 40850 58158 40852 58210
rect 40796 56980 40852 58158
rect 41132 58212 41188 58222
rect 41188 58156 41524 58212
rect 41132 58118 41188 58156
rect 41244 57540 41300 57550
rect 41244 57446 41300 57484
rect 40908 56980 40964 56990
rect 40796 56924 40908 56980
rect 40684 56814 40686 56866
rect 40738 56814 40740 56866
rect 40684 56802 40740 56814
rect 40908 56866 40964 56924
rect 41356 56980 41412 56990
rect 41356 56886 41412 56924
rect 40908 56814 40910 56866
rect 40962 56814 40964 56866
rect 40908 56802 40964 56814
rect 41468 56866 41524 58156
rect 42252 57876 42308 57886
rect 42252 57782 42308 57820
rect 43708 57874 43764 58380
rect 47516 58324 47572 58334
rect 44380 58212 44436 58222
rect 44492 58212 44548 58222
rect 44380 58210 44492 58212
rect 44380 58158 44382 58210
rect 44434 58158 44492 58210
rect 44380 58156 44492 58158
rect 44380 58146 44436 58156
rect 43708 57822 43710 57874
rect 43762 57822 43764 57874
rect 43708 57810 43764 57822
rect 41804 57540 41860 57550
rect 41468 56814 41470 56866
rect 41522 56814 41524 56866
rect 41468 56802 41524 56814
rect 41580 57538 41860 57540
rect 41580 57486 41806 57538
rect 41858 57486 41860 57538
rect 41580 57484 41860 57486
rect 40572 55246 40574 55298
rect 40626 55246 40628 55298
rect 40572 55234 40628 55246
rect 40796 56642 40852 56654
rect 40796 56590 40798 56642
rect 40850 56590 40852 56642
rect 40796 55300 40852 56590
rect 41020 55970 41076 55982
rect 41020 55918 41022 55970
rect 41074 55918 41076 55970
rect 41020 55748 41076 55918
rect 41468 55972 41524 55982
rect 41468 55878 41524 55916
rect 41020 55682 41076 55692
rect 41020 55524 41076 55534
rect 41020 55430 41076 55468
rect 40796 55234 40852 55244
rect 41356 54514 41412 54526
rect 41356 54462 41358 54514
rect 41410 54462 41412 54514
rect 41132 54404 41188 54414
rect 40460 53890 40516 53900
rect 41020 54402 41188 54404
rect 41020 54350 41134 54402
rect 41186 54350 41188 54402
rect 41020 54348 41188 54350
rect 40348 53676 40852 53732
rect 40348 52164 40404 53676
rect 40796 53620 40852 53676
rect 40908 53620 40964 53630
rect 40796 53618 40964 53620
rect 40796 53566 40910 53618
rect 40962 53566 40964 53618
rect 40796 53564 40964 53566
rect 40908 53554 40964 53564
rect 40684 53506 40740 53518
rect 40684 53454 40686 53506
rect 40738 53454 40740 53506
rect 40348 52162 40516 52164
rect 40348 52110 40350 52162
rect 40402 52110 40516 52162
rect 40348 52108 40516 52110
rect 40348 52098 40404 52108
rect 40236 51550 40238 51602
rect 40290 51550 40292 51602
rect 39788 50820 39844 50830
rect 39788 50706 39844 50764
rect 39788 50654 39790 50706
rect 39842 50654 39844 50706
rect 39788 50642 39844 50654
rect 40124 50820 40180 50830
rect 40012 50594 40068 50606
rect 40012 50542 40014 50594
rect 40066 50542 40068 50594
rect 40012 50484 40068 50542
rect 39676 50428 40068 50484
rect 39676 49586 39732 50428
rect 39900 49812 39956 49822
rect 40124 49812 40180 50764
rect 39900 49810 40180 49812
rect 39900 49758 39902 49810
rect 39954 49758 40180 49810
rect 39900 49756 40180 49758
rect 39900 49746 39956 49756
rect 39676 49534 39678 49586
rect 39730 49534 39732 49586
rect 39676 48692 39732 49534
rect 39676 48626 39732 48636
rect 40236 48580 40292 51550
rect 40348 50706 40404 50718
rect 40348 50654 40350 50706
rect 40402 50654 40404 50706
rect 40348 50372 40404 50654
rect 40348 50306 40404 50316
rect 40348 49924 40404 49934
rect 40348 49830 40404 49868
rect 40236 48514 40292 48524
rect 40124 48468 40180 48478
rect 40012 48356 40068 48394
rect 40124 48374 40180 48412
rect 40012 48290 40068 48300
rect 39564 48150 39620 48188
rect 40348 48244 40404 48254
rect 40348 48150 40404 48188
rect 39228 48130 39284 48142
rect 39228 48078 39230 48130
rect 39282 48078 39284 48130
rect 39228 47572 39284 48078
rect 40012 48132 40068 48142
rect 40012 48038 40068 48076
rect 39228 47506 39284 47516
rect 40236 47908 40292 47918
rect 40012 47460 40068 47470
rect 39116 47348 39172 47358
rect 38892 47292 39116 47348
rect 39116 47254 39172 47292
rect 38108 45106 38164 45118
rect 38108 45054 38110 45106
rect 38162 45054 38164 45106
rect 37996 44884 38052 44894
rect 37884 44548 37940 44558
rect 37884 44434 37940 44492
rect 37884 44382 37886 44434
rect 37938 44382 37940 44434
rect 37884 44370 37940 44382
rect 37548 44034 37604 44044
rect 37660 44322 37828 44324
rect 37660 44270 37774 44322
rect 37826 44270 37828 44322
rect 37660 44268 37828 44270
rect 37324 43540 37380 43550
rect 37212 43538 37380 43540
rect 37212 43486 37326 43538
rect 37378 43486 37380 43538
rect 37212 43484 37380 43486
rect 37324 43474 37380 43484
rect 37660 43540 37716 44268
rect 37772 44258 37828 44268
rect 37884 44212 37940 44222
rect 37660 42754 37716 43484
rect 37660 42702 37662 42754
rect 37714 42702 37716 42754
rect 37660 42690 37716 42702
rect 37772 43652 37828 43662
rect 37772 42642 37828 43596
rect 37884 43650 37940 44156
rect 37996 43762 38052 44828
rect 38108 44772 38164 45054
rect 38108 44324 38164 44716
rect 38108 44258 38164 44268
rect 37996 43710 37998 43762
rect 38050 43710 38052 43762
rect 37996 43698 38052 43710
rect 37884 43598 37886 43650
rect 37938 43598 37940 43650
rect 37884 42756 37940 43598
rect 38108 43538 38164 43550
rect 38108 43486 38110 43538
rect 38162 43486 38164 43538
rect 38108 43204 38164 43486
rect 38108 43138 38164 43148
rect 37884 42690 37940 42700
rect 37772 42590 37774 42642
rect 37826 42590 37828 42642
rect 37772 42578 37828 42590
rect 36988 41188 37044 41356
rect 37772 41972 37828 41982
rect 37772 41300 37828 41916
rect 38108 41412 38164 41422
rect 38108 41318 38164 41356
rect 37772 41234 37828 41244
rect 36876 41132 37044 41188
rect 37884 41188 37940 41198
rect 36540 40964 36596 40974
rect 36540 40962 36708 40964
rect 36540 40910 36542 40962
rect 36594 40910 36708 40962
rect 36540 40908 36708 40910
rect 36540 40898 36596 40908
rect 36428 39778 36484 39788
rect 36540 40514 36596 40526
rect 36540 40462 36542 40514
rect 36594 40462 36596 40514
rect 36428 38834 36484 38846
rect 36428 38782 36430 38834
rect 36482 38782 36484 38834
rect 36428 38668 36484 38782
rect 36092 37958 36148 37996
rect 36204 38612 36484 38668
rect 35868 37828 35924 37838
rect 36204 37828 36260 38612
rect 35756 37826 36260 37828
rect 35756 37774 35870 37826
rect 35922 37774 36260 37826
rect 35756 37772 36260 37774
rect 35084 34972 35308 35028
rect 35364 34972 35588 35028
rect 35644 36484 35700 36494
rect 35084 34914 35140 34972
rect 35308 34962 35364 34972
rect 35084 34862 35086 34914
rect 35138 34862 35140 34914
rect 35084 34850 35140 34862
rect 35532 34802 35588 34814
rect 35532 34750 35534 34802
rect 35586 34750 35588 34802
rect 35084 34690 35140 34702
rect 35084 34638 35086 34690
rect 35138 34638 35140 34690
rect 35084 33572 35140 34638
rect 35532 34244 35588 34750
rect 35532 34178 35588 34188
rect 35644 34130 35700 36428
rect 35756 36372 35812 37772
rect 35868 37762 35924 37772
rect 36540 37492 36596 40462
rect 36092 37436 36596 37492
rect 35980 37044 36036 37054
rect 36092 37044 36148 37436
rect 36540 37380 36596 37436
rect 36540 37314 36596 37324
rect 36652 39396 36708 40908
rect 36876 40852 36932 41132
rect 37884 41094 37940 41132
rect 37212 41076 37268 41086
rect 37212 40982 37268 41020
rect 36988 40964 37044 40974
rect 36988 40870 37044 40908
rect 37100 40962 37156 40974
rect 37100 40910 37102 40962
rect 37154 40910 37156 40962
rect 36876 40786 36932 40796
rect 36316 37268 36372 37278
rect 35980 37042 36148 37044
rect 35980 36990 35982 37042
rect 36034 36990 36148 37042
rect 35980 36988 36148 36990
rect 36204 37154 36260 37166
rect 36204 37102 36206 37154
rect 36258 37102 36260 37154
rect 35756 36306 35812 36316
rect 35868 36482 35924 36494
rect 35868 36430 35870 36482
rect 35922 36430 35924 36482
rect 35868 35308 35924 36430
rect 35756 35252 35924 35308
rect 35756 34244 35812 35252
rect 35868 34804 35924 34814
rect 35980 34804 36036 36988
rect 36204 36932 36260 37102
rect 36204 36148 36260 36876
rect 36204 35364 36260 36092
rect 36316 35698 36372 37212
rect 36428 37266 36484 37278
rect 36428 37214 36430 37266
rect 36482 37214 36484 37266
rect 36428 36372 36484 37214
rect 36428 36278 36484 36316
rect 36540 37044 36596 37054
rect 36316 35646 36318 35698
rect 36370 35646 36372 35698
rect 36316 35634 36372 35646
rect 36540 35586 36596 36988
rect 36652 36932 36708 39340
rect 36876 40404 36932 40414
rect 36876 38946 36932 40348
rect 37100 39844 37156 40910
rect 37436 40964 37492 40974
rect 37212 40516 37268 40526
rect 37212 40422 37268 40460
rect 37436 40404 37492 40908
rect 37436 40338 37492 40348
rect 36876 38894 36878 38946
rect 36930 38894 36932 38946
rect 36876 38882 36932 38894
rect 36988 39788 37156 39844
rect 36876 37826 36932 37838
rect 36876 37774 36878 37826
rect 36930 37774 36932 37826
rect 36876 37268 36932 37774
rect 36988 37492 37044 39788
rect 37212 39620 37268 39630
rect 37212 39618 37380 39620
rect 37212 39566 37214 39618
rect 37266 39566 37380 39618
rect 37212 39564 37380 39566
rect 37212 39554 37268 39564
rect 37324 38612 37380 39564
rect 37884 39506 37940 39518
rect 37884 39454 37886 39506
rect 37938 39454 37940 39506
rect 37212 37938 37268 37950
rect 37212 37886 37214 37938
rect 37266 37886 37268 37938
rect 37100 37828 37156 37838
rect 37100 37734 37156 37772
rect 36988 37426 37044 37436
rect 36876 37202 36932 37212
rect 36652 36866 36708 36876
rect 36876 37044 36932 37054
rect 36652 36260 36708 36270
rect 36652 35698 36708 36204
rect 36652 35646 36654 35698
rect 36706 35646 36708 35698
rect 36652 35634 36708 35646
rect 36540 35534 36542 35586
rect 36594 35534 36596 35586
rect 36204 35308 36372 35364
rect 35868 34802 36036 34804
rect 35868 34750 35870 34802
rect 35922 34750 36036 34802
rect 35868 34748 36036 34750
rect 36204 35140 36260 35150
rect 35868 34738 35924 34748
rect 36092 34692 36148 34702
rect 35980 34636 36092 34692
rect 35868 34244 35924 34254
rect 35756 34188 35868 34244
rect 35868 34178 35924 34188
rect 35980 34242 36036 34636
rect 36092 34626 36148 34636
rect 36204 34354 36260 35084
rect 36204 34302 36206 34354
rect 36258 34302 36260 34354
rect 36204 34290 36260 34302
rect 35980 34190 35982 34242
rect 36034 34190 36036 34242
rect 35980 34178 36036 34190
rect 36092 34244 36148 34254
rect 35644 34078 35646 34130
rect 35698 34078 35700 34130
rect 35644 34066 35700 34078
rect 35308 33908 35364 33918
rect 35308 33906 35588 33908
rect 35308 33854 35310 33906
rect 35362 33854 35588 33906
rect 35308 33852 35588 33854
rect 35308 33842 35364 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35084 33516 35252 33572
rect 35084 33346 35140 33358
rect 35084 33294 35086 33346
rect 35138 33294 35140 33346
rect 35084 32900 35140 33294
rect 35084 32834 35140 32844
rect 35196 32340 35252 33516
rect 35420 33348 35476 33358
rect 35420 33254 35476 33292
rect 35532 32900 35588 33852
rect 36092 33348 36148 34188
rect 36316 34132 36372 35308
rect 36540 35308 36596 35534
rect 36540 35252 36820 35308
rect 36316 34038 36372 34076
rect 36540 34468 36596 34478
rect 35980 33292 36148 33348
rect 36204 33458 36260 33470
rect 36204 33406 36206 33458
rect 36258 33406 36260 33458
rect 35532 32834 35588 32844
rect 35868 33234 35924 33246
rect 35868 33182 35870 33234
rect 35922 33182 35924 33234
rect 35084 32284 35252 32340
rect 34972 31892 35028 31902
rect 34972 31798 35028 31836
rect 34748 31778 34804 31790
rect 34748 31726 34750 31778
rect 34802 31726 34804 31778
rect 34748 31556 34804 31726
rect 34748 31490 34804 31500
rect 33516 30146 33572 30156
rect 33964 31052 34692 31108
rect 32060 30034 32116 30044
rect 33852 30100 33908 30110
rect 31948 29922 32004 29932
rect 33180 29986 33236 29998
rect 33180 29934 33182 29986
rect 33234 29934 33236 29986
rect 31948 29652 32004 29662
rect 31836 29650 32004 29652
rect 31836 29598 31950 29650
rect 32002 29598 32004 29650
rect 31836 29596 32004 29598
rect 31948 29586 32004 29596
rect 32396 29652 32452 29662
rect 32396 29558 32452 29596
rect 33180 29652 33236 29934
rect 33404 29988 33460 29998
rect 33628 29988 33684 29998
rect 33404 29986 33572 29988
rect 33404 29934 33406 29986
rect 33458 29934 33572 29986
rect 33404 29932 33572 29934
rect 33404 29922 33460 29932
rect 33180 29586 33236 29596
rect 33404 29650 33460 29662
rect 33404 29598 33406 29650
rect 33458 29598 33460 29650
rect 31276 29540 31332 29550
rect 31276 29446 31332 29484
rect 33068 29540 33124 29550
rect 31164 29374 31166 29426
rect 31218 29374 31220 29426
rect 31052 28868 31108 28878
rect 31052 28774 31108 28812
rect 31164 28644 31220 29374
rect 32508 29426 32564 29438
rect 32508 29374 32510 29426
rect 32562 29374 32564 29426
rect 32508 28756 32564 29374
rect 33068 28980 33124 29484
rect 33292 29538 33348 29550
rect 33292 29486 33294 29538
rect 33346 29486 33348 29538
rect 33180 29426 33236 29438
rect 33180 29374 33182 29426
rect 33234 29374 33236 29426
rect 33180 29204 33236 29374
rect 33180 29138 33236 29148
rect 33068 28924 33236 28980
rect 32508 28690 32564 28700
rect 32620 28868 32676 28878
rect 31164 28550 31220 28588
rect 31388 28644 31444 28654
rect 31164 28420 31220 28430
rect 31164 28082 31220 28364
rect 31164 28030 31166 28082
rect 31218 28030 31220 28082
rect 31164 27188 31220 28030
rect 31388 28082 31444 28588
rect 31724 28530 31780 28542
rect 32620 28532 32676 28812
rect 33068 28754 33124 28766
rect 33068 28702 33070 28754
rect 33122 28702 33124 28754
rect 31724 28478 31726 28530
rect 31778 28478 31780 28530
rect 31388 28030 31390 28082
rect 31442 28030 31444 28082
rect 31276 27748 31332 27758
rect 31276 27654 31332 27692
rect 30828 25396 30884 26796
rect 30828 25172 30884 25340
rect 30828 25106 30884 25116
rect 30940 27186 31220 27188
rect 30940 27134 31166 27186
rect 31218 27134 31220 27186
rect 30940 27132 31220 27134
rect 30940 24948 30996 27132
rect 31164 27122 31220 27132
rect 31388 27074 31444 28030
rect 31500 28308 31556 28318
rect 31500 27636 31556 28252
rect 31500 27570 31556 27580
rect 31612 27858 31668 27870
rect 31612 27806 31614 27858
rect 31666 27806 31668 27858
rect 31612 27412 31668 27806
rect 31612 27346 31668 27356
rect 31724 27860 31780 28478
rect 32508 28476 32676 28532
rect 32956 28642 33012 28654
rect 32956 28590 32958 28642
rect 33010 28590 33012 28642
rect 32396 28420 32452 28430
rect 31388 27022 31390 27074
rect 31442 27022 31444 27074
rect 31388 27010 31444 27022
rect 31500 26962 31556 26974
rect 31500 26910 31502 26962
rect 31554 26910 31556 26962
rect 31164 26292 31220 26302
rect 30156 23884 30772 23940
rect 30828 24892 30996 24948
rect 31052 26236 31164 26292
rect 30828 23940 30884 24892
rect 30940 24722 30996 24734
rect 30940 24670 30942 24722
rect 30994 24670 30996 24722
rect 30940 24610 30996 24670
rect 30940 24558 30942 24610
rect 30994 24558 30996 24610
rect 30940 24546 30996 24558
rect 30828 23884 30996 23940
rect 29820 23660 29988 23716
rect 30044 23716 30100 23726
rect 29596 23154 29652 23166
rect 29596 23102 29598 23154
rect 29650 23102 29652 23154
rect 29596 23044 29652 23102
rect 29596 22978 29652 22988
rect 29708 23156 29764 23166
rect 29316 22876 29540 22932
rect 29260 22838 29316 22876
rect 29148 22418 29204 22428
rect 29372 22482 29428 22494
rect 29372 22430 29374 22482
rect 29426 22430 29428 22482
rect 29372 22372 29428 22430
rect 29372 22306 29428 22316
rect 29708 21810 29764 23100
rect 29820 22596 29876 23660
rect 29932 23380 29988 23390
rect 29932 23286 29988 23324
rect 29932 22596 29988 22606
rect 29820 22540 29932 22596
rect 29932 22530 29988 22540
rect 30044 22372 30100 23660
rect 29708 21758 29710 21810
rect 29762 21758 29764 21810
rect 29708 21746 29764 21758
rect 29820 22370 30100 22372
rect 29820 22318 30046 22370
rect 30098 22318 30100 22370
rect 29820 22316 30100 22318
rect 29820 21588 29876 22316
rect 30044 22306 30100 22316
rect 29372 21532 29876 21588
rect 29260 21476 29316 21486
rect 29260 20804 29316 21420
rect 29372 21026 29428 21532
rect 30044 21476 30100 21486
rect 30044 21382 30100 21420
rect 29372 20974 29374 21026
rect 29426 20974 29428 21026
rect 29372 20962 29428 20974
rect 29932 21364 29988 21374
rect 29932 20914 29988 21308
rect 30156 20916 30212 23884
rect 30380 23714 30436 23726
rect 30380 23662 30382 23714
rect 30434 23662 30436 23714
rect 30268 23380 30324 23390
rect 30268 21700 30324 23324
rect 30380 23156 30436 23662
rect 30604 23716 30660 23726
rect 30604 23622 30660 23660
rect 30716 23714 30772 23726
rect 30716 23662 30718 23714
rect 30770 23662 30772 23714
rect 30380 23090 30436 23100
rect 30492 23604 30548 23614
rect 30492 23044 30548 23548
rect 30492 22370 30548 22988
rect 30492 22318 30494 22370
rect 30546 22318 30548 22370
rect 30492 22306 30548 22318
rect 30716 22148 30772 23662
rect 30828 23716 30884 23726
rect 30828 23622 30884 23660
rect 30716 22082 30772 22092
rect 30940 22036 30996 23884
rect 31052 23380 31108 26236
rect 31164 26198 31220 26236
rect 31388 26180 31444 26190
rect 31388 25730 31444 26124
rect 31388 25678 31390 25730
rect 31442 25678 31444 25730
rect 31388 25666 31444 25678
rect 31276 25172 31332 25182
rect 31164 25116 31276 25172
rect 31164 25060 31220 25116
rect 31276 25106 31332 25116
rect 31164 24610 31220 25004
rect 31500 24948 31556 26910
rect 31724 26514 31780 27804
rect 31724 26462 31726 26514
rect 31778 26462 31780 26514
rect 31724 26450 31780 26462
rect 31948 28308 32004 28318
rect 31948 27858 32004 28252
rect 32396 27970 32452 28364
rect 32508 28082 32564 28476
rect 32956 28308 33012 28590
rect 32956 28242 33012 28252
rect 33068 28084 33124 28702
rect 32508 28030 32510 28082
rect 32562 28030 32564 28082
rect 32508 28018 32564 28030
rect 32844 28082 33124 28084
rect 32844 28030 33070 28082
rect 33122 28030 33124 28082
rect 32844 28028 33124 28030
rect 32396 27918 32398 27970
rect 32450 27918 32452 27970
rect 32396 27906 32452 27918
rect 31948 27806 31950 27858
rect 32002 27806 32004 27858
rect 31948 27188 32004 27806
rect 31164 24558 31166 24610
rect 31218 24558 31220 24610
rect 31164 24546 31220 24558
rect 31276 24892 31556 24948
rect 31052 23314 31108 23324
rect 31276 23044 31332 24892
rect 31836 24836 31892 24846
rect 31388 24724 31444 24734
rect 31724 24724 31780 24734
rect 31388 24630 31444 24668
rect 31500 24722 31780 24724
rect 31500 24670 31726 24722
rect 31778 24670 31780 24722
rect 31500 24668 31780 24670
rect 31388 23714 31444 23726
rect 31388 23662 31390 23714
rect 31442 23662 31444 23714
rect 31388 23604 31444 23662
rect 31388 23538 31444 23548
rect 31164 22988 31332 23044
rect 30828 21980 30996 22036
rect 31052 22820 31108 22830
rect 30828 21924 30884 21980
rect 30268 21606 30324 21644
rect 30604 21868 30884 21924
rect 29932 20862 29934 20914
rect 29986 20862 29988 20914
rect 29932 20850 29988 20862
rect 30044 20860 30212 20916
rect 29260 20802 29540 20804
rect 29260 20750 29262 20802
rect 29314 20750 29540 20802
rect 29260 20748 29540 20750
rect 29260 20738 29316 20748
rect 29372 19908 29428 19918
rect 29036 19794 29092 19806
rect 29036 19742 29038 19794
rect 29090 19742 29092 19794
rect 29036 19012 29092 19742
rect 29372 19346 29428 19852
rect 29372 19294 29374 19346
rect 29426 19294 29428 19346
rect 29372 19282 29428 19294
rect 29484 19236 29540 20748
rect 29820 20690 29876 20702
rect 29820 20638 29822 20690
rect 29874 20638 29876 20690
rect 29820 20244 29876 20638
rect 29820 20178 29876 20188
rect 29708 20130 29764 20142
rect 29708 20078 29710 20130
rect 29762 20078 29764 20130
rect 29596 19236 29652 19246
rect 29484 19234 29652 19236
rect 29484 19182 29598 19234
rect 29650 19182 29652 19234
rect 29484 19180 29652 19182
rect 29596 19170 29652 19180
rect 29036 18946 29092 18956
rect 29708 18788 29764 20078
rect 29820 20020 29876 20030
rect 29820 19926 29876 19964
rect 29708 18722 29764 18732
rect 29820 19460 29876 19470
rect 29484 18452 29540 18462
rect 28924 18396 29428 18452
rect 28700 18338 29092 18340
rect 28700 18286 28702 18338
rect 28754 18286 29092 18338
rect 28700 18284 29092 18286
rect 28700 18274 28756 18284
rect 28476 17574 28532 17612
rect 28252 16566 28308 16604
rect 28924 17108 28980 17118
rect 28924 16884 28980 17052
rect 28028 16370 28084 16380
rect 27916 16156 28308 16212
rect 27356 15986 27412 15998
rect 27356 15934 27358 15986
rect 27410 15934 27412 15986
rect 27356 14756 27412 15934
rect 27692 15988 27748 15998
rect 27916 15988 27972 16156
rect 27692 15986 27972 15988
rect 27692 15934 27694 15986
rect 27746 15934 27972 15986
rect 27692 15932 27972 15934
rect 28028 15986 28084 15998
rect 28028 15934 28030 15986
rect 28082 15934 28084 15986
rect 27692 15922 27748 15932
rect 28028 15876 28084 15934
rect 28028 15810 28084 15820
rect 28140 15874 28196 15886
rect 28140 15822 28142 15874
rect 28194 15822 28196 15874
rect 28140 15540 28196 15822
rect 27580 15484 28196 15540
rect 27356 14690 27412 14700
rect 27468 15314 27524 15326
rect 27468 15262 27470 15314
rect 27522 15262 27524 15314
rect 27356 14420 27412 14430
rect 27468 14420 27524 15262
rect 27412 14364 27524 14420
rect 27356 14354 27412 14364
rect 27244 13906 27300 13916
rect 26460 13858 26628 13860
rect 26460 13806 26462 13858
rect 26514 13806 26628 13858
rect 26460 13804 26628 13806
rect 27580 13858 27636 15484
rect 27916 15316 27972 15326
rect 27692 15202 27748 15214
rect 27692 15150 27694 15202
rect 27746 15150 27748 15202
rect 27692 15092 27748 15150
rect 27692 15026 27748 15036
rect 27580 13806 27582 13858
rect 27634 13806 27636 13858
rect 26460 13794 26516 13804
rect 27580 13794 27636 13806
rect 27804 14644 27860 14654
rect 26236 13694 26238 13746
rect 26290 13694 26292 13746
rect 26236 13682 26292 13694
rect 26908 13746 26964 13758
rect 26908 13694 26910 13746
rect 26962 13694 26964 13746
rect 25900 13234 25956 13244
rect 25676 12898 25732 12908
rect 25900 12962 25956 12974
rect 25900 12910 25902 12962
rect 25954 12910 25956 12962
rect 25788 12738 25844 12750
rect 25788 12686 25790 12738
rect 25842 12686 25844 12738
rect 25676 12180 25732 12190
rect 25676 12086 25732 12124
rect 25788 11844 25844 12686
rect 25900 12740 25956 12910
rect 26348 12740 26404 12750
rect 25900 12738 26404 12740
rect 25900 12686 26350 12738
rect 26402 12686 26404 12738
rect 25900 12684 26404 12686
rect 25900 12404 25956 12414
rect 26124 12404 26180 12414
rect 25956 12348 26068 12404
rect 25900 12338 25956 12348
rect 25788 11778 25844 11788
rect 25900 12178 25956 12190
rect 25900 12126 25902 12178
rect 25954 12126 25956 12178
rect 25900 11508 25956 12126
rect 25788 11452 25956 11508
rect 25676 11396 25732 11406
rect 25676 11302 25732 11340
rect 25340 9214 25342 9266
rect 25394 9214 25396 9266
rect 25340 9202 25396 9214
rect 25452 10108 25620 10164
rect 25676 10610 25732 10622
rect 25676 10558 25678 10610
rect 25730 10558 25732 10610
rect 25676 10500 25732 10558
rect 25452 9268 25508 10108
rect 25564 9828 25620 9838
rect 25676 9828 25732 10444
rect 25564 9826 25732 9828
rect 25564 9774 25566 9826
rect 25618 9774 25732 9826
rect 25564 9772 25732 9774
rect 25564 9762 25620 9772
rect 25564 9268 25620 9278
rect 25452 9266 25620 9268
rect 25452 9214 25566 9266
rect 25618 9214 25620 9266
rect 25452 9212 25620 9214
rect 25564 9202 25620 9212
rect 25228 9102 25230 9154
rect 25282 9102 25284 9154
rect 25228 9090 25284 9102
rect 25116 8194 25172 8204
rect 25676 8036 25732 9772
rect 25788 9716 25844 11452
rect 25900 11282 25956 11294
rect 25900 11230 25902 11282
rect 25954 11230 25956 11282
rect 25900 10836 25956 11230
rect 25900 10770 25956 10780
rect 26012 10612 26068 12348
rect 26124 12290 26180 12348
rect 26124 12238 26126 12290
rect 26178 12238 26180 12290
rect 26124 12226 26180 12238
rect 26236 11956 26292 11966
rect 26236 10836 26292 11900
rect 26348 11172 26404 12684
rect 26908 12740 26964 13694
rect 27804 12852 27860 14588
rect 26908 12674 26964 12684
rect 27132 12850 27860 12852
rect 27132 12798 27806 12850
rect 27858 12798 27860 12850
rect 27132 12796 27860 12798
rect 26348 11078 26404 11116
rect 26460 12628 26516 12638
rect 26348 10836 26404 10846
rect 26236 10834 26404 10836
rect 26236 10782 26350 10834
rect 26402 10782 26404 10834
rect 26236 10780 26404 10782
rect 26348 10770 26404 10780
rect 26460 10722 26516 12572
rect 27132 12402 27188 12796
rect 27804 12786 27860 12796
rect 27356 12628 27412 12638
rect 27132 12350 27134 12402
rect 27186 12350 27188 12402
rect 27132 12338 27188 12350
rect 27244 12572 27356 12628
rect 26796 11956 26852 11966
rect 26572 11396 26628 11406
rect 26572 11302 26628 11340
rect 26796 11394 26852 11900
rect 26796 11342 26798 11394
rect 26850 11342 26852 11394
rect 26796 11330 26852 11342
rect 27020 11844 27076 11854
rect 26684 11170 26740 11182
rect 27020 11172 27076 11788
rect 27244 11284 27300 12572
rect 27356 12562 27412 12572
rect 27468 12516 27524 12526
rect 26684 11118 26686 11170
rect 26738 11118 26740 11170
rect 26460 10670 26462 10722
rect 26514 10670 26516 10722
rect 26460 10658 26516 10670
rect 26572 10724 26628 10734
rect 26012 10610 26404 10612
rect 26012 10558 26014 10610
rect 26066 10558 26404 10610
rect 26012 10556 26404 10558
rect 26012 10546 26068 10556
rect 25900 10388 25956 10398
rect 25956 10332 26180 10388
rect 25900 10322 25956 10332
rect 25788 9650 25844 9660
rect 25900 9826 25956 9838
rect 25900 9774 25902 9826
rect 25954 9774 25956 9826
rect 25900 9268 25956 9774
rect 25900 9202 25956 9212
rect 25900 9042 25956 9054
rect 25900 8990 25902 9042
rect 25954 8990 25956 9042
rect 25900 8820 25956 8990
rect 26124 9042 26180 10332
rect 26236 9940 26292 9950
rect 26236 9846 26292 9884
rect 26124 8990 26126 9042
rect 26178 8990 26180 9042
rect 26124 8978 26180 8990
rect 26348 9266 26404 10556
rect 26572 9716 26628 10668
rect 26684 10612 26740 11118
rect 26684 10546 26740 10556
rect 26796 11116 27076 11172
rect 27132 11282 27300 11284
rect 27132 11230 27246 11282
rect 27298 11230 27300 11282
rect 27132 11228 27300 11230
rect 26796 10052 26852 11116
rect 27020 10724 27076 10734
rect 27020 10610 27076 10668
rect 27020 10558 27022 10610
rect 27074 10558 27076 10610
rect 27020 10546 27076 10558
rect 27132 10164 27188 11228
rect 27244 11218 27300 11228
rect 27356 11732 27412 11742
rect 27356 11394 27412 11676
rect 27356 11342 27358 11394
rect 27410 11342 27412 11394
rect 27356 11060 27412 11342
rect 26796 9986 26852 9996
rect 27020 10108 27188 10164
rect 27244 11004 27412 11060
rect 27020 9828 27076 10108
rect 27020 9772 27188 9828
rect 26348 9214 26350 9266
rect 26402 9214 26404 9266
rect 25900 8754 25956 8764
rect 26236 8930 26292 8942
rect 26236 8878 26238 8930
rect 26290 8878 26292 8930
rect 25228 7980 25732 8036
rect 26124 8036 26180 8046
rect 25228 6692 25284 7980
rect 26124 7942 26180 7980
rect 25676 7588 25732 7598
rect 26236 7588 26292 8878
rect 26348 8596 26404 9214
rect 26348 8530 26404 8540
rect 26460 9660 26628 9716
rect 26796 9716 26852 9726
rect 25676 7586 26292 7588
rect 25676 7534 25678 7586
rect 25730 7534 26292 7586
rect 25676 7532 26292 7534
rect 25676 7522 25732 7532
rect 25116 6636 25284 6692
rect 25564 7364 25620 7374
rect 25004 6580 25060 6590
rect 25004 6486 25060 6524
rect 24892 6402 24948 6412
rect 24780 6132 24836 6142
rect 24780 6038 24836 6076
rect 24780 5684 24836 5694
rect 24780 5682 25060 5684
rect 24780 5630 24782 5682
rect 24834 5630 25060 5682
rect 24780 5628 25060 5630
rect 24780 5618 24836 5628
rect 24668 5236 24724 5246
rect 24668 5142 24724 5180
rect 25004 5234 25060 5628
rect 25116 5346 25172 6636
rect 25340 6578 25396 6590
rect 25340 6526 25342 6578
rect 25394 6526 25396 6578
rect 25228 6466 25284 6478
rect 25228 6414 25230 6466
rect 25282 6414 25284 6466
rect 25228 6020 25284 6414
rect 25228 5954 25284 5964
rect 25340 6244 25396 6526
rect 25116 5294 25118 5346
rect 25170 5294 25172 5346
rect 25116 5282 25172 5294
rect 25004 5182 25006 5234
rect 25058 5182 25060 5234
rect 25004 5170 25060 5182
rect 24668 4564 24724 4574
rect 24556 4508 24668 4564
rect 24108 4498 24164 4508
rect 24220 4470 24276 4508
rect 24668 4470 24724 4508
rect 24108 3668 24164 3678
rect 24780 3668 24836 3678
rect 23996 3666 24836 3668
rect 23996 3614 24110 3666
rect 24162 3614 24782 3666
rect 24834 3614 24836 3666
rect 23996 3612 24836 3614
rect 24108 3602 24164 3612
rect 24780 3602 24836 3612
rect 25228 3668 25284 3678
rect 25340 3668 25396 6188
rect 25452 6468 25508 6478
rect 25452 6130 25508 6412
rect 25564 6244 25620 7308
rect 26460 6914 26516 9660
rect 26796 9268 26852 9660
rect 26796 9156 26852 9212
rect 26908 9156 26964 9166
rect 26796 9154 26964 9156
rect 26796 9102 26910 9154
rect 26962 9102 26964 9154
rect 26796 9100 26964 9102
rect 26908 9090 26964 9100
rect 26572 9044 26628 9054
rect 26572 8950 26628 8988
rect 27132 8428 27188 9772
rect 27244 9266 27300 11004
rect 27356 10836 27412 10846
rect 27356 10722 27412 10780
rect 27356 10670 27358 10722
rect 27410 10670 27412 10722
rect 27356 10276 27412 10670
rect 27356 10210 27412 10220
rect 27244 9214 27246 9266
rect 27298 9214 27300 9266
rect 27244 9202 27300 9214
rect 27020 8372 27188 8428
rect 27020 8260 27076 8372
rect 26908 8204 27076 8260
rect 27132 8258 27188 8270
rect 27132 8206 27134 8258
rect 27186 8206 27188 8258
rect 26572 8036 26628 8046
rect 26628 7980 26852 8036
rect 26572 7970 26628 7980
rect 26460 6862 26462 6914
rect 26514 6862 26516 6914
rect 26460 6850 26516 6862
rect 26572 7812 26628 7822
rect 25676 6580 25732 6590
rect 25676 6486 25732 6524
rect 26012 6578 26068 6590
rect 26012 6526 26014 6578
rect 26066 6526 26068 6578
rect 25564 6178 25620 6188
rect 25452 6078 25454 6130
rect 25506 6078 25508 6130
rect 25452 6066 25508 6078
rect 25900 5684 25956 5694
rect 25676 5346 25732 5358
rect 25676 5294 25678 5346
rect 25730 5294 25732 5346
rect 25676 5234 25732 5294
rect 25676 5182 25678 5234
rect 25730 5182 25732 5234
rect 25676 5170 25732 5182
rect 25900 5348 25956 5628
rect 25452 4564 25508 4574
rect 25452 4470 25508 4508
rect 25900 4562 25956 5292
rect 26012 5124 26068 6526
rect 26348 6580 26404 6590
rect 26348 6130 26404 6524
rect 26572 6468 26628 7756
rect 26348 6078 26350 6130
rect 26402 6078 26404 6130
rect 26348 6066 26404 6078
rect 26460 6412 26628 6468
rect 26796 6914 26852 7980
rect 26796 6862 26798 6914
rect 26850 6862 26852 6914
rect 26796 6580 26852 6862
rect 26012 5058 26068 5068
rect 26124 4900 26180 4910
rect 26124 4806 26180 4844
rect 26460 4900 26516 6412
rect 26684 6244 26740 6254
rect 26572 5236 26628 5246
rect 26684 5236 26740 6188
rect 26796 6020 26852 6524
rect 26796 5954 26852 5964
rect 26796 5348 26852 5358
rect 26908 5348 26964 8204
rect 27132 8148 27188 8206
rect 27356 8260 27412 8270
rect 27356 8166 27412 8204
rect 27020 8092 27132 8148
rect 27020 6916 27076 8092
rect 27132 8082 27188 8092
rect 27468 7924 27524 12460
rect 27916 11788 27972 15260
rect 28140 14530 28196 14542
rect 28140 14478 28142 14530
rect 28194 14478 28196 14530
rect 28140 13972 28196 14478
rect 27804 11732 27972 11788
rect 28028 12068 28084 12078
rect 27692 9042 27748 9054
rect 27692 8990 27694 9042
rect 27746 8990 27748 9042
rect 27692 8932 27748 8990
rect 27692 8866 27748 8876
rect 27692 8036 27748 8046
rect 27692 7942 27748 7980
rect 27020 6850 27076 6860
rect 27132 7868 27524 7924
rect 26796 5346 26964 5348
rect 26796 5294 26798 5346
rect 26850 5294 26964 5346
rect 26796 5292 26964 5294
rect 26796 5282 26852 5292
rect 26572 5234 26684 5236
rect 26572 5182 26574 5234
rect 26626 5182 26684 5234
rect 26572 5180 26684 5182
rect 26572 5170 26628 5180
rect 26684 5170 26740 5180
rect 26460 4834 26516 4844
rect 26684 4900 26740 4910
rect 25900 4510 25902 4562
rect 25954 4510 25956 4562
rect 25900 4498 25956 4510
rect 26684 4562 26740 4844
rect 26684 4510 26686 4562
rect 26738 4510 26740 4562
rect 26684 4498 26740 4510
rect 26908 4564 26964 5292
rect 26908 4498 26964 4508
rect 27020 5236 27076 5246
rect 27020 4562 27076 5180
rect 27132 5234 27188 7868
rect 27804 7700 27860 11732
rect 28028 11618 28084 12012
rect 28028 11566 28030 11618
rect 28082 11566 28084 11618
rect 28028 11554 28084 11566
rect 28140 11284 28196 13916
rect 28252 12404 28308 16156
rect 28364 16100 28420 16110
rect 28364 16006 28420 16044
rect 28476 16098 28532 16110
rect 28476 16046 28478 16098
rect 28530 16046 28532 16098
rect 28364 14532 28420 14542
rect 28364 14438 28420 14476
rect 28476 14306 28532 16046
rect 28812 16100 28868 16110
rect 28700 15428 28756 15438
rect 28700 15334 28756 15372
rect 28476 14254 28478 14306
rect 28530 14254 28532 14306
rect 28476 14242 28532 14254
rect 28588 14530 28644 14542
rect 28588 14478 28590 14530
rect 28642 14478 28644 14530
rect 28588 14308 28644 14478
rect 28588 14242 28644 14252
rect 28252 12310 28308 12348
rect 28700 12628 28756 12638
rect 28140 11218 28196 11228
rect 28252 12180 28308 12190
rect 27916 10724 27972 10734
rect 27972 10668 28084 10724
rect 27916 10658 27972 10668
rect 27692 7644 27804 7700
rect 27468 7250 27524 7262
rect 27468 7198 27470 7250
rect 27522 7198 27524 7250
rect 27132 5182 27134 5234
rect 27186 5182 27188 5234
rect 27132 5170 27188 5182
rect 27244 6692 27300 6702
rect 27244 6356 27300 6636
rect 27468 6580 27524 7198
rect 27692 7028 27748 7644
rect 27804 7634 27860 7644
rect 27916 10276 27972 10286
rect 27916 9716 27972 10220
rect 28028 9938 28084 10668
rect 28252 10498 28308 12124
rect 28700 11956 28756 12572
rect 28700 11890 28756 11900
rect 28364 11620 28420 11630
rect 28364 11526 28420 11564
rect 28588 10948 28644 10958
rect 28588 10610 28644 10892
rect 28588 10558 28590 10610
rect 28642 10558 28644 10610
rect 28588 10546 28644 10558
rect 28252 10446 28254 10498
rect 28306 10446 28308 10498
rect 28252 10434 28308 10446
rect 28028 9886 28030 9938
rect 28082 9886 28084 9938
rect 28028 9874 28084 9886
rect 28588 10052 28644 10062
rect 28140 9826 28196 9838
rect 28140 9774 28142 9826
rect 28194 9774 28196 9826
rect 28140 9716 28196 9774
rect 27916 9660 28196 9716
rect 28252 9828 28308 9838
rect 27804 7476 27860 7486
rect 27916 7476 27972 9660
rect 28028 9156 28084 9166
rect 28028 9042 28084 9100
rect 28028 8990 28030 9042
rect 28082 8990 28084 9042
rect 28028 8596 28084 8990
rect 28140 8932 28196 8942
rect 28140 8838 28196 8876
rect 28028 8530 28084 8540
rect 28252 8484 28308 9772
rect 28364 9716 28420 9726
rect 28364 9044 28420 9660
rect 28588 9266 28644 9996
rect 28812 9716 28868 16044
rect 28924 15314 28980 16828
rect 29036 16882 29092 18284
rect 29148 18228 29204 18238
rect 29148 17666 29204 18172
rect 29148 17614 29150 17666
rect 29202 17614 29204 17666
rect 29148 17602 29204 17614
rect 29260 18116 29316 18126
rect 29036 16830 29038 16882
rect 29090 16830 29092 16882
rect 29036 16818 29092 16830
rect 29148 17444 29204 17454
rect 29148 16098 29204 17388
rect 29148 16046 29150 16098
rect 29202 16046 29204 16098
rect 29148 16034 29204 16046
rect 29260 15986 29316 18060
rect 29260 15934 29262 15986
rect 29314 15934 29316 15986
rect 29260 15922 29316 15934
rect 28924 15262 28926 15314
rect 28978 15262 28980 15314
rect 28924 15250 28980 15262
rect 29148 15876 29204 15886
rect 29148 15148 29204 15820
rect 28924 15092 29204 15148
rect 29372 15148 29428 18396
rect 29484 16098 29540 18396
rect 29596 18116 29652 18126
rect 29596 17778 29652 18060
rect 29596 17726 29598 17778
rect 29650 17726 29652 17778
rect 29596 17714 29652 17726
rect 29708 17892 29764 17902
rect 29708 17556 29764 17836
rect 29484 16046 29486 16098
rect 29538 16046 29540 16098
rect 29484 16034 29540 16046
rect 29596 17500 29764 17556
rect 29596 16098 29652 17500
rect 29708 16660 29764 16670
rect 29708 16566 29764 16604
rect 29596 16046 29598 16098
rect 29650 16046 29652 16098
rect 29596 16034 29652 16046
rect 29708 16436 29764 16446
rect 29708 15988 29764 16380
rect 29820 16100 29876 19404
rect 29932 16884 29988 16894
rect 29932 16790 29988 16828
rect 29932 16100 29988 16110
rect 29820 16098 29988 16100
rect 29820 16046 29934 16098
rect 29986 16046 29988 16098
rect 29820 16044 29988 16046
rect 29932 16034 29988 16044
rect 29708 15932 29876 15988
rect 29708 15540 29764 15550
rect 29372 15092 29540 15148
rect 28924 12740 28980 15092
rect 29260 14644 29316 14654
rect 29260 14550 29316 14588
rect 29372 14532 29428 14542
rect 29148 14308 29204 14318
rect 28924 12178 28980 12684
rect 28924 12126 28926 12178
rect 28978 12126 28980 12178
rect 28924 12114 28980 12126
rect 29036 14306 29204 14308
rect 29036 14254 29150 14306
rect 29202 14254 29204 14306
rect 29036 14252 29204 14254
rect 29036 12516 29092 14252
rect 29148 14242 29204 14252
rect 29260 13076 29316 13086
rect 29372 13076 29428 14476
rect 29260 13074 29428 13076
rect 29260 13022 29262 13074
rect 29314 13022 29428 13074
rect 29260 13020 29428 13022
rect 29260 13010 29316 13020
rect 29148 12738 29204 12750
rect 29148 12686 29150 12738
rect 29202 12686 29204 12738
rect 29148 12628 29204 12686
rect 29148 12562 29204 12572
rect 29372 12740 29428 12750
rect 29036 11844 29092 12460
rect 29036 11778 29092 11788
rect 29148 12404 29204 12414
rect 29148 11394 29204 12348
rect 29260 12290 29316 12302
rect 29260 12238 29262 12290
rect 29314 12238 29316 12290
rect 29260 11732 29316 12238
rect 29260 11666 29316 11676
rect 29148 11342 29150 11394
rect 29202 11342 29204 11394
rect 29148 11330 29204 11342
rect 29372 11396 29428 12684
rect 29372 11330 29428 11340
rect 29372 9828 29428 9838
rect 29372 9734 29428 9772
rect 28812 9660 29092 9716
rect 28588 9214 28590 9266
rect 28642 9214 28644 9266
rect 28588 9202 28644 9214
rect 28812 9268 28868 9278
rect 28812 9174 28868 9212
rect 28700 9044 28756 9054
rect 28364 9042 28644 9044
rect 28364 8990 28366 9042
rect 28418 8990 28644 9042
rect 28364 8988 28644 8990
rect 28364 8978 28420 8988
rect 28588 8708 28644 8988
rect 28700 8950 28756 8988
rect 28588 8652 28868 8708
rect 28028 7700 28084 7710
rect 28252 7700 28308 8428
rect 28588 8258 28644 8270
rect 28588 8206 28590 8258
rect 28642 8206 28644 8258
rect 28588 8148 28644 8206
rect 28700 8148 28756 8158
rect 28588 8092 28700 8148
rect 28700 8082 28756 8092
rect 28028 7698 28308 7700
rect 28028 7646 28030 7698
rect 28082 7646 28308 7698
rect 28028 7644 28308 7646
rect 28364 8034 28420 8046
rect 28364 7982 28366 8034
rect 28418 7982 28420 8034
rect 28364 7700 28420 7982
rect 28476 8036 28532 8046
rect 28476 7942 28532 7980
rect 28028 7634 28084 7644
rect 28364 7634 28420 7644
rect 28476 7588 28532 7598
rect 28476 7494 28532 7532
rect 28812 7586 28868 8652
rect 28812 7534 28814 7586
rect 28866 7534 28868 7586
rect 28812 7522 28868 7534
rect 27804 7474 27972 7476
rect 27804 7422 27806 7474
rect 27858 7422 27972 7474
rect 27804 7420 27972 7422
rect 27804 7410 27860 7420
rect 28924 7364 28980 7374
rect 27692 6962 27748 6972
rect 28252 7362 28980 7364
rect 28252 7310 28926 7362
rect 28978 7310 28980 7362
rect 28252 7308 28980 7310
rect 28140 6692 28196 6702
rect 27580 6580 27636 6590
rect 27468 6578 27636 6580
rect 27468 6526 27582 6578
rect 27634 6526 27636 6578
rect 27468 6524 27636 6526
rect 27580 6468 27636 6524
rect 27580 6402 27636 6412
rect 28140 6356 28196 6636
rect 28252 6578 28308 7308
rect 28924 7298 28980 7308
rect 28476 7140 28532 7150
rect 28476 7028 28532 7084
rect 28476 6972 28644 7028
rect 28252 6526 28254 6578
rect 28306 6526 28308 6578
rect 28252 6514 28308 6526
rect 28476 6802 28532 6814
rect 28476 6750 28478 6802
rect 28530 6750 28532 6802
rect 28476 6580 28532 6750
rect 28476 6514 28532 6524
rect 28364 6466 28420 6478
rect 28364 6414 28366 6466
rect 28418 6414 28420 6466
rect 28140 6300 28308 6356
rect 27244 5012 27300 6300
rect 28140 6020 28196 6030
rect 28140 5926 28196 5964
rect 27468 5908 27524 5918
rect 28028 5908 28084 5918
rect 27468 5906 28084 5908
rect 27468 5854 27470 5906
rect 27522 5854 28030 5906
rect 28082 5854 28084 5906
rect 27468 5852 28084 5854
rect 27468 5842 27524 5852
rect 27692 5122 27748 5852
rect 28028 5842 28084 5852
rect 27692 5070 27694 5122
rect 27746 5070 27748 5122
rect 27692 5058 27748 5070
rect 28028 5124 28084 5134
rect 27356 5012 27412 5022
rect 27244 5010 27412 5012
rect 27244 4958 27358 5010
rect 27410 4958 27412 5010
rect 27244 4956 27412 4958
rect 27356 4946 27412 4956
rect 28028 5010 28084 5068
rect 28252 5122 28308 6300
rect 28364 5684 28420 6414
rect 28588 6356 28644 6972
rect 28364 5618 28420 5628
rect 28476 6300 28644 6356
rect 28812 6468 28868 6478
rect 28476 6132 28532 6300
rect 28252 5070 28254 5122
rect 28306 5070 28308 5122
rect 28252 5058 28308 5070
rect 28028 4958 28030 5010
rect 28082 4958 28084 5010
rect 28028 4946 28084 4958
rect 27020 4510 27022 4562
rect 27074 4510 27076 4562
rect 27020 4498 27076 4510
rect 27468 4676 27524 4686
rect 27468 3892 27524 4620
rect 27916 4564 27972 4574
rect 27972 4508 28084 4564
rect 27916 4498 27972 4508
rect 27916 4340 27972 4350
rect 27916 4246 27972 4284
rect 27580 4226 27636 4238
rect 27580 4174 27582 4226
rect 27634 4174 27636 4226
rect 27580 4114 27636 4174
rect 27580 4062 27582 4114
rect 27634 4062 27636 4114
rect 27580 4050 27636 4062
rect 27020 3780 27076 3790
rect 25228 3666 25396 3668
rect 25228 3614 25230 3666
rect 25282 3614 25396 3666
rect 25228 3612 25396 3614
rect 26124 3668 26180 3678
rect 25228 3602 25284 3612
rect 26124 3574 26180 3612
rect 25676 3556 25732 3566
rect 25676 3462 25732 3500
rect 23100 3332 23492 3388
rect 26572 3444 26628 3482
rect 26572 3378 26628 3388
rect 27020 3442 27076 3724
rect 27468 3666 27524 3836
rect 27468 3614 27470 3666
rect 27522 3614 27524 3666
rect 27468 3602 27524 3614
rect 27916 3668 27972 3678
rect 28028 3668 28084 4508
rect 28476 4562 28532 6076
rect 28812 5906 28868 6412
rect 28812 5854 28814 5906
rect 28866 5854 28868 5906
rect 28812 5842 28868 5854
rect 28476 4510 28478 4562
rect 28530 4510 28532 4562
rect 28476 4114 28532 4510
rect 28924 4564 28980 4574
rect 29036 4564 29092 9660
rect 29260 9268 29316 9278
rect 29260 9042 29316 9212
rect 29484 9154 29540 15092
rect 29596 14756 29652 14766
rect 29596 14530 29652 14700
rect 29596 14478 29598 14530
rect 29650 14478 29652 14530
rect 29596 14466 29652 14478
rect 29596 14308 29652 14318
rect 29596 14214 29652 14252
rect 29708 13634 29764 15484
rect 29708 13582 29710 13634
rect 29762 13582 29764 13634
rect 29708 13570 29764 13582
rect 29708 12962 29764 12974
rect 29708 12910 29710 12962
rect 29762 12910 29764 12962
rect 29708 12852 29764 12910
rect 29708 12786 29764 12796
rect 29596 12292 29652 12302
rect 29596 11506 29652 12236
rect 29596 11454 29598 11506
rect 29650 11454 29652 11506
rect 29596 11442 29652 11454
rect 29484 9102 29486 9154
rect 29538 9102 29540 9154
rect 29484 9090 29540 9102
rect 29596 11284 29652 11294
rect 29260 8990 29262 9042
rect 29314 8990 29316 9042
rect 29260 8978 29316 8990
rect 29260 8596 29316 8606
rect 29148 8258 29204 8270
rect 29148 8206 29150 8258
rect 29202 8206 29204 8258
rect 29148 7812 29204 8206
rect 29148 7746 29204 7756
rect 29148 7588 29204 7598
rect 29260 7588 29316 8540
rect 29148 7586 29316 7588
rect 29148 7534 29150 7586
rect 29202 7534 29316 7586
rect 29148 7532 29316 7534
rect 29148 7522 29204 7532
rect 29372 7476 29428 7486
rect 29372 7382 29428 7420
rect 29596 7252 29652 11228
rect 29820 10388 29876 15932
rect 30044 15876 30100 20860
rect 30156 20690 30212 20702
rect 30156 20638 30158 20690
rect 30210 20638 30212 20690
rect 30156 20356 30212 20638
rect 30380 20692 30436 20702
rect 30380 20598 30436 20636
rect 30156 20290 30212 20300
rect 30604 20580 30660 21868
rect 30940 21812 30996 21822
rect 30828 21756 30940 21812
rect 30492 20132 30548 20142
rect 30492 20038 30548 20076
rect 30380 20018 30436 20030
rect 30380 19966 30382 20018
rect 30434 19966 30436 20018
rect 30380 19684 30436 19966
rect 30156 19348 30212 19358
rect 30156 19254 30212 19292
rect 30380 18004 30436 19628
rect 30492 19124 30548 19134
rect 30492 18676 30548 19068
rect 30492 18450 30548 18620
rect 30492 18398 30494 18450
rect 30546 18398 30548 18450
rect 30492 18386 30548 18398
rect 30380 17948 30548 18004
rect 30380 17780 30436 17790
rect 30380 17686 30436 17724
rect 30268 17666 30324 17678
rect 30268 17614 30270 17666
rect 30322 17614 30324 17666
rect 30156 16772 30212 16782
rect 30156 15986 30212 16716
rect 30268 16322 30324 17614
rect 30380 17108 30436 17118
rect 30380 17014 30436 17052
rect 30268 16270 30270 16322
rect 30322 16270 30324 16322
rect 30268 16258 30324 16270
rect 30156 15934 30158 15986
rect 30210 15934 30212 15986
rect 30156 15922 30212 15934
rect 30044 15810 30100 15820
rect 30492 15316 30548 17948
rect 30604 16212 30660 20524
rect 30716 20690 30772 20702
rect 30716 20638 30718 20690
rect 30770 20638 30772 20690
rect 30716 20468 30772 20638
rect 30716 20402 30772 20412
rect 30716 20132 30772 20142
rect 30828 20132 30884 21756
rect 30940 21746 30996 21756
rect 31052 21810 31108 22764
rect 31052 21758 31054 21810
rect 31106 21758 31108 21810
rect 31052 21746 31108 21758
rect 31164 21588 31220 22988
rect 31500 22820 31556 24668
rect 31724 24658 31780 24668
rect 31836 24052 31892 24780
rect 31948 24834 32004 27132
rect 32508 27412 32564 27422
rect 32172 27074 32228 27086
rect 32172 27022 32174 27074
rect 32226 27022 32228 27074
rect 32172 26290 32228 27022
rect 32508 27074 32564 27356
rect 32508 27022 32510 27074
rect 32562 27022 32564 27074
rect 32508 27010 32564 27022
rect 32172 26238 32174 26290
rect 32226 26238 32228 26290
rect 32172 26180 32228 26238
rect 32172 26114 32228 26124
rect 32396 26178 32452 26190
rect 32396 26126 32398 26178
rect 32450 26126 32452 26178
rect 32396 25956 32452 26126
rect 32396 25506 32452 25900
rect 32396 25454 32398 25506
rect 32450 25454 32452 25506
rect 32396 25442 32452 25454
rect 32844 25508 32900 28028
rect 33068 28018 33124 28028
rect 33180 28082 33236 28924
rect 33292 28644 33348 29486
rect 33292 28578 33348 28588
rect 33180 28030 33182 28082
rect 33234 28030 33236 28082
rect 33180 28018 33236 28030
rect 33292 27860 33348 27870
rect 32956 27858 33348 27860
rect 32956 27806 33294 27858
rect 33346 27806 33348 27858
rect 32956 27804 33348 27806
rect 32956 27074 33012 27804
rect 33292 27794 33348 27804
rect 33404 27412 33460 29598
rect 33404 27346 33460 27356
rect 33516 28084 33572 29932
rect 33628 29986 33796 29988
rect 33628 29934 33630 29986
rect 33682 29934 33796 29986
rect 33628 29932 33796 29934
rect 33628 29922 33684 29932
rect 33404 27188 33460 27198
rect 33404 27094 33460 27132
rect 32956 27022 32958 27074
rect 33010 27022 33012 27074
rect 32956 25956 33012 27022
rect 33516 26908 33572 28028
rect 33740 29876 33796 29932
rect 33628 27860 33684 27870
rect 33628 27766 33684 27804
rect 33740 27748 33796 29820
rect 33852 29538 33908 30044
rect 33852 29486 33854 29538
rect 33906 29486 33908 29538
rect 33852 29474 33908 29486
rect 33852 28756 33908 28766
rect 33852 28082 33908 28700
rect 33852 28030 33854 28082
rect 33906 28030 33908 28082
rect 33852 28018 33908 28030
rect 33964 27860 34020 31052
rect 34188 30982 34244 30994
rect 34188 30930 34190 30982
rect 34242 30930 34244 30982
rect 34188 30884 34244 30930
rect 34972 30884 35028 30894
rect 34188 30818 34244 30828
rect 34524 30882 35028 30884
rect 34524 30830 34974 30882
rect 35026 30830 35028 30882
rect 34524 30828 35028 30830
rect 34188 30660 34244 30670
rect 34188 30210 34244 30604
rect 34524 30548 34580 30828
rect 34972 30818 35028 30828
rect 34300 30492 34580 30548
rect 34300 30322 34356 30492
rect 35084 30436 35140 32284
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35532 31780 35588 31790
rect 35532 31686 35588 31724
rect 35756 31778 35812 31790
rect 35756 31726 35758 31778
rect 35810 31726 35812 31778
rect 35756 31556 35812 31726
rect 35756 31490 35812 31500
rect 35868 31554 35924 33182
rect 35980 32340 36036 33292
rect 36092 33122 36148 33134
rect 36092 33070 36094 33122
rect 36146 33070 36148 33122
rect 36092 32788 36148 33070
rect 36092 32722 36148 32732
rect 36204 32674 36260 33406
rect 36204 32622 36206 32674
rect 36258 32622 36260 32674
rect 36204 32610 36260 32622
rect 35980 32274 36036 32284
rect 35980 31892 36036 31902
rect 35980 31778 36036 31836
rect 35980 31726 35982 31778
rect 36034 31726 36036 31778
rect 35980 31714 36036 31726
rect 36428 31890 36484 31902
rect 36428 31838 36430 31890
rect 36482 31838 36484 31890
rect 36428 31780 36484 31838
rect 36428 31714 36484 31724
rect 36316 31668 36372 31678
rect 36316 31574 36372 31612
rect 35868 31502 35870 31554
rect 35922 31502 35924 31554
rect 35868 31490 35924 31502
rect 36540 30996 36596 34412
rect 36652 34242 36708 34254
rect 36652 34190 36654 34242
rect 36706 34190 36708 34242
rect 36652 33012 36708 34190
rect 36652 32946 36708 32956
rect 36540 30930 36596 30940
rect 35644 30772 35700 30782
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34300 30270 34302 30322
rect 34354 30270 34356 30322
rect 34300 30258 34356 30270
rect 34524 30380 35140 30436
rect 34188 30158 34190 30210
rect 34242 30158 34244 30210
rect 34188 30146 34244 30158
rect 34412 30212 34468 30222
rect 34412 30118 34468 30156
rect 34524 29988 34580 30380
rect 34748 30212 34804 30222
rect 34972 30212 35028 30222
rect 34748 30210 35028 30212
rect 34748 30158 34750 30210
rect 34802 30158 34974 30210
rect 35026 30158 35028 30210
rect 34748 30156 35028 30158
rect 34748 30146 34804 30156
rect 34972 30146 35028 30156
rect 35644 30210 35700 30716
rect 36092 30212 36148 30222
rect 35644 30158 35646 30210
rect 35698 30158 35700 30210
rect 34412 29932 34580 29988
rect 34972 29988 35028 29998
rect 34300 28308 34356 28318
rect 34076 28084 34132 28094
rect 34076 27990 34132 28028
rect 33740 26908 33796 27692
rect 32956 25890 33012 25900
rect 33068 26852 33124 26862
rect 33068 26402 33124 26796
rect 33180 26852 33572 26908
rect 33628 26852 33796 26908
rect 33852 27804 34020 27860
rect 34188 27858 34244 27870
rect 34188 27806 34190 27858
rect 34242 27806 34244 27858
rect 33180 26514 33236 26852
rect 33180 26462 33182 26514
rect 33234 26462 33236 26514
rect 33180 26450 33236 26462
rect 33068 26350 33070 26402
rect 33122 26350 33124 26402
rect 33068 25732 33124 26350
rect 33628 26178 33684 26852
rect 33628 26126 33630 26178
rect 33682 26126 33684 26178
rect 33068 25676 33348 25732
rect 33068 25508 33124 25518
rect 32844 25506 33236 25508
rect 32844 25454 33070 25506
rect 33122 25454 33236 25506
rect 32844 25452 33236 25454
rect 33068 25442 33124 25452
rect 32732 25172 32788 25182
rect 31948 24782 31950 24834
rect 32002 24782 32004 24834
rect 31948 24612 32004 24782
rect 32060 24836 32116 24846
rect 32060 24742 32116 24780
rect 31948 24546 32004 24556
rect 32172 24722 32228 24734
rect 32172 24670 32174 24722
rect 32226 24670 32228 24722
rect 32172 24164 32228 24670
rect 32172 24098 32228 24108
rect 31612 23996 31892 24052
rect 31612 23940 31668 23996
rect 32060 23940 32116 23950
rect 31612 23846 31668 23884
rect 31948 23938 32116 23940
rect 31948 23886 32062 23938
rect 32114 23886 32116 23938
rect 31948 23884 32116 23886
rect 31836 23826 31892 23838
rect 31836 23774 31838 23826
rect 31890 23774 31892 23826
rect 31836 23492 31892 23774
rect 31500 22754 31556 22764
rect 31612 23436 31892 23492
rect 31052 20804 31108 20814
rect 31164 20804 31220 21532
rect 31052 20802 31220 20804
rect 31052 20750 31054 20802
rect 31106 20750 31220 20802
rect 31052 20748 31220 20750
rect 31276 22708 31332 22718
rect 31052 20738 31108 20748
rect 31276 20690 31332 22652
rect 31500 22372 31556 22382
rect 31500 22278 31556 22316
rect 31612 21698 31668 23436
rect 31612 21646 31614 21698
rect 31666 21646 31668 21698
rect 31388 21364 31444 21374
rect 31388 21270 31444 21308
rect 31612 21140 31668 21646
rect 31612 21074 31668 21084
rect 31724 23266 31780 23278
rect 31724 23214 31726 23266
rect 31778 23214 31780 23266
rect 31724 20914 31780 23214
rect 31836 22258 31892 22270
rect 31836 22206 31838 22258
rect 31890 22206 31892 22258
rect 31836 21812 31892 22206
rect 31948 22036 32004 23884
rect 32060 23874 32116 23884
rect 32172 23938 32228 23950
rect 32172 23886 32174 23938
rect 32226 23886 32228 23938
rect 32172 22708 32228 23886
rect 32172 22642 32228 22652
rect 32284 23940 32340 23950
rect 32060 22596 32116 22606
rect 32060 22370 32116 22540
rect 32060 22318 32062 22370
rect 32114 22318 32116 22370
rect 32060 22306 32116 22318
rect 32172 22258 32228 22270
rect 32172 22206 32174 22258
rect 32226 22206 32228 22258
rect 32060 22036 32116 22046
rect 31948 21980 32060 22036
rect 31836 21746 31892 21756
rect 32060 21476 32116 21980
rect 32172 21924 32228 22206
rect 32172 21858 32228 21868
rect 32284 22260 32340 23884
rect 32396 23716 32452 23726
rect 32396 23714 32676 23716
rect 32396 23662 32398 23714
rect 32450 23662 32676 23714
rect 32396 23660 32676 23662
rect 32396 23650 32452 23660
rect 32620 22594 32676 23660
rect 32620 22542 32622 22594
rect 32674 22542 32676 22594
rect 32620 22530 32676 22542
rect 32732 22484 32788 25116
rect 33180 24162 33236 25452
rect 33180 24110 33182 24162
rect 33234 24110 33236 24162
rect 33180 24098 33236 24110
rect 33180 23268 33236 23278
rect 33180 23174 33236 23212
rect 33068 22930 33124 22942
rect 33068 22878 33070 22930
rect 33122 22878 33124 22930
rect 33068 22708 33124 22878
rect 33068 22642 33124 22652
rect 32732 22418 32788 22428
rect 33292 22484 33348 25676
rect 33516 25394 33572 25406
rect 33516 25342 33518 25394
rect 33570 25342 33572 25394
rect 33404 24836 33460 24846
rect 33404 24742 33460 24780
rect 33516 24500 33572 25342
rect 33516 24434 33572 24444
rect 33516 23940 33572 23950
rect 33516 23846 33572 23884
rect 33292 22418 33348 22428
rect 33404 23604 33460 23614
rect 33628 23604 33684 26126
rect 33460 23548 33684 23604
rect 32172 21700 32228 21710
rect 32284 21700 32340 22204
rect 32396 22370 32452 22382
rect 32396 22318 32398 22370
rect 32450 22318 32452 22370
rect 32396 21812 32452 22318
rect 33068 22260 33124 22270
rect 33292 22260 33348 22270
rect 33068 22166 33124 22204
rect 33180 22258 33348 22260
rect 33180 22206 33294 22258
rect 33346 22206 33348 22258
rect 33180 22204 33348 22206
rect 32396 21746 32452 21756
rect 32732 21924 32788 21934
rect 32172 21698 32340 21700
rect 32172 21646 32174 21698
rect 32226 21646 32340 21698
rect 32172 21644 32340 21646
rect 32732 21700 32788 21868
rect 32732 21644 33012 21700
rect 32172 21634 32228 21644
rect 31724 20862 31726 20914
rect 31778 20862 31780 20914
rect 31724 20850 31780 20862
rect 31836 21420 32116 21476
rect 31276 20638 31278 20690
rect 31330 20638 31332 20690
rect 31276 20626 31332 20638
rect 31612 20802 31668 20814
rect 31612 20750 31614 20802
rect 31666 20750 31668 20802
rect 30940 20580 30996 20590
rect 30940 20486 30996 20524
rect 31500 20580 31556 20590
rect 31612 20580 31668 20750
rect 31556 20524 31668 20580
rect 31500 20514 31556 20524
rect 31052 20356 31108 20366
rect 30716 20130 30884 20132
rect 30716 20078 30718 20130
rect 30770 20078 30884 20130
rect 30716 20076 30884 20078
rect 30940 20244 30996 20254
rect 30716 20066 30772 20076
rect 30940 20020 30996 20188
rect 30828 20018 30996 20020
rect 30828 19966 30942 20018
rect 30994 19966 30996 20018
rect 30828 19964 30996 19966
rect 30716 18452 30772 18462
rect 30716 18358 30772 18396
rect 30828 18228 30884 19964
rect 30940 19954 30996 19964
rect 31052 20130 31108 20300
rect 31052 20078 31054 20130
rect 31106 20078 31108 20130
rect 30716 18172 30884 18228
rect 30940 18452 30996 18462
rect 30716 17778 30772 18172
rect 30716 17726 30718 17778
rect 30770 17726 30772 17778
rect 30716 16660 30772 17726
rect 30828 17668 30884 17678
rect 30828 16772 30884 17612
rect 30940 16882 30996 18396
rect 31052 17668 31108 20078
rect 31164 20132 31220 20142
rect 31164 19122 31220 20076
rect 31724 20132 31780 20142
rect 31836 20132 31892 21420
rect 32620 21364 32676 21374
rect 32060 21140 32116 21150
rect 31948 20916 32004 20926
rect 31948 20822 32004 20860
rect 31724 20130 31892 20132
rect 31724 20078 31726 20130
rect 31778 20078 31892 20130
rect 31724 20076 31892 20078
rect 31724 20066 31780 20076
rect 31948 20020 32004 20030
rect 32060 20020 32116 21084
rect 32396 20804 32452 20814
rect 32396 20710 32452 20748
rect 31948 20018 32116 20020
rect 31948 19966 31950 20018
rect 32002 19966 32116 20018
rect 31948 19964 32116 19966
rect 32508 20692 32564 20702
rect 32508 20244 32564 20636
rect 32620 20468 32676 21308
rect 32956 20916 33012 21644
rect 33068 21586 33124 21598
rect 33068 21534 33070 21586
rect 33122 21534 33124 21586
rect 33068 21364 33124 21534
rect 33068 21298 33124 21308
rect 33068 21140 33124 21150
rect 33180 21140 33236 22204
rect 33292 22194 33348 22204
rect 33292 21812 33348 21822
rect 33292 21718 33348 21756
rect 33292 21588 33348 21598
rect 33292 21494 33348 21532
rect 33124 21084 33236 21140
rect 33068 21074 33124 21084
rect 33068 20916 33124 20926
rect 32956 20914 33124 20916
rect 32956 20862 33070 20914
rect 33122 20862 33124 20914
rect 32956 20860 33124 20862
rect 33068 20850 33124 20860
rect 33404 20580 33460 23548
rect 33852 23492 33908 27804
rect 34188 27748 34244 27806
rect 34188 27682 34244 27692
rect 34076 27300 34132 27310
rect 33964 26964 34020 26974
rect 33964 26870 34020 26908
rect 34076 25844 34132 27244
rect 34300 26908 34356 28252
rect 34188 26852 34356 26908
rect 34188 26178 34244 26852
rect 34188 26126 34190 26178
rect 34242 26126 34244 26178
rect 34188 25844 34244 26126
rect 34412 26068 34468 29932
rect 34524 29540 34580 29550
rect 34524 27972 34580 29484
rect 34748 29426 34804 29438
rect 34748 29374 34750 29426
rect 34802 29374 34804 29426
rect 34636 28420 34692 28430
rect 34636 28326 34692 28364
rect 34748 28308 34804 29374
rect 34972 28868 35028 29932
rect 35084 29986 35140 29998
rect 35084 29934 35086 29986
rect 35138 29934 35140 29986
rect 35084 29540 35140 29934
rect 35084 29474 35140 29484
rect 35308 29986 35364 29998
rect 35308 29934 35310 29986
rect 35362 29934 35364 29986
rect 35308 29540 35364 29934
rect 35532 29652 35588 29662
rect 35308 29474 35364 29484
rect 35420 29596 35532 29652
rect 34748 28242 34804 28252
rect 34860 28812 35028 28868
rect 35084 29316 35140 29326
rect 34748 27972 34804 27982
rect 34524 27970 34804 27972
rect 34524 27918 34750 27970
rect 34802 27918 34804 27970
rect 34524 27916 34804 27918
rect 34748 27906 34804 27916
rect 34860 27970 34916 28812
rect 34972 28644 35028 28654
rect 35084 28644 35140 29260
rect 35196 29314 35252 29326
rect 35196 29262 35198 29314
rect 35250 29262 35252 29314
rect 35196 29204 35252 29262
rect 35308 29316 35364 29326
rect 35420 29316 35476 29596
rect 35532 29586 35588 29596
rect 35644 29540 35700 30158
rect 35868 30210 36148 30212
rect 35868 30158 36094 30210
rect 36146 30158 36148 30210
rect 35868 30156 36148 30158
rect 35756 29988 35812 29998
rect 35756 29894 35812 29932
rect 35868 29876 35924 30156
rect 36092 30146 36148 30156
rect 35980 29988 36036 29998
rect 35980 29986 36372 29988
rect 35980 29934 35982 29986
rect 36034 29934 36372 29986
rect 35980 29932 36372 29934
rect 35980 29922 36036 29932
rect 35868 29810 35924 29820
rect 35980 29652 36036 29662
rect 35644 29484 35812 29540
rect 35308 29314 35476 29316
rect 35308 29262 35310 29314
rect 35362 29262 35476 29314
rect 35308 29260 35476 29262
rect 35532 29426 35588 29438
rect 35532 29374 35534 29426
rect 35586 29374 35588 29426
rect 35532 29316 35588 29374
rect 35644 29316 35700 29326
rect 35532 29260 35644 29316
rect 35308 29250 35364 29260
rect 35644 29250 35700 29260
rect 35196 29138 35252 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34972 28642 35140 28644
rect 34972 28590 34974 28642
rect 35026 28590 35140 28642
rect 34972 28588 35140 28590
rect 35196 28868 35252 28878
rect 35756 28868 35812 29484
rect 35980 29428 36036 29596
rect 35980 29426 36148 29428
rect 35980 29374 35982 29426
rect 36034 29374 36148 29426
rect 35980 29372 36148 29374
rect 35980 29362 36036 29372
rect 35196 28754 35252 28812
rect 35196 28702 35198 28754
rect 35250 28702 35252 28754
rect 35196 28644 35252 28702
rect 34972 28578 35028 28588
rect 35196 28578 35252 28588
rect 35420 28812 35812 28868
rect 35868 28868 35924 28878
rect 34860 27918 34862 27970
rect 34914 27918 34916 27970
rect 34860 27906 34916 27918
rect 34972 28420 35028 28430
rect 34860 27188 34916 27198
rect 34972 27188 35028 28364
rect 35420 27636 35476 28812
rect 35532 28642 35588 28654
rect 35532 28590 35534 28642
rect 35586 28590 35588 28642
rect 35532 28308 35588 28590
rect 35532 28242 35588 28252
rect 35756 28642 35812 28654
rect 35756 28590 35758 28642
rect 35810 28590 35812 28642
rect 35756 28084 35812 28590
rect 35532 28028 35812 28084
rect 35532 27860 35588 28028
rect 35532 27766 35588 27804
rect 35756 27858 35812 27870
rect 35756 27806 35758 27858
rect 35810 27806 35812 27858
rect 35756 27748 35812 27806
rect 35868 27860 35924 28812
rect 35980 28644 36036 28654
rect 35980 28550 36036 28588
rect 36092 28308 36148 29372
rect 36204 29426 36260 29438
rect 36204 29374 36206 29426
rect 36258 29374 36260 29426
rect 36204 29092 36260 29374
rect 36204 29026 36260 29036
rect 36092 28242 36148 28252
rect 36204 28420 36260 28430
rect 35980 27860 36036 27870
rect 35868 27858 36036 27860
rect 35868 27806 35982 27858
rect 36034 27806 36036 27858
rect 35868 27804 36036 27806
rect 35980 27794 36036 27804
rect 35756 27692 35924 27748
rect 34916 27132 35028 27188
rect 35084 27580 35476 27636
rect 34860 27074 34916 27132
rect 34860 27022 34862 27074
rect 34914 27022 34916 27074
rect 34860 27010 34916 27022
rect 34524 26964 34580 27002
rect 35084 26908 35140 27580
rect 35868 27524 35924 27692
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35756 27076 35812 27086
rect 34524 26898 34580 26908
rect 34972 26852 35140 26908
rect 35196 26964 35252 27002
rect 35196 26898 35252 26908
rect 34524 26292 34580 26302
rect 34524 26198 34580 26236
rect 34748 26180 34804 26190
rect 34748 26086 34804 26124
rect 34412 26012 34580 26068
rect 34188 25788 34468 25844
rect 34076 25778 34132 25788
rect 34412 25730 34468 25788
rect 34412 25678 34414 25730
rect 34466 25678 34468 25730
rect 34412 25666 34468 25678
rect 34300 25620 34356 25630
rect 34188 25564 34300 25620
rect 34188 25506 34244 25564
rect 34300 25554 34356 25564
rect 34188 25454 34190 25506
rect 34242 25454 34244 25506
rect 34188 25442 34244 25454
rect 34412 25284 34468 25294
rect 34300 24164 34356 24174
rect 34188 23938 34244 23950
rect 34188 23886 34190 23938
rect 34242 23886 34244 23938
rect 33852 23436 34132 23492
rect 33852 23268 33908 23278
rect 33516 22370 33572 22382
rect 33852 22372 33908 23212
rect 33516 22318 33518 22370
rect 33570 22318 33572 22370
rect 33516 22036 33572 22318
rect 33516 21970 33572 21980
rect 33628 22370 33908 22372
rect 33628 22318 33854 22370
rect 33906 22318 33908 22370
rect 33628 22316 33908 22318
rect 33628 21698 33684 22316
rect 33852 22306 33908 22316
rect 33964 22372 34020 22382
rect 33628 21646 33630 21698
rect 33682 21646 33684 21698
rect 33628 21634 33684 21646
rect 33852 22146 33908 22158
rect 33852 22094 33854 22146
rect 33906 22094 33908 22146
rect 33852 20916 33908 22094
rect 33964 21810 34020 22316
rect 34076 22148 34132 23436
rect 34188 23268 34244 23886
rect 34300 23826 34356 24108
rect 34300 23774 34302 23826
rect 34354 23774 34356 23826
rect 34300 23762 34356 23774
rect 34300 23380 34356 23390
rect 34412 23380 34468 25228
rect 34300 23378 34468 23380
rect 34300 23326 34302 23378
rect 34354 23326 34468 23378
rect 34300 23324 34468 23326
rect 34300 23314 34356 23324
rect 34188 23202 34244 23212
rect 34524 22820 34580 26012
rect 34524 22754 34580 22764
rect 34748 25730 34804 25742
rect 34748 25678 34750 25730
rect 34802 25678 34804 25730
rect 34748 24948 34804 25678
rect 34860 25620 34916 25630
rect 34972 25620 35028 26852
rect 35532 26850 35588 26862
rect 35532 26798 35534 26850
rect 35586 26798 35588 26850
rect 34860 25618 35028 25620
rect 34860 25566 34862 25618
rect 34914 25566 35028 25618
rect 34860 25564 35028 25566
rect 35084 26066 35140 26078
rect 35084 26014 35086 26066
rect 35138 26014 35140 26066
rect 35084 25620 35140 26014
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34860 25554 34916 25564
rect 35084 25554 35140 25564
rect 35420 25508 35476 25518
rect 35420 25414 35476 25452
rect 35084 25396 35140 25406
rect 35084 25302 35140 25340
rect 34524 22596 34580 22606
rect 34524 22260 34580 22540
rect 34412 22258 34580 22260
rect 34412 22206 34526 22258
rect 34578 22206 34580 22258
rect 34412 22204 34580 22206
rect 34188 22148 34244 22158
rect 34076 22146 34244 22148
rect 34076 22094 34190 22146
rect 34242 22094 34244 22146
rect 34076 22092 34244 22094
rect 33964 21758 33966 21810
rect 34018 21758 34020 21810
rect 33964 21746 34020 21758
rect 34188 21252 34244 22092
rect 34300 21476 34356 21486
rect 34300 21382 34356 21420
rect 34188 21196 34356 21252
rect 33852 20850 33908 20860
rect 32620 20402 32676 20412
rect 32844 20524 33460 20580
rect 32508 20018 32564 20188
rect 32508 19966 32510 20018
rect 32562 19966 32564 20018
rect 31948 19348 32004 19964
rect 32508 19954 32564 19966
rect 31948 19282 32004 19292
rect 32732 19908 32788 19918
rect 31164 19070 31166 19122
rect 31218 19070 31220 19122
rect 31164 19058 31220 19070
rect 32508 19010 32564 19022
rect 32508 18958 32510 19010
rect 32562 18958 32564 19010
rect 32396 18452 32452 18462
rect 32508 18452 32564 18958
rect 32732 18564 32788 19852
rect 32732 18498 32788 18508
rect 32452 18396 32564 18452
rect 32396 18358 32452 18396
rect 31052 17602 31108 17612
rect 31948 18338 32004 18350
rect 31948 18286 31950 18338
rect 32002 18286 32004 18338
rect 31948 17668 32004 18286
rect 31948 17602 32004 17612
rect 32396 17556 32452 17566
rect 32396 17462 32452 17500
rect 32172 17444 32228 17454
rect 31612 16994 31668 17006
rect 31612 16942 31614 16994
rect 31666 16942 31668 16994
rect 31276 16884 31332 16894
rect 30940 16830 30942 16882
rect 30994 16830 30996 16882
rect 30940 16818 30996 16830
rect 31052 16882 31332 16884
rect 31052 16830 31278 16882
rect 31330 16830 31332 16882
rect 31052 16828 31332 16830
rect 30828 16706 30884 16716
rect 30716 16594 30772 16604
rect 30716 16212 30772 16222
rect 31052 16212 31108 16828
rect 31276 16818 31332 16828
rect 30604 16210 30772 16212
rect 30604 16158 30718 16210
rect 30770 16158 30772 16210
rect 30604 16156 30772 16158
rect 30716 16146 30772 16156
rect 30828 16156 31108 16212
rect 30716 15540 30772 15550
rect 30828 15540 30884 16156
rect 31500 16098 31556 16110
rect 31500 16046 31502 16098
rect 31554 16046 31556 16098
rect 30772 15484 30884 15540
rect 30940 15986 30996 15998
rect 30940 15934 30942 15986
rect 30994 15934 30996 15986
rect 30716 15446 30772 15484
rect 30492 15250 30548 15260
rect 30940 15148 30996 15934
rect 30716 15092 30996 15148
rect 31500 15428 31556 16046
rect 30604 14756 30660 14766
rect 29932 14532 29988 14542
rect 29932 14530 30100 14532
rect 29932 14478 29934 14530
rect 29986 14478 30100 14530
rect 29932 14476 30100 14478
rect 29932 14466 29988 14476
rect 29932 13748 29988 13758
rect 29932 13654 29988 13692
rect 30044 13524 30100 14476
rect 30156 14420 30212 14430
rect 30156 13748 30212 14364
rect 30380 14418 30436 14430
rect 30380 14366 30382 14418
rect 30434 14366 30436 14418
rect 30380 14308 30436 14366
rect 30380 14242 30436 14252
rect 30156 13692 30324 13748
rect 30044 13458 30100 13468
rect 30268 13300 30324 13692
rect 30492 13746 30548 13758
rect 30492 13694 30494 13746
rect 30546 13694 30548 13746
rect 30156 13244 30324 13300
rect 30380 13634 30436 13646
rect 30380 13582 30382 13634
rect 30434 13582 30436 13634
rect 30156 13074 30212 13244
rect 30156 13022 30158 13074
rect 30210 13022 30212 13074
rect 30156 13010 30212 13022
rect 30268 13076 30324 13086
rect 29932 12628 29988 12638
rect 29932 12404 29988 12572
rect 29932 12310 29988 12348
rect 30268 12068 30324 13020
rect 29932 11732 29988 11742
rect 29932 10610 29988 11676
rect 30268 11284 30324 12012
rect 30380 11508 30436 13582
rect 30492 11620 30548 13694
rect 30604 13076 30660 14700
rect 30716 13524 30772 15092
rect 31164 14756 31220 14766
rect 31164 14662 31220 14700
rect 30716 13458 30772 13468
rect 30828 14306 30884 14318
rect 30828 14254 30830 14306
rect 30882 14254 30884 14306
rect 30828 13746 30884 14254
rect 30828 13694 30830 13746
rect 30882 13694 30884 13746
rect 30828 13300 30884 13694
rect 30828 13234 30884 13244
rect 30940 13748 30996 13758
rect 30604 13010 30660 13020
rect 30604 12852 30660 12862
rect 30604 12758 30660 12796
rect 30604 12180 30660 12190
rect 30604 12086 30660 12124
rect 30604 11620 30660 11630
rect 30492 11564 30604 11620
rect 30604 11526 30660 11564
rect 30828 11620 30884 11630
rect 30380 11452 30548 11508
rect 30380 11284 30436 11294
rect 30268 11282 30436 11284
rect 30268 11230 30382 11282
rect 30434 11230 30436 11282
rect 30268 11228 30436 11230
rect 30380 11218 30436 11228
rect 29932 10558 29934 10610
rect 29986 10558 29988 10610
rect 29932 10546 29988 10558
rect 29820 10332 30212 10388
rect 29820 9714 29876 9726
rect 29820 9662 29822 9714
rect 29874 9662 29876 9714
rect 29708 9492 29764 9502
rect 29708 9154 29764 9436
rect 29820 9268 29876 9662
rect 29932 9716 29988 9726
rect 29932 9622 29988 9660
rect 29820 9202 29876 9212
rect 29708 9102 29710 9154
rect 29762 9102 29764 9154
rect 29708 9090 29764 9102
rect 29820 8930 29876 8942
rect 29820 8878 29822 8930
rect 29874 8878 29876 8930
rect 29820 8372 29876 8878
rect 30044 8818 30100 8830
rect 30044 8766 30046 8818
rect 30098 8766 30100 8818
rect 29932 8372 29988 8382
rect 29820 8370 29988 8372
rect 29820 8318 29934 8370
rect 29986 8318 29988 8370
rect 29820 8316 29988 8318
rect 29932 8306 29988 8316
rect 29372 7196 29652 7252
rect 29708 8148 29764 8158
rect 29708 7474 29764 8092
rect 29932 7700 29988 7710
rect 29932 7588 29988 7644
rect 30044 7698 30100 8766
rect 30044 7646 30046 7698
rect 30098 7646 30100 7698
rect 30044 7634 30100 7646
rect 29708 7422 29710 7474
rect 29762 7422 29764 7474
rect 29148 5796 29204 5806
rect 29148 5702 29204 5740
rect 28924 4562 29092 4564
rect 28924 4510 28926 4562
rect 28978 4510 29092 4562
rect 28924 4508 29092 4510
rect 29260 4564 29316 4574
rect 28924 4498 28980 4508
rect 29260 4470 29316 4508
rect 28476 4062 28478 4114
rect 28530 4062 28532 4114
rect 28476 4050 28532 4062
rect 27916 3666 28084 3668
rect 27916 3614 27918 3666
rect 27970 3614 28084 3666
rect 27916 3612 28084 3614
rect 28924 3668 28980 3678
rect 29372 3668 29428 7196
rect 29484 6578 29540 6590
rect 29484 6526 29486 6578
rect 29538 6526 29540 6578
rect 29484 6356 29540 6526
rect 29596 6580 29652 6590
rect 29596 6486 29652 6524
rect 29708 6356 29764 7422
rect 29820 7586 29988 7588
rect 29820 7534 29934 7586
rect 29986 7534 29988 7586
rect 29820 7532 29988 7534
rect 29820 6804 29876 7532
rect 29932 7522 29988 7532
rect 30156 7476 30212 10332
rect 30492 10052 30548 11452
rect 30716 10612 30772 10622
rect 30716 10518 30772 10556
rect 30492 9938 30548 9996
rect 30492 9886 30494 9938
rect 30546 9886 30548 9938
rect 30492 9874 30548 9886
rect 30268 9826 30324 9838
rect 30268 9774 30270 9826
rect 30322 9774 30324 9826
rect 30268 9380 30324 9774
rect 30268 9314 30324 9324
rect 30268 8932 30324 8942
rect 30268 8838 30324 8876
rect 30828 8260 30884 11564
rect 30940 9266 30996 13692
rect 31164 13524 31220 13534
rect 31052 12964 31108 12974
rect 31164 12964 31220 13468
rect 31388 13300 31444 13310
rect 31052 12962 31220 12964
rect 31052 12910 31054 12962
rect 31106 12910 31220 12962
rect 31052 12908 31220 12910
rect 31276 12964 31332 12974
rect 31052 12898 31108 12908
rect 31164 12740 31220 12750
rect 31052 12404 31108 12414
rect 31052 10050 31108 12348
rect 31052 9998 31054 10050
rect 31106 9998 31108 10050
rect 31052 9986 31108 9998
rect 31164 9716 31220 12684
rect 31276 12292 31332 12908
rect 31276 12226 31332 12236
rect 31388 11394 31444 13244
rect 31388 11342 31390 11394
rect 31442 11342 31444 11394
rect 31388 11330 31444 11342
rect 31388 11172 31444 11182
rect 31388 10724 31444 11116
rect 31500 10836 31556 15372
rect 31612 15988 31668 16942
rect 32060 16996 32116 17006
rect 32060 16902 32116 16940
rect 32172 16994 32228 17388
rect 32172 16942 32174 16994
rect 32226 16942 32228 16994
rect 32172 16930 32228 16942
rect 31948 16884 32004 16894
rect 31948 16660 32004 16828
rect 32060 16660 32116 16670
rect 31948 16658 32116 16660
rect 31948 16606 32062 16658
rect 32114 16606 32116 16658
rect 31948 16604 32116 16606
rect 32060 16594 32116 16604
rect 31724 16100 31780 16110
rect 32060 16100 32116 16110
rect 31724 16098 32116 16100
rect 31724 16046 31726 16098
rect 31778 16046 32062 16098
rect 32114 16046 32116 16098
rect 31724 16044 32116 16046
rect 31724 16034 31780 16044
rect 31612 14644 31668 15932
rect 31612 14578 31668 14588
rect 31836 14530 31892 16044
rect 32060 15538 32116 16044
rect 32060 15486 32062 15538
rect 32114 15486 32116 15538
rect 32060 15474 32116 15486
rect 32620 16098 32676 16110
rect 32620 16046 32622 16098
rect 32674 16046 32676 16098
rect 31836 14478 31838 14530
rect 31890 14478 31892 14530
rect 31836 14466 31892 14478
rect 32284 14532 32340 14542
rect 32284 14438 32340 14476
rect 31724 14418 31780 14430
rect 31724 14366 31726 14418
rect 31778 14366 31780 14418
rect 31724 14308 31780 14366
rect 31836 14308 31892 14318
rect 31724 14252 31836 14308
rect 31836 14242 31892 14252
rect 32284 13972 32340 13982
rect 32172 13916 32284 13972
rect 31724 13748 31780 13758
rect 31724 11508 31780 13692
rect 31836 13746 31892 13758
rect 31836 13694 31838 13746
rect 31890 13694 31892 13746
rect 31836 12964 31892 13694
rect 31836 12898 31892 12908
rect 31948 12180 32004 12190
rect 31836 12178 32004 12180
rect 31836 12126 31950 12178
rect 32002 12126 32004 12178
rect 31836 12124 32004 12126
rect 31836 12068 31892 12124
rect 31948 12114 32004 12124
rect 31836 12002 31892 12012
rect 31836 11508 31892 11518
rect 31724 11506 31892 11508
rect 31724 11454 31838 11506
rect 31890 11454 31892 11506
rect 31724 11452 31892 11454
rect 31836 11442 31892 11452
rect 32172 11172 32228 13916
rect 32284 13878 32340 13916
rect 32620 12852 32676 16046
rect 32620 12786 32676 12796
rect 32844 12404 32900 20524
rect 32956 20244 33012 20254
rect 32956 18676 33012 20188
rect 33516 20020 33572 20030
rect 33516 19906 33572 19964
rect 33516 19854 33518 19906
rect 33570 19854 33572 19906
rect 33516 19842 33572 19854
rect 33628 20018 33684 20030
rect 33628 19966 33630 20018
rect 33682 19966 33684 20018
rect 33292 19460 33348 19470
rect 33068 19236 33124 19246
rect 33068 19234 33236 19236
rect 33068 19182 33070 19234
rect 33122 19182 33236 19234
rect 33068 19180 33236 19182
rect 33068 19170 33124 19180
rect 33180 18900 33236 19180
rect 33292 19124 33348 19404
rect 33628 19348 33684 19966
rect 34188 20020 34244 20030
rect 34188 19926 34244 19964
rect 34076 19794 34132 19806
rect 34076 19742 34078 19794
rect 34130 19742 34132 19794
rect 33852 19348 33908 19358
rect 33628 19292 33852 19348
rect 33852 19124 33908 19292
rect 34076 19124 34132 19742
rect 34188 19236 34244 19246
rect 34188 19142 34244 19180
rect 33292 19122 33796 19124
rect 33292 19070 33294 19122
rect 33346 19070 33796 19122
rect 33292 19068 33796 19070
rect 33292 19058 33348 19068
rect 33180 18844 33572 18900
rect 33180 18676 33236 18686
rect 32956 18674 33236 18676
rect 32956 18622 33182 18674
rect 33234 18622 33236 18674
rect 32956 18620 33236 18622
rect 33180 18610 33236 18620
rect 33068 18452 33124 18462
rect 33068 18358 33124 18396
rect 33516 18452 33572 18844
rect 33740 18562 33796 19068
rect 33852 19122 34020 19124
rect 33852 19070 33854 19122
rect 33906 19070 34020 19122
rect 33852 19068 34020 19070
rect 33852 19058 33908 19068
rect 33740 18510 33742 18562
rect 33794 18510 33796 18562
rect 33740 18498 33796 18510
rect 33628 18452 33684 18462
rect 33516 18450 33684 18452
rect 33516 18398 33630 18450
rect 33682 18398 33684 18450
rect 33516 18396 33684 18398
rect 33516 17892 33572 18396
rect 33628 18386 33684 18396
rect 33516 17826 33572 17836
rect 33740 18340 33796 18350
rect 33292 17108 33348 17118
rect 33292 16884 33348 17052
rect 33180 16882 33348 16884
rect 33180 16830 33294 16882
rect 33346 16830 33348 16882
rect 33180 16828 33348 16830
rect 32956 16436 33012 16446
rect 32956 16098 33012 16380
rect 32956 16046 32958 16098
rect 33010 16046 33012 16098
rect 32956 16034 33012 16046
rect 33068 15988 33124 15998
rect 33068 15894 33124 15932
rect 33180 15764 33236 16828
rect 33292 16818 33348 16828
rect 33516 16994 33572 17006
rect 33516 16942 33518 16994
rect 33570 16942 33572 16994
rect 33516 16212 33572 16942
rect 33516 16098 33572 16156
rect 33516 16046 33518 16098
rect 33570 16046 33572 16098
rect 33516 16034 33572 16046
rect 33628 16660 33684 16670
rect 33292 15876 33348 15886
rect 33292 15874 33572 15876
rect 33292 15822 33294 15874
rect 33346 15822 33572 15874
rect 33292 15820 33572 15822
rect 33292 15810 33348 15820
rect 32956 15708 33236 15764
rect 32956 14980 33012 15708
rect 33180 15428 33236 15438
rect 33180 15334 33236 15372
rect 33516 15426 33572 15820
rect 33516 15374 33518 15426
rect 33570 15374 33572 15426
rect 33516 15362 33572 15374
rect 33628 15764 33684 16604
rect 33628 15314 33684 15708
rect 33628 15262 33630 15314
rect 33682 15262 33684 15314
rect 33628 15250 33684 15262
rect 32956 14914 33012 14924
rect 33068 15090 33124 15102
rect 33068 15038 33070 15090
rect 33122 15038 33124 15090
rect 33068 14756 33124 15038
rect 33068 14690 33124 14700
rect 33404 14756 33460 14766
rect 33404 14662 33460 14700
rect 33292 14642 33348 14654
rect 33292 14590 33294 14642
rect 33346 14590 33348 14642
rect 33068 14530 33124 14542
rect 33068 14478 33070 14530
rect 33122 14478 33124 14530
rect 33068 14420 33124 14478
rect 33068 14354 33124 14364
rect 33292 13748 33348 14590
rect 33404 14420 33460 14430
rect 33404 13860 33460 14364
rect 33404 13766 33460 13804
rect 33292 13654 33348 13692
rect 33292 12516 33348 12526
rect 33740 12516 33796 18284
rect 33852 18228 33908 18238
rect 33852 17106 33908 18172
rect 33964 17890 34020 19068
rect 34076 19058 34132 19068
rect 34300 19012 34356 21196
rect 34300 18946 34356 18956
rect 33964 17838 33966 17890
rect 34018 17838 34020 17890
rect 33964 17826 34020 17838
rect 34076 18452 34132 18462
rect 33852 17054 33854 17106
rect 33906 17054 33908 17106
rect 33852 17042 33908 17054
rect 34076 17106 34132 18396
rect 34076 17054 34078 17106
rect 34130 17054 34132 17106
rect 34076 17042 34132 17054
rect 34412 17108 34468 22204
rect 34524 22194 34580 22204
rect 34524 21700 34580 21710
rect 34524 21586 34580 21644
rect 34524 21534 34526 21586
rect 34578 21534 34580 21586
rect 34524 21522 34580 21534
rect 34748 21588 34804 24892
rect 35532 24724 35588 26798
rect 35756 25508 35812 27020
rect 35868 26964 35924 27468
rect 35868 26898 35924 26908
rect 35756 25442 35812 25452
rect 36092 25394 36148 25406
rect 36092 25342 36094 25394
rect 36146 25342 36148 25394
rect 35756 25284 35812 25294
rect 35756 25190 35812 25228
rect 35308 24500 35364 24510
rect 35084 24498 35364 24500
rect 35084 24446 35310 24498
rect 35362 24446 35364 24498
rect 35084 24444 35364 24446
rect 35084 24164 35140 24444
rect 35308 24434 35364 24444
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 24164 35252 24174
rect 35140 24162 35252 24164
rect 35140 24110 35198 24162
rect 35250 24110 35252 24162
rect 35140 24108 35252 24110
rect 35084 24070 35140 24108
rect 35196 24098 35252 24108
rect 35420 23826 35476 23838
rect 35420 23774 35422 23826
rect 35474 23774 35476 23826
rect 34860 23716 34916 23726
rect 34860 23622 34916 23660
rect 35084 23716 35140 23726
rect 34860 22146 34916 22158
rect 34860 22094 34862 22146
rect 34914 22094 34916 22146
rect 34860 21588 34916 22094
rect 34972 21588 35028 21598
rect 34860 21586 35028 21588
rect 34860 21534 34974 21586
rect 35026 21534 35028 21586
rect 34860 21532 35028 21534
rect 34748 21522 34804 21532
rect 34972 20804 35028 21532
rect 35084 20916 35140 23660
rect 35420 23378 35476 23774
rect 35420 23326 35422 23378
rect 35474 23326 35476 23378
rect 35420 23156 35476 23326
rect 35420 23090 35476 23100
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 22596 35252 22606
rect 35196 22370 35252 22540
rect 35196 22318 35198 22370
rect 35250 22318 35252 22370
rect 35196 22306 35252 22318
rect 35532 21700 35588 24668
rect 35756 23940 35812 23950
rect 35756 23826 35812 23884
rect 35756 23774 35758 23826
rect 35810 23774 35812 23826
rect 35756 23762 35812 23774
rect 36092 23716 36148 25342
rect 36092 23650 36148 23660
rect 35868 23268 35924 23278
rect 35868 23174 35924 23212
rect 36092 23156 36148 23166
rect 36092 23062 36148 23100
rect 35868 22932 35924 22942
rect 35868 22370 35924 22876
rect 35868 22318 35870 22370
rect 35922 22318 35924 22370
rect 35868 22306 35924 22318
rect 35532 21634 35588 21644
rect 35980 22146 36036 22158
rect 35980 22094 35982 22146
rect 36034 22094 36036 22146
rect 35756 21588 35812 21598
rect 35756 21494 35812 21532
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 20916 35252 20926
rect 35084 20914 35252 20916
rect 35084 20862 35198 20914
rect 35250 20862 35252 20914
rect 35084 20860 35252 20862
rect 35196 20850 35252 20860
rect 34972 20692 35028 20748
rect 35084 20692 35140 20702
rect 34972 20636 35084 20692
rect 35084 20626 35140 20636
rect 35868 20690 35924 20702
rect 35868 20638 35870 20690
rect 35922 20638 35924 20690
rect 35532 20578 35588 20590
rect 35532 20526 35534 20578
rect 35586 20526 35588 20578
rect 35308 20244 35364 20254
rect 35532 20244 35588 20526
rect 35364 20188 35588 20244
rect 35756 20578 35812 20590
rect 35756 20526 35758 20578
rect 35810 20526 35812 20578
rect 35308 20178 35364 20188
rect 34748 20132 34804 20142
rect 34748 19122 34804 20076
rect 34748 19070 34750 19122
rect 34802 19070 34804 19122
rect 34748 18676 34804 19070
rect 34860 20130 34916 20142
rect 34860 20078 34862 20130
rect 34914 20078 34916 20130
rect 34860 18788 34916 20078
rect 34972 20132 35028 20142
rect 34972 19348 35028 20076
rect 35756 20132 35812 20526
rect 35756 20066 35812 20076
rect 35196 19908 35252 19918
rect 35252 19852 35700 19908
rect 35196 19842 35252 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34972 19234 35028 19292
rect 34972 19182 34974 19234
rect 35026 19182 35028 19234
rect 34972 19170 35028 19182
rect 35420 19348 35476 19358
rect 34860 18732 35252 18788
rect 34748 18610 34804 18620
rect 35084 18452 35140 18490
rect 35084 18386 35140 18396
rect 35196 18340 35252 18732
rect 35196 18274 35252 18284
rect 35420 18338 35476 19292
rect 35420 18286 35422 18338
rect 35474 18286 35476 18338
rect 35084 18228 35140 18238
rect 34972 18226 35140 18228
rect 34972 18174 35086 18226
rect 35138 18174 35140 18226
rect 34972 18172 35140 18174
rect 34412 17042 34468 17052
rect 34524 17780 34580 17790
rect 34524 16882 34580 17724
rect 34972 17668 35028 18172
rect 35084 18162 35140 18172
rect 35420 18228 35476 18286
rect 35420 18162 35476 18172
rect 35532 18788 35588 18798
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35532 17780 35588 18732
rect 35644 18564 35700 19852
rect 35756 19236 35812 19246
rect 35868 19236 35924 20638
rect 35980 20132 36036 22094
rect 36204 21140 36260 28364
rect 36316 27186 36372 29932
rect 36652 29652 36708 29662
rect 36652 29558 36708 29596
rect 36540 29540 36596 29550
rect 36540 29446 36596 29484
rect 36428 29428 36484 29438
rect 36428 28866 36484 29372
rect 36764 29204 36820 35252
rect 36876 34692 36932 36988
rect 37212 36932 37268 37886
rect 37212 36866 37268 36876
rect 37100 35700 37156 35710
rect 37100 35026 37156 35644
rect 37100 34974 37102 35026
rect 37154 34974 37156 35026
rect 37100 34962 37156 34974
rect 36876 34626 36932 34636
rect 37212 34580 37268 34590
rect 36876 34130 36932 34142
rect 36876 34078 36878 34130
rect 36930 34078 36932 34130
rect 36876 31444 36932 34078
rect 37212 34132 37268 34524
rect 37324 34468 37380 38556
rect 37436 38610 37492 38622
rect 37436 38558 37438 38610
rect 37490 38558 37492 38610
rect 37436 37378 37492 38558
rect 37436 37326 37438 37378
rect 37490 37326 37492 37378
rect 37436 37044 37492 37326
rect 37436 36978 37492 36988
rect 37660 37826 37716 37838
rect 37660 37774 37662 37826
rect 37714 37774 37716 37826
rect 37436 36484 37492 36494
rect 37660 36484 37716 37774
rect 37884 37268 37940 39454
rect 38220 39508 38276 45276
rect 38780 45108 38836 46732
rect 40012 46674 40068 47404
rect 40236 46900 40292 47852
rect 40460 47460 40516 52108
rect 40572 51604 40628 51614
rect 40572 49924 40628 51548
rect 40572 49026 40628 49868
rect 40572 48974 40574 49026
rect 40626 48974 40628 49026
rect 40572 48962 40628 48974
rect 40684 47684 40740 53454
rect 40908 53060 40964 53070
rect 40908 52966 40964 53004
rect 41020 52388 41076 54348
rect 41132 54338 41188 54348
rect 41356 53844 41412 54462
rect 41356 53778 41412 53788
rect 41244 53620 41300 53630
rect 41580 53620 41636 57484
rect 41804 57474 41860 57484
rect 44044 57316 44100 57326
rect 42700 56978 42756 56990
rect 42700 56926 42702 56978
rect 42754 56926 42756 56978
rect 42588 56866 42644 56878
rect 42588 56814 42590 56866
rect 42642 56814 42644 56866
rect 42252 56756 42308 56766
rect 42252 56662 42308 56700
rect 42588 56308 42644 56814
rect 42588 56242 42644 56252
rect 42252 55970 42308 55982
rect 42252 55918 42254 55970
rect 42306 55918 42308 55970
rect 42252 55748 42308 55918
rect 42028 55692 42252 55748
rect 41916 55076 41972 55086
rect 41244 53618 41636 53620
rect 41244 53566 41246 53618
rect 41298 53566 41582 53618
rect 41634 53566 41636 53618
rect 41244 53564 41636 53566
rect 41244 53554 41300 53564
rect 41132 53284 41188 53294
rect 41132 52946 41188 53228
rect 41132 52894 41134 52946
rect 41186 52894 41188 52946
rect 41132 52882 41188 52894
rect 40908 52332 41076 52388
rect 40796 50482 40852 50494
rect 40796 50430 40798 50482
rect 40850 50430 40852 50482
rect 40796 50372 40852 50430
rect 40796 49812 40852 50316
rect 40796 49746 40852 49756
rect 40684 47618 40740 47628
rect 40908 47572 40964 52332
rect 41020 52052 41076 52062
rect 41020 51958 41076 51996
rect 41020 51268 41076 51278
rect 41020 51266 41412 51268
rect 41020 51214 41022 51266
rect 41074 51214 41412 51266
rect 41020 51212 41412 51214
rect 41020 51202 41076 51212
rect 41244 50596 41300 50606
rect 41020 50484 41076 50522
rect 41020 50418 41076 50428
rect 41132 50370 41188 50382
rect 41132 50318 41134 50370
rect 41186 50318 41188 50370
rect 41020 49810 41076 49822
rect 41020 49758 41022 49810
rect 41074 49758 41076 49810
rect 41020 48916 41076 49758
rect 41132 49252 41188 50318
rect 41132 49186 41188 49196
rect 41132 48916 41188 48926
rect 41244 48916 41300 50540
rect 41356 49700 41412 51212
rect 41580 50428 41636 53564
rect 41804 55074 41972 55076
rect 41804 55022 41918 55074
rect 41970 55022 41972 55074
rect 41804 55020 41972 55022
rect 41692 52834 41748 52846
rect 41692 52782 41694 52834
rect 41746 52782 41748 52834
rect 41692 51492 41748 52782
rect 41692 51426 41748 51436
rect 41692 50708 41748 50718
rect 41692 50614 41748 50652
rect 41804 50428 41860 55020
rect 41916 55010 41972 55020
rect 41916 53506 41972 53518
rect 41916 53454 41918 53506
rect 41970 53454 41972 53506
rect 41916 53284 41972 53454
rect 41916 53218 41972 53228
rect 42028 52612 42084 55692
rect 42252 55682 42308 55692
rect 42588 55300 42644 55310
rect 42588 55206 42644 55244
rect 42252 55074 42308 55086
rect 42252 55022 42254 55074
rect 42306 55022 42308 55074
rect 42252 54740 42308 55022
rect 42140 54404 42196 54414
rect 42140 54310 42196 54348
rect 42252 53732 42308 54684
rect 42252 53666 42308 53676
rect 42700 53732 42756 56926
rect 43484 56644 43540 56654
rect 43484 56642 43652 56644
rect 43484 56590 43486 56642
rect 43538 56590 43652 56642
rect 43484 56588 43652 56590
rect 43484 56578 43540 56588
rect 42812 56308 42868 56318
rect 42812 55186 42868 56252
rect 42924 56194 42980 56206
rect 42924 56142 42926 56194
rect 42978 56142 42980 56194
rect 42924 55410 42980 56142
rect 42924 55358 42926 55410
rect 42978 55358 42980 55410
rect 42924 55346 42980 55358
rect 43596 55972 43652 56588
rect 43372 55298 43428 55310
rect 43372 55246 43374 55298
rect 43426 55246 43428 55298
rect 42812 55134 42814 55186
rect 42866 55134 42868 55186
rect 42812 55122 42868 55134
rect 42924 55188 42980 55198
rect 42924 55094 42980 55132
rect 43372 54068 43428 55246
rect 43372 54002 43428 54012
rect 42700 53666 42756 53676
rect 43260 53730 43316 53742
rect 43260 53678 43262 53730
rect 43314 53678 43316 53730
rect 42364 53506 42420 53518
rect 42364 53454 42366 53506
rect 42418 53454 42420 53506
rect 42364 53396 42420 53454
rect 43036 53506 43092 53518
rect 43036 53454 43038 53506
rect 43090 53454 43092 53506
rect 42364 53330 42420 53340
rect 42812 53396 42868 53406
rect 42700 53058 42756 53070
rect 42700 53006 42702 53058
rect 42754 53006 42756 53058
rect 42028 52556 42196 52612
rect 42028 52388 42084 52398
rect 41916 52332 42028 52388
rect 41916 51490 41972 52332
rect 42028 52322 42084 52332
rect 42140 52164 42196 52556
rect 42700 52388 42756 53006
rect 42700 52322 42756 52332
rect 41916 51438 41918 51490
rect 41970 51438 41972 51490
rect 41916 51426 41972 51438
rect 42028 52108 42196 52164
rect 41580 50372 41748 50428
rect 41804 50372 41972 50428
rect 41356 49634 41412 49644
rect 41020 48914 41300 48916
rect 41020 48862 41134 48914
rect 41186 48862 41300 48914
rect 41020 48860 41300 48862
rect 41132 48850 41188 48860
rect 41468 48804 41524 48814
rect 41132 48692 41188 48702
rect 41132 48242 41188 48636
rect 41132 48190 41134 48242
rect 41186 48190 41188 48242
rect 41132 48178 41188 48190
rect 41468 48130 41524 48748
rect 41580 48356 41636 48366
rect 41580 48262 41636 48300
rect 41468 48078 41470 48130
rect 41522 48078 41524 48130
rect 41468 48066 41524 48078
rect 41580 47684 41636 47694
rect 41580 47590 41636 47628
rect 40908 47516 41412 47572
rect 40460 47404 40852 47460
rect 40796 47348 40852 47404
rect 40796 47292 41076 47348
rect 40572 47236 40628 47246
rect 40236 46834 40292 46844
rect 40348 47234 40628 47236
rect 40348 47182 40574 47234
rect 40626 47182 40628 47234
rect 40348 47180 40628 47182
rect 40012 46622 40014 46674
rect 40066 46622 40068 46674
rect 38780 45042 38836 45052
rect 39004 46452 39060 46462
rect 39004 45780 39060 46396
rect 39676 46116 39732 46126
rect 39676 46022 39732 46060
rect 38332 44884 38388 44894
rect 38332 44882 38500 44884
rect 38332 44830 38334 44882
rect 38386 44830 38500 44882
rect 38332 44828 38500 44830
rect 38332 44818 38388 44828
rect 38332 44098 38388 44110
rect 38332 44046 38334 44098
rect 38386 44046 38388 44098
rect 38332 42644 38388 44046
rect 38444 43652 38500 44828
rect 38444 43586 38500 43596
rect 38668 44322 38724 44334
rect 38668 44270 38670 44322
rect 38722 44270 38724 44322
rect 38556 43540 38612 43550
rect 38556 42644 38612 43484
rect 38332 42588 38500 42644
rect 38444 41972 38500 42588
rect 38556 42578 38612 42588
rect 38444 41906 38500 41916
rect 38332 41858 38388 41870
rect 38332 41806 38334 41858
rect 38386 41806 38388 41858
rect 38332 40516 38388 41806
rect 38668 41412 38724 44270
rect 38892 42756 38948 42766
rect 38892 42662 38948 42700
rect 38780 41412 38836 41422
rect 38668 41410 38836 41412
rect 38668 41358 38782 41410
rect 38834 41358 38836 41410
rect 38668 41356 38836 41358
rect 39004 41412 39060 45724
rect 39340 45666 39396 45678
rect 39340 45614 39342 45666
rect 39394 45614 39396 45666
rect 39228 45108 39284 45118
rect 39228 45014 39284 45052
rect 39340 44436 39396 45614
rect 39676 44994 39732 45006
rect 39676 44942 39678 44994
rect 39730 44942 39732 44994
rect 39676 44548 39732 44942
rect 39900 44884 39956 44894
rect 39900 44790 39956 44828
rect 39676 44482 39732 44492
rect 39228 44434 39396 44436
rect 39228 44382 39342 44434
rect 39394 44382 39396 44434
rect 39228 44380 39396 44382
rect 39116 44210 39172 44222
rect 39116 44158 39118 44210
rect 39170 44158 39172 44210
rect 39116 43540 39172 44158
rect 39116 43474 39172 43484
rect 39116 43316 39172 43326
rect 39228 43316 39284 44380
rect 39340 44370 39396 44380
rect 39564 44436 39620 44446
rect 39564 43538 39620 44380
rect 40012 43876 40068 46622
rect 40348 46004 40404 47180
rect 40572 47170 40628 47180
rect 40236 45948 40404 46004
rect 40460 46788 40516 46798
rect 40236 45892 40292 45948
rect 40124 45890 40292 45892
rect 40124 45838 40238 45890
rect 40290 45838 40292 45890
rect 40124 45836 40292 45838
rect 40124 44660 40180 45836
rect 40236 45826 40292 45836
rect 40348 45778 40404 45790
rect 40348 45726 40350 45778
rect 40402 45726 40404 45778
rect 40236 45444 40292 45454
rect 40236 45330 40292 45388
rect 40236 45278 40238 45330
rect 40290 45278 40292 45330
rect 40236 45266 40292 45278
rect 40348 45108 40404 45726
rect 40124 44594 40180 44604
rect 40236 44996 40292 45006
rect 40124 44436 40180 44446
rect 40124 44342 40180 44380
rect 40124 43876 40180 43886
rect 40012 43820 40124 43876
rect 39564 43486 39566 43538
rect 39618 43486 39620 43538
rect 39564 43474 39620 43486
rect 39116 43314 39284 43316
rect 39116 43262 39118 43314
rect 39170 43262 39284 43314
rect 39116 43260 39284 43262
rect 40012 43426 40068 43438
rect 40012 43374 40014 43426
rect 40066 43374 40068 43426
rect 39116 43250 39172 43260
rect 39900 43092 39956 43102
rect 39900 42978 39956 43036
rect 39900 42926 39902 42978
rect 39954 42926 39956 42978
rect 39900 42914 39956 42926
rect 39340 42644 39396 42654
rect 39396 42588 39508 42644
rect 39340 42578 39396 42588
rect 39116 41412 39172 41422
rect 39004 41410 39172 41412
rect 39004 41358 39118 41410
rect 39170 41358 39172 41410
rect 39004 41356 39172 41358
rect 38780 41346 38836 41356
rect 39116 41346 39172 41356
rect 39340 41300 39396 41310
rect 39452 41300 39508 42588
rect 39676 41970 39732 41982
rect 39676 41918 39678 41970
rect 39730 41918 39732 41970
rect 39340 41298 39508 41300
rect 39340 41246 39342 41298
rect 39394 41246 39508 41298
rect 39340 41244 39508 41246
rect 39564 41746 39620 41758
rect 39564 41694 39566 41746
rect 39618 41694 39620 41746
rect 39340 41234 39396 41244
rect 38444 40964 38500 40974
rect 38444 40870 38500 40908
rect 38332 40450 38388 40460
rect 39228 40514 39284 40526
rect 39228 40462 39230 40514
rect 39282 40462 39284 40514
rect 38220 39442 38276 39452
rect 38668 39844 38724 39854
rect 38668 39058 38724 39788
rect 39228 39844 39284 40462
rect 39564 40068 39620 41694
rect 39676 40964 39732 41918
rect 39676 40898 39732 40908
rect 39788 41860 39844 41870
rect 40012 41860 40068 43374
rect 39788 41858 40068 41860
rect 39788 41806 39790 41858
rect 39842 41806 40068 41858
rect 39788 41804 40068 41806
rect 39788 40852 39844 41804
rect 39788 40786 39844 40796
rect 40124 41186 40180 43820
rect 40236 43538 40292 44940
rect 40348 44548 40404 45052
rect 40348 44482 40404 44492
rect 40460 44210 40516 46732
rect 40908 46788 40964 46798
rect 40908 46694 40964 46732
rect 40796 46564 40852 46574
rect 40796 45332 40852 46508
rect 41020 45892 41076 47292
rect 41356 46676 41412 47516
rect 41692 46676 41748 50372
rect 41804 47460 41860 47470
rect 41804 47366 41860 47404
rect 41916 47012 41972 50372
rect 41916 46946 41972 46956
rect 42028 48468 42084 52108
rect 42476 50594 42532 50606
rect 42476 50542 42478 50594
rect 42530 50542 42532 50594
rect 42476 50428 42532 50542
rect 42700 50594 42756 50606
rect 42700 50542 42702 50594
rect 42754 50542 42756 50594
rect 42700 50428 42756 50542
rect 42812 50596 42868 53340
rect 43036 52388 43092 53454
rect 43036 52322 43092 52332
rect 43148 52276 43204 52286
rect 43260 52276 43316 53678
rect 43204 52220 43316 52276
rect 43148 52182 43204 52220
rect 42812 50530 42868 50540
rect 43036 52052 43092 52062
rect 43484 52052 43540 52062
rect 43036 50482 43092 51996
rect 43372 52050 43540 52052
rect 43372 51998 43486 52050
rect 43538 51998 43540 52050
rect 43372 51996 43540 51998
rect 43148 51604 43204 51614
rect 43148 51510 43204 51548
rect 43036 50430 43038 50482
rect 43090 50430 43092 50482
rect 42140 50372 42196 50382
rect 42476 50372 42644 50428
rect 42700 50372 42980 50428
rect 43036 50418 43092 50430
rect 43260 50594 43316 50606
rect 43260 50542 43262 50594
rect 43314 50542 43316 50594
rect 42140 50370 42308 50372
rect 42140 50318 42142 50370
rect 42194 50318 42308 50370
rect 42140 50316 42308 50318
rect 42140 50306 42196 50316
rect 42140 49924 42196 49934
rect 42140 49810 42196 49868
rect 42140 49758 42142 49810
rect 42194 49758 42196 49810
rect 42140 49746 42196 49758
rect 42252 49476 42308 50316
rect 42252 49420 42532 49476
rect 42364 49028 42420 49038
rect 42364 48934 42420 48972
rect 42364 48580 42420 48590
rect 42028 48242 42084 48412
rect 42028 48190 42030 48242
rect 42082 48190 42084 48242
rect 41356 46620 41636 46676
rect 41132 46452 41188 46462
rect 41132 46358 41188 46396
rect 41468 46450 41524 46462
rect 41468 46398 41470 46450
rect 41522 46398 41524 46450
rect 41356 45892 41412 45902
rect 41020 45890 41412 45892
rect 41020 45838 41358 45890
rect 41410 45838 41412 45890
rect 41020 45836 41412 45838
rect 41356 45826 41412 45836
rect 41132 45668 41188 45678
rect 41132 45666 41300 45668
rect 41132 45614 41134 45666
rect 41186 45614 41300 45666
rect 41132 45612 41300 45614
rect 41132 45602 41188 45612
rect 40908 45332 40964 45342
rect 40796 45330 40964 45332
rect 40796 45278 40910 45330
rect 40962 45278 40964 45330
rect 40796 45276 40964 45278
rect 40908 45266 40964 45276
rect 41132 45220 41188 45230
rect 41132 45106 41188 45164
rect 41132 45054 41134 45106
rect 41186 45054 41188 45106
rect 41132 45042 41188 45054
rect 41020 44436 41076 44446
rect 41020 44342 41076 44380
rect 40460 44158 40462 44210
rect 40514 44158 40516 44210
rect 40460 44146 40516 44158
rect 40908 43652 40964 43662
rect 40236 43486 40238 43538
rect 40290 43486 40292 43538
rect 40236 43474 40292 43486
rect 40796 43540 40852 43550
rect 40236 43204 40292 43214
rect 40236 42756 40292 43148
rect 40236 42662 40292 42700
rect 40796 42754 40852 43484
rect 40796 42702 40798 42754
rect 40850 42702 40852 42754
rect 40796 42690 40852 42702
rect 40908 42084 40964 43596
rect 41132 43538 41188 43550
rect 41132 43486 41134 43538
rect 41186 43486 41188 43538
rect 41132 43092 41188 43486
rect 41020 42980 41076 43018
rect 41020 42914 41076 42924
rect 40460 41970 40516 41982
rect 40460 41918 40462 41970
rect 40514 41918 40516 41970
rect 40460 41412 40516 41918
rect 40908 41970 40964 42028
rect 40908 41918 40910 41970
rect 40962 41918 40964 41970
rect 40908 41906 40964 41918
rect 41132 42082 41188 43036
rect 41132 42030 41134 42082
rect 41186 42030 41188 42082
rect 40796 41412 40852 41422
rect 40460 41410 40852 41412
rect 40460 41358 40798 41410
rect 40850 41358 40852 41410
rect 40460 41356 40852 41358
rect 40796 41346 40852 41356
rect 40124 41134 40126 41186
rect 40178 41134 40180 41186
rect 40124 40740 40180 41134
rect 40348 41244 40740 41300
rect 40348 41186 40404 41244
rect 40348 41134 40350 41186
rect 40402 41134 40404 41186
rect 40348 41122 40404 41134
rect 40684 41188 40740 41244
rect 41132 41188 41188 42030
rect 40684 41186 41188 41188
rect 40684 41134 41134 41186
rect 41186 41134 41188 41186
rect 40684 41132 41188 41134
rect 41132 41122 41188 41132
rect 40572 41076 40628 41086
rect 40572 40982 40628 41020
rect 40460 40962 40516 40974
rect 40460 40910 40462 40962
rect 40514 40910 40516 40962
rect 40124 40684 40404 40740
rect 40236 40514 40292 40526
rect 40236 40462 40238 40514
rect 40290 40462 40292 40514
rect 40124 40404 40180 40414
rect 39564 40002 39620 40012
rect 39676 40402 40180 40404
rect 39676 40350 40126 40402
rect 40178 40350 40180 40402
rect 39676 40348 40180 40350
rect 39228 39778 39284 39788
rect 38668 39006 38670 39058
rect 38722 39006 38724 39058
rect 38668 38994 38724 39006
rect 39676 38668 39732 40348
rect 40124 40338 40180 40348
rect 40236 40068 40292 40462
rect 40348 40292 40404 40684
rect 40460 40628 40516 40910
rect 40908 40964 40964 40974
rect 40964 40908 41188 40964
rect 40908 40870 40964 40908
rect 40460 40562 40516 40572
rect 40796 40852 40852 40862
rect 40460 40404 40516 40414
rect 40460 40402 40740 40404
rect 40460 40350 40462 40402
rect 40514 40350 40740 40402
rect 40460 40348 40740 40350
rect 40460 40338 40516 40348
rect 40348 40226 40404 40236
rect 39564 38612 39732 38668
rect 39900 40012 40292 40068
rect 37996 38052 38052 38062
rect 37996 38050 38164 38052
rect 37996 37998 37998 38050
rect 38050 37998 38164 38050
rect 37996 37996 38164 37998
rect 37996 37986 38052 37996
rect 37884 37202 37940 37212
rect 37996 37266 38052 37278
rect 37996 37214 37998 37266
rect 38050 37214 38052 37266
rect 37996 36932 38052 37214
rect 37884 36594 37940 36606
rect 37884 36542 37886 36594
rect 37938 36542 37940 36594
rect 37436 36482 37716 36484
rect 37436 36430 37438 36482
rect 37490 36430 37716 36482
rect 37436 36428 37716 36430
rect 37772 36484 37828 36494
rect 37436 35700 37492 36428
rect 37772 36390 37828 36428
rect 37884 36260 37940 36542
rect 37884 36194 37940 36204
rect 37996 35812 38052 36876
rect 37996 35746 38052 35756
rect 38108 36036 38164 37996
rect 37436 35634 37492 35644
rect 37548 34916 37604 34926
rect 37548 34822 37604 34860
rect 38108 34914 38164 35980
rect 38108 34862 38110 34914
rect 38162 34862 38164 34914
rect 38108 34850 38164 34862
rect 38220 37938 38276 37950
rect 38220 37886 38222 37938
rect 38274 37886 38276 37938
rect 38220 34916 38276 37886
rect 38668 37938 38724 37950
rect 38668 37886 38670 37938
rect 38722 37886 38724 37938
rect 38220 34850 38276 34860
rect 38332 36260 38388 36270
rect 37772 34692 37828 34702
rect 37772 34690 37940 34692
rect 37772 34638 37774 34690
rect 37826 34638 37940 34690
rect 37772 34636 37940 34638
rect 37772 34626 37828 34636
rect 37324 34402 37380 34412
rect 37100 33908 37156 33918
rect 37100 33570 37156 33852
rect 37100 33518 37102 33570
rect 37154 33518 37156 33570
rect 37100 33506 37156 33518
rect 36988 33124 37044 33134
rect 36988 33030 37044 33068
rect 37100 32450 37156 32462
rect 37100 32398 37102 32450
rect 37154 32398 37156 32450
rect 37100 32340 37156 32398
rect 37100 32274 37156 32284
rect 36876 31388 37156 31444
rect 37100 30996 37156 31388
rect 37100 30882 37156 30940
rect 37100 30830 37102 30882
rect 37154 30830 37156 30882
rect 37100 30818 37156 30830
rect 37212 30660 37268 34076
rect 37772 34130 37828 34142
rect 37772 34078 37774 34130
rect 37826 34078 37828 34130
rect 37548 33796 37604 33806
rect 37324 33740 37548 33796
rect 37324 33570 37380 33740
rect 37548 33730 37604 33740
rect 37324 33518 37326 33570
rect 37378 33518 37380 33570
rect 37324 33506 37380 33518
rect 37772 33348 37828 34078
rect 37884 34020 37940 34636
rect 38332 34580 38388 36204
rect 38556 35812 38612 35822
rect 38556 35698 38612 35756
rect 38556 35646 38558 35698
rect 38610 35646 38612 35698
rect 38556 35634 38612 35646
rect 38668 35140 38724 37886
rect 39452 37716 39508 37726
rect 39340 37266 39396 37278
rect 39340 37214 39342 37266
rect 39394 37214 39396 37266
rect 38780 37156 38836 37166
rect 38780 37062 38836 37100
rect 38780 35700 38836 35710
rect 38780 35606 38836 35644
rect 38220 34524 38388 34580
rect 38444 35084 38724 35140
rect 39340 35140 39396 37214
rect 37884 33954 37940 33964
rect 37996 34132 38052 34142
rect 37884 33572 37940 33582
rect 37996 33572 38052 34076
rect 38220 34018 38276 34524
rect 38220 33966 38222 34018
rect 38274 33966 38276 34018
rect 38220 33796 38276 33966
rect 38220 33730 38276 33740
rect 38332 34018 38388 34030
rect 38332 33966 38334 34018
rect 38386 33966 38388 34018
rect 38332 33572 38388 33966
rect 37884 33570 38052 33572
rect 37884 33518 37886 33570
rect 37938 33518 38052 33570
rect 37884 33516 38052 33518
rect 38108 33516 38388 33572
rect 37884 33506 37940 33516
rect 37772 33292 38052 33348
rect 37660 33234 37716 33246
rect 37660 33182 37662 33234
rect 37714 33182 37716 33234
rect 37660 32564 37716 33182
rect 37436 32338 37492 32350
rect 37436 32286 37438 32338
rect 37490 32286 37492 32338
rect 37436 31892 37492 32286
rect 37436 31826 37492 31836
rect 37324 31668 37380 31678
rect 37380 31612 37604 31668
rect 37324 31574 37380 31612
rect 37548 31218 37604 31612
rect 37660 31666 37716 32508
rect 37772 33124 37828 33134
rect 37772 32562 37828 33068
rect 37772 32510 37774 32562
rect 37826 32510 37828 32562
rect 37772 32498 37828 32510
rect 37996 32676 38052 33292
rect 37996 32562 38052 32620
rect 37996 32510 37998 32562
rect 38050 32510 38052 32562
rect 37996 32498 38052 32510
rect 37884 32452 37940 32462
rect 37884 31780 37940 32396
rect 38108 32228 38164 33516
rect 38220 33348 38276 33358
rect 38276 33292 38388 33348
rect 38220 33254 38276 33292
rect 38332 32786 38388 33292
rect 38332 32734 38334 32786
rect 38386 32734 38388 32786
rect 38332 32228 38388 32734
rect 38444 32786 38500 35084
rect 39340 35074 39396 35084
rect 38668 34468 38724 34478
rect 38668 33684 38724 34412
rect 38892 34468 38948 34478
rect 38892 34242 38948 34412
rect 39340 34244 39396 34254
rect 38892 34190 38894 34242
rect 38946 34190 38948 34242
rect 38892 34020 38948 34190
rect 39004 34188 39340 34244
rect 39004 34130 39060 34188
rect 39340 34178 39396 34188
rect 39004 34078 39006 34130
rect 39058 34078 39060 34130
rect 39004 34066 39060 34078
rect 38892 33954 38948 33964
rect 39340 33908 39396 33918
rect 39340 33814 39396 33852
rect 39452 33796 39508 37660
rect 39564 35364 39620 38612
rect 39788 38610 39844 38622
rect 39788 38558 39790 38610
rect 39842 38558 39844 38610
rect 39788 37492 39844 38558
rect 39788 37426 39844 37436
rect 39676 37380 39732 37390
rect 39676 37044 39732 37324
rect 39676 36978 39732 36988
rect 39788 37154 39844 37166
rect 39788 37102 39790 37154
rect 39842 37102 39844 37154
rect 39788 36596 39844 37102
rect 39900 37044 39956 40012
rect 40012 39844 40068 39854
rect 40012 39730 40068 39788
rect 40012 39678 40014 39730
rect 40066 39678 40068 39730
rect 40012 38948 40068 39678
rect 40460 39396 40516 39406
rect 40460 39302 40516 39340
rect 40236 38948 40292 38958
rect 40012 38946 40292 38948
rect 40012 38894 40238 38946
rect 40290 38894 40292 38946
rect 40012 38892 40292 38894
rect 40012 37938 40068 38892
rect 40236 38882 40292 38892
rect 40348 38948 40404 38958
rect 40012 37886 40014 37938
rect 40066 37886 40068 37938
rect 40012 37874 40068 37886
rect 40348 37828 40404 38892
rect 40684 38668 40740 40348
rect 40796 40402 40852 40796
rect 40796 40350 40798 40402
rect 40850 40350 40852 40402
rect 40796 39618 40852 40350
rect 40796 39566 40798 39618
rect 40850 39566 40852 39618
rect 40796 39554 40852 39566
rect 40908 40516 40964 40526
rect 40684 38612 40852 38668
rect 40348 37762 40404 37772
rect 40796 37492 40852 38612
rect 40908 37940 40964 40460
rect 41132 40402 41188 40908
rect 41244 40852 41300 45612
rect 41468 44996 41524 46398
rect 41468 44930 41524 44940
rect 41580 44772 41636 46620
rect 41692 46004 41748 46620
rect 42028 46340 42084 48190
rect 42252 48524 42364 48580
rect 42028 46274 42084 46284
rect 42140 48132 42196 48142
rect 42140 46004 42196 48076
rect 42252 46898 42308 48524
rect 42364 48514 42420 48524
rect 42252 46846 42254 46898
rect 42306 46846 42308 46898
rect 42252 46834 42308 46846
rect 42364 47234 42420 47246
rect 42364 47182 42366 47234
rect 42418 47182 42420 47234
rect 41692 45948 41972 46004
rect 41692 45780 41748 45790
rect 41692 45218 41748 45724
rect 41692 45166 41694 45218
rect 41746 45166 41748 45218
rect 41692 45154 41748 45166
rect 41356 44716 41636 44772
rect 41356 44546 41412 44716
rect 41356 44494 41358 44546
rect 41410 44494 41412 44546
rect 41356 43988 41412 44494
rect 41356 43922 41412 43932
rect 41580 44210 41636 44222
rect 41580 44158 41582 44210
rect 41634 44158 41636 44210
rect 41580 43876 41636 44158
rect 41580 43810 41636 43820
rect 41356 43652 41412 43662
rect 41580 43652 41860 43708
rect 41356 43650 41636 43652
rect 41356 43598 41358 43650
rect 41410 43598 41636 43650
rect 41356 43596 41636 43598
rect 41804 43650 41860 43652
rect 41804 43598 41806 43650
rect 41858 43598 41860 43650
rect 41356 42754 41412 43596
rect 41804 43586 41860 43598
rect 41692 43540 41748 43550
rect 41692 43446 41748 43484
rect 41916 43428 41972 45948
rect 42140 45938 42196 45948
rect 42140 45780 42196 45790
rect 42140 45778 42308 45780
rect 42140 45726 42142 45778
rect 42194 45726 42308 45778
rect 42140 45724 42308 45726
rect 42140 45714 42196 45724
rect 42140 45556 42196 45566
rect 42140 45106 42196 45500
rect 42140 45054 42142 45106
rect 42194 45054 42196 45106
rect 42140 45042 42196 45054
rect 42252 44436 42308 45724
rect 42364 44548 42420 47182
rect 42476 46676 42532 49420
rect 42588 48468 42644 50372
rect 42812 49812 42868 49822
rect 42812 49718 42868 49756
rect 42700 49252 42756 49262
rect 42700 49158 42756 49196
rect 42924 49140 42980 50372
rect 43260 49140 43316 50542
rect 43372 49812 43428 51996
rect 43484 51986 43540 51996
rect 43596 50428 43652 55916
rect 44044 56642 44100 57260
rect 44268 56644 44324 56654
rect 44044 56590 44046 56642
rect 44098 56590 44100 56642
rect 44044 55300 44100 56590
rect 43820 55244 44100 55300
rect 44156 56588 44268 56644
rect 43708 53732 43764 53742
rect 43708 53638 43764 53676
rect 43820 53508 43876 55244
rect 43932 55076 43988 55086
rect 43932 54982 43988 55020
rect 44156 54404 44212 56588
rect 44268 56578 44324 56588
rect 44268 55076 44324 55086
rect 44268 55074 44436 55076
rect 44268 55022 44270 55074
rect 44322 55022 44436 55074
rect 44268 55020 44436 55022
rect 44268 55010 44324 55020
rect 44268 54404 44324 54414
rect 44156 54402 44324 54404
rect 44156 54350 44270 54402
rect 44322 54350 44324 54402
rect 44156 54348 44324 54350
rect 44268 54338 44324 54348
rect 43708 53452 43876 53508
rect 43932 53844 43988 53854
rect 43932 53506 43988 53788
rect 44268 53732 44324 53742
rect 44268 53638 44324 53676
rect 43932 53454 43934 53506
rect 43986 53454 43988 53506
rect 43708 52500 43764 53452
rect 43932 53442 43988 53454
rect 44044 53618 44100 53630
rect 44044 53566 44046 53618
rect 44098 53566 44100 53618
rect 44044 52948 44100 53566
rect 44044 52882 44100 52892
rect 44268 52834 44324 52846
rect 44268 52782 44270 52834
rect 44322 52782 44324 52834
rect 43708 52434 43764 52444
rect 43820 52722 43876 52734
rect 43820 52670 43822 52722
rect 43874 52670 43876 52722
rect 43820 52612 43876 52670
rect 44268 52612 44324 52782
rect 43820 52556 44324 52612
rect 43708 52162 43764 52174
rect 43708 52110 43710 52162
rect 43762 52110 43764 52162
rect 43708 51604 43764 52110
rect 43708 50594 43764 51548
rect 43820 51378 43876 52556
rect 44268 52276 44324 52286
rect 44380 52276 44436 55020
rect 44492 54628 44548 58156
rect 45164 58210 45220 58222
rect 45164 58158 45166 58210
rect 45218 58158 45220 58210
rect 44716 57762 44772 57774
rect 44716 57710 44718 57762
rect 44770 57710 44772 57762
rect 44716 56532 44772 57710
rect 44940 57316 44996 57326
rect 44940 56978 44996 57260
rect 44940 56926 44942 56978
rect 44994 56926 44996 56978
rect 44940 56914 44996 56926
rect 44716 56466 44772 56476
rect 45164 56756 45220 58158
rect 45612 58212 45668 58222
rect 45612 58118 45668 58156
rect 46060 58212 46116 58222
rect 46060 58118 46116 58156
rect 47516 57874 47572 58268
rect 47516 57822 47518 57874
rect 47570 57822 47572 57874
rect 47516 57810 47572 57822
rect 47628 58210 47684 58222
rect 47628 58158 47630 58210
rect 47682 58158 47684 58210
rect 46508 57540 46564 57550
rect 46396 57538 46564 57540
rect 46396 57486 46510 57538
rect 46562 57486 46564 57538
rect 46396 57484 46564 57486
rect 45836 57428 45892 57438
rect 46172 57428 46228 57438
rect 45164 56084 45220 56700
rect 45724 57426 46228 57428
rect 45724 57374 45838 57426
rect 45890 57374 46174 57426
rect 46226 57374 46228 57426
rect 45724 57372 46228 57374
rect 45500 56642 45556 56654
rect 45500 56590 45502 56642
rect 45554 56590 45556 56642
rect 45500 56532 45556 56590
rect 44492 52612 44548 54572
rect 44604 56028 45220 56084
rect 45276 56194 45332 56206
rect 45276 56142 45278 56194
rect 45330 56142 45332 56194
rect 44604 53172 44660 56028
rect 44828 55860 44884 55870
rect 45276 55860 45332 56142
rect 44828 55858 45332 55860
rect 44828 55806 44830 55858
rect 44882 55806 45332 55858
rect 44828 55804 45332 55806
rect 44828 55794 44884 55804
rect 45052 55636 45108 55646
rect 44716 55188 44772 55198
rect 44716 54738 44772 55132
rect 44940 55076 44996 55086
rect 44716 54686 44718 54738
rect 44770 54686 44772 54738
rect 44716 54674 44772 54686
rect 44828 55074 44996 55076
rect 44828 55022 44942 55074
rect 44994 55022 44996 55074
rect 44828 55020 44996 55022
rect 44828 53956 44884 55020
rect 44940 55010 44996 55020
rect 45052 54514 45108 55580
rect 45276 55412 45332 55804
rect 45388 55412 45444 55422
rect 45276 55356 45388 55412
rect 45388 55346 45444 55356
rect 45500 55186 45556 56476
rect 45500 55134 45502 55186
rect 45554 55134 45556 55186
rect 45500 55122 45556 55134
rect 45612 56194 45668 56206
rect 45612 56142 45614 56194
rect 45666 56142 45668 56194
rect 45612 54964 45668 56142
rect 45724 55298 45780 57372
rect 45836 57362 45892 57372
rect 46172 57362 46228 57372
rect 45836 56756 45892 56766
rect 45836 56662 45892 56700
rect 46172 56644 46228 56654
rect 46172 56550 46228 56588
rect 45948 56532 46004 56542
rect 45948 56082 46004 56476
rect 45948 56030 45950 56082
rect 46002 56030 46004 56082
rect 45948 56018 46004 56030
rect 46284 55858 46340 55870
rect 46284 55806 46286 55858
rect 46338 55806 46340 55858
rect 46172 55412 46228 55422
rect 46172 55318 46228 55356
rect 45724 55246 45726 55298
rect 45778 55246 45780 55298
rect 45724 55234 45780 55246
rect 45612 54908 45892 54964
rect 45612 54628 45668 54638
rect 45388 54516 45444 54526
rect 45052 54462 45054 54514
rect 45106 54462 45108 54514
rect 45052 54450 45108 54462
rect 45276 54460 45388 54516
rect 44716 53900 44884 53956
rect 44940 54404 44996 54414
rect 44940 53954 44996 54348
rect 44940 53902 44942 53954
rect 44994 53902 44996 53954
rect 44716 53396 44772 53900
rect 44940 53890 44996 53902
rect 44828 53620 44884 53630
rect 45052 53620 45108 53630
rect 44828 53618 44996 53620
rect 44828 53566 44830 53618
rect 44882 53566 44996 53618
rect 44828 53564 44996 53566
rect 44828 53554 44884 53564
rect 44716 53330 44772 53340
rect 44604 53116 44772 53172
rect 44604 52836 44660 52846
rect 44604 52742 44660 52780
rect 44604 52612 44660 52622
rect 44492 52556 44604 52612
rect 44604 52546 44660 52556
rect 44268 52274 44436 52276
rect 44268 52222 44270 52274
rect 44322 52222 44436 52274
rect 44268 52220 44436 52222
rect 44268 52164 44324 52220
rect 43820 51326 43822 51378
rect 43874 51326 43876 51378
rect 43820 51314 43876 51326
rect 43932 52108 44324 52164
rect 43708 50542 43710 50594
rect 43762 50542 43764 50594
rect 43708 50530 43764 50542
rect 43820 51156 43876 51166
rect 43484 50372 43652 50428
rect 43484 50036 43540 50372
rect 43484 49970 43540 49980
rect 43372 49756 43540 49812
rect 43484 49700 43540 49756
rect 43596 49810 43652 49822
rect 43596 49758 43598 49810
rect 43650 49758 43652 49810
rect 43596 49700 43652 49758
rect 43484 49644 43652 49700
rect 42924 49084 43092 49140
rect 42588 48412 42980 48468
rect 42588 48244 42644 48254
rect 42588 48150 42644 48188
rect 42700 47572 42756 47582
rect 42924 47572 42980 48412
rect 43036 48356 43092 49084
rect 43148 49084 43316 49140
rect 43372 49588 43428 49598
rect 43148 48580 43204 49084
rect 43260 48916 43316 48954
rect 43260 48850 43316 48860
rect 43148 48514 43204 48524
rect 43260 48692 43316 48702
rect 43036 48300 43204 48356
rect 43036 48132 43092 48142
rect 43036 48038 43092 48076
rect 43036 47572 43092 47582
rect 42924 47570 43092 47572
rect 42924 47518 43038 47570
rect 43090 47518 43092 47570
rect 42924 47516 43092 47518
rect 42588 47348 42644 47358
rect 42588 47254 42644 47292
rect 42700 47346 42756 47516
rect 43036 47506 43092 47516
rect 42700 47294 42702 47346
rect 42754 47294 42756 47346
rect 42588 46676 42644 46686
rect 42476 46674 42644 46676
rect 42476 46622 42590 46674
rect 42642 46622 42644 46674
rect 42476 46620 42644 46622
rect 42588 46610 42644 46620
rect 42700 44884 42756 47294
rect 43148 47124 43204 48300
rect 43148 47058 43204 47068
rect 42812 47012 42868 47022
rect 42812 46786 42868 46956
rect 42812 46734 42814 46786
rect 42866 46734 42868 46786
rect 42812 46722 42868 46734
rect 43260 46900 43316 48636
rect 43372 48244 43428 49532
rect 43484 49026 43540 49038
rect 43484 48974 43486 49026
rect 43538 48974 43540 49026
rect 43484 48916 43540 48974
rect 43484 48850 43540 48860
rect 43372 48178 43428 48188
rect 43596 48132 43652 49644
rect 43484 47460 43540 47470
rect 43372 47348 43428 47358
rect 43372 47254 43428 47292
rect 43484 47346 43540 47404
rect 43484 47294 43486 47346
rect 43538 47294 43540 47346
rect 43484 47282 43540 47294
rect 43596 47346 43652 48076
rect 43820 48804 43876 51100
rect 43596 47294 43598 47346
rect 43650 47294 43652 47346
rect 43596 47282 43652 47294
rect 43708 47796 43764 47806
rect 43260 45556 43316 46844
rect 43372 46786 43428 46798
rect 43372 46734 43374 46786
rect 43426 46734 43428 46786
rect 43372 46564 43428 46734
rect 43372 46498 43428 46508
rect 43260 45490 43316 45500
rect 43260 45332 43316 45342
rect 43260 45218 43316 45276
rect 43260 45166 43262 45218
rect 43314 45166 43316 45218
rect 43260 45154 43316 45166
rect 43372 45220 43428 45230
rect 43036 45106 43092 45118
rect 43036 45054 43038 45106
rect 43090 45054 43092 45106
rect 42700 44828 42980 44884
rect 42588 44548 42644 44558
rect 42364 44546 42644 44548
rect 42364 44494 42590 44546
rect 42642 44494 42644 44546
rect 42364 44492 42644 44494
rect 42588 44482 42644 44492
rect 42700 44546 42756 44558
rect 42700 44494 42702 44546
rect 42754 44494 42756 44546
rect 42252 44380 42532 44436
rect 42476 44324 42532 44380
rect 42700 44324 42756 44494
rect 42476 44268 42756 44324
rect 41804 43372 41972 43428
rect 42140 44210 42196 44222
rect 42140 44158 42142 44210
rect 42194 44158 42196 44210
rect 41468 43316 41524 43326
rect 41468 43314 41636 43316
rect 41468 43262 41470 43314
rect 41522 43262 41636 43314
rect 41468 43260 41636 43262
rect 41468 43250 41524 43260
rect 41356 42702 41358 42754
rect 41410 42702 41412 42754
rect 41356 41972 41412 42702
rect 41580 42756 41636 43260
rect 41692 42756 41748 42766
rect 41580 42754 41748 42756
rect 41580 42702 41694 42754
rect 41746 42702 41748 42754
rect 41580 42700 41748 42702
rect 41692 42690 41748 42700
rect 41356 41906 41412 41916
rect 41468 42084 41524 42094
rect 41468 41186 41524 42028
rect 41468 41134 41470 41186
rect 41522 41134 41524 41186
rect 41468 41076 41524 41134
rect 41468 41010 41524 41020
rect 41804 40964 41860 43372
rect 42140 42756 42196 44158
rect 42812 44212 42868 44222
rect 42812 44118 42868 44156
rect 42924 43988 42980 44828
rect 42364 43932 42980 43988
rect 42252 43764 42308 43774
rect 42252 43670 42308 43708
rect 41916 42196 41972 42206
rect 41916 42102 41972 42140
rect 42028 42084 42084 42094
rect 42028 41970 42084 42028
rect 42028 41918 42030 41970
rect 42082 41918 42084 41970
rect 42028 41906 42084 41918
rect 42140 41748 42196 42700
rect 42252 43540 42308 43550
rect 42252 41970 42308 43484
rect 42252 41918 42254 41970
rect 42306 41918 42308 41970
rect 42252 41906 42308 41918
rect 42140 41692 42308 41748
rect 41804 40962 42196 40964
rect 41804 40910 41806 40962
rect 41858 40910 42196 40962
rect 41804 40908 42196 40910
rect 41804 40898 41860 40908
rect 41244 40796 41748 40852
rect 41244 40628 41300 40638
rect 41300 40572 41412 40628
rect 41244 40562 41300 40572
rect 41132 40350 41134 40402
rect 41186 40350 41188 40402
rect 41020 40290 41076 40302
rect 41020 40238 41022 40290
rect 41074 40238 41076 40290
rect 41020 38052 41076 40238
rect 41132 39508 41188 40350
rect 41356 40402 41412 40572
rect 41356 40350 41358 40402
rect 41410 40350 41412 40402
rect 41356 40292 41412 40350
rect 41356 40236 41636 40292
rect 41580 39730 41636 40236
rect 41580 39678 41582 39730
rect 41634 39678 41636 39730
rect 41580 39666 41636 39678
rect 41132 39414 41188 39452
rect 41468 39506 41524 39518
rect 41468 39454 41470 39506
rect 41522 39454 41524 39506
rect 41132 39060 41188 39070
rect 41132 38966 41188 39004
rect 41356 38948 41412 38958
rect 41356 38854 41412 38892
rect 41244 38724 41300 38762
rect 41244 38658 41300 38668
rect 41468 38276 41524 39454
rect 41580 38836 41636 38846
rect 41580 38722 41636 38780
rect 41580 38670 41582 38722
rect 41634 38670 41636 38722
rect 41580 38658 41636 38670
rect 41692 38276 41748 40796
rect 42028 40516 42084 40526
rect 42028 40404 42084 40460
rect 41916 40348 42084 40404
rect 41916 40290 41972 40348
rect 41916 40238 41918 40290
rect 41970 40238 41972 40290
rect 41916 40226 41972 40238
rect 41916 39620 41972 39630
rect 41916 39618 42084 39620
rect 41916 39566 41918 39618
rect 41970 39566 42084 39618
rect 41916 39564 42084 39566
rect 41916 39554 41972 39564
rect 42028 39172 42084 39564
rect 42028 39106 42084 39116
rect 42140 38834 42196 40908
rect 42140 38782 42142 38834
rect 42194 38782 42196 38834
rect 41804 38610 41860 38622
rect 41804 38558 41806 38610
rect 41858 38558 41860 38610
rect 41804 38500 41860 38558
rect 42140 38612 42196 38782
rect 42140 38546 42196 38556
rect 41804 38434 41860 38444
rect 42028 38388 42084 38398
rect 41692 38220 41972 38276
rect 41468 38210 41524 38220
rect 41020 37996 41300 38052
rect 40908 37884 41188 37940
rect 40908 37492 40964 37502
rect 40796 37490 40964 37492
rect 40796 37438 40910 37490
rect 40962 37438 40964 37490
rect 40796 37436 40964 37438
rect 40908 37426 40964 37436
rect 41132 37490 41188 37884
rect 41132 37438 41134 37490
rect 41186 37438 41188 37490
rect 41132 37426 41188 37438
rect 40348 37266 40404 37278
rect 40348 37214 40350 37266
rect 40402 37214 40404 37266
rect 40348 37156 40404 37214
rect 41020 37268 41076 37278
rect 41020 37174 41076 37212
rect 40348 37090 40404 37100
rect 41132 37156 41188 37166
rect 39900 36988 40292 37044
rect 39788 36530 39844 36540
rect 39900 36482 39956 36494
rect 39900 36430 39902 36482
rect 39954 36430 39956 36482
rect 39564 35298 39620 35308
rect 39676 36370 39732 36382
rect 39676 36318 39678 36370
rect 39730 36318 39732 36370
rect 39564 34916 39620 34926
rect 39564 34822 39620 34860
rect 39676 34244 39732 36318
rect 39788 36372 39844 36382
rect 39788 35812 39844 36316
rect 39900 35924 39956 36430
rect 39900 35858 39956 35868
rect 40124 36148 40180 36158
rect 40124 35922 40180 36092
rect 40124 35870 40126 35922
rect 40178 35870 40180 35922
rect 39788 35718 39844 35756
rect 40012 35810 40068 35822
rect 40012 35758 40014 35810
rect 40066 35758 40068 35810
rect 39900 35364 39956 35374
rect 39788 35308 39900 35364
rect 39788 34580 39844 35308
rect 39900 35298 39956 35308
rect 40012 35140 40068 35758
rect 40124 35364 40180 35870
rect 40236 35922 40292 36988
rect 41020 36820 41076 36830
rect 40796 36764 41020 36820
rect 40236 35870 40238 35922
rect 40290 35870 40292 35922
rect 40236 35858 40292 35870
rect 40684 35924 40740 35934
rect 40348 35812 40404 35822
rect 40348 35718 40404 35756
rect 40124 35298 40180 35308
rect 40572 35140 40628 35150
rect 40684 35140 40740 35868
rect 40012 35084 40404 35140
rect 40012 34916 40068 34926
rect 39788 34524 39956 34580
rect 39900 34468 39956 34524
rect 39788 34244 39844 34254
rect 39676 34188 39788 34244
rect 39676 34130 39732 34188
rect 39788 34178 39844 34188
rect 39676 34078 39678 34130
rect 39730 34078 39732 34130
rect 39676 34066 39732 34078
rect 39900 34130 39956 34412
rect 39900 34078 39902 34130
rect 39954 34078 39956 34130
rect 39900 34066 39956 34078
rect 40012 34020 40068 34860
rect 40348 34804 40404 35084
rect 40628 35084 40740 35140
rect 40572 35046 40628 35084
rect 40572 34804 40628 34814
rect 40348 34802 40628 34804
rect 40348 34750 40574 34802
rect 40626 34750 40628 34802
rect 40348 34748 40628 34750
rect 40348 34356 40404 34366
rect 40348 34262 40404 34300
rect 40012 33954 40068 33964
rect 40348 33908 40404 33918
rect 39452 33740 39620 33796
rect 38668 33618 38724 33628
rect 39452 33572 39508 33582
rect 38444 32734 38446 32786
rect 38498 32734 38500 32786
rect 38444 32722 38500 32734
rect 38780 32788 38836 32798
rect 38780 32694 38836 32732
rect 38556 32676 38612 32686
rect 38556 32582 38612 32620
rect 39452 32564 39508 33516
rect 39452 32470 39508 32508
rect 39228 32452 39284 32462
rect 39228 32358 39284 32396
rect 38108 32172 38276 32228
rect 38332 32172 38612 32228
rect 38220 32116 38276 32172
rect 38220 32060 38388 32116
rect 37996 31780 38052 31790
rect 37884 31778 38052 31780
rect 37884 31726 37998 31778
rect 38050 31726 38052 31778
rect 37884 31724 38052 31726
rect 37996 31714 38052 31724
rect 38220 31778 38276 31790
rect 38220 31726 38222 31778
rect 38274 31726 38276 31778
rect 37660 31614 37662 31666
rect 37714 31614 37716 31666
rect 37660 31556 37716 31614
rect 38220 31556 38276 31726
rect 37660 31500 38276 31556
rect 38332 31556 38388 32060
rect 38556 31948 38612 32172
rect 38556 31892 38724 31948
rect 38556 31780 38612 31790
rect 38556 31686 38612 31724
rect 38668 31668 38724 31892
rect 38892 31668 38948 31678
rect 38668 31666 38948 31668
rect 38668 31614 38894 31666
rect 38946 31614 38948 31666
rect 38668 31612 38948 31614
rect 38892 31602 38948 31612
rect 38332 31490 38388 31500
rect 37548 31166 37550 31218
rect 37602 31166 37604 31218
rect 37548 31154 37604 31166
rect 38780 31220 38836 31230
rect 37660 31108 37716 31118
rect 38780 31108 38836 31164
rect 37100 30604 37268 30660
rect 37324 30660 37380 30670
rect 36876 29426 36932 29438
rect 36876 29374 36878 29426
rect 36930 29374 36932 29426
rect 36876 29316 36932 29374
rect 36876 29250 36932 29260
rect 36428 28814 36430 28866
rect 36482 28814 36484 28866
rect 36428 28802 36484 28814
rect 36540 29148 36820 29204
rect 36428 28308 36484 28318
rect 36428 27858 36484 28252
rect 36428 27806 36430 27858
rect 36482 27806 36484 27858
rect 36428 27794 36484 27806
rect 36540 27636 36596 29148
rect 36988 29092 37044 29102
rect 36652 28980 36708 28990
rect 36652 28082 36708 28924
rect 36988 28644 37044 29036
rect 36988 28550 37044 28588
rect 37100 28420 37156 30604
rect 37212 30210 37268 30222
rect 37212 30158 37214 30210
rect 37266 30158 37268 30210
rect 37212 29988 37268 30158
rect 37212 29922 37268 29932
rect 37212 29428 37268 29438
rect 37212 29334 37268 29372
rect 37212 28868 37268 28878
rect 37212 28754 37268 28812
rect 37324 28866 37380 30604
rect 37660 30210 37716 31052
rect 38444 31106 38836 31108
rect 38444 31054 38782 31106
rect 38834 31054 38836 31106
rect 38444 31052 38836 31054
rect 38108 30996 38164 31006
rect 37660 30158 37662 30210
rect 37714 30158 37716 30210
rect 37660 30146 37716 30158
rect 37772 30884 37828 30894
rect 37324 28814 37326 28866
rect 37378 28814 37380 28866
rect 37324 28802 37380 28814
rect 37436 29988 37492 29998
rect 37212 28702 37214 28754
rect 37266 28702 37268 28754
rect 37212 28690 37268 28702
rect 36652 28030 36654 28082
rect 36706 28030 36708 28082
rect 36652 28018 36708 28030
rect 36988 28364 37156 28420
rect 36316 27134 36318 27186
rect 36370 27134 36372 27186
rect 36316 26852 36372 27134
rect 36316 26786 36372 26796
rect 36428 27580 36596 27636
rect 36764 27860 36820 27870
rect 36764 27634 36820 27804
rect 36764 27582 36766 27634
rect 36818 27582 36820 27634
rect 36316 26402 36372 26414
rect 36316 26350 36318 26402
rect 36370 26350 36372 26402
rect 36316 24834 36372 26350
rect 36316 24782 36318 24834
rect 36370 24782 36372 24834
rect 36316 22372 36372 24782
rect 36428 22372 36484 27580
rect 36764 26404 36820 27582
rect 36988 26908 37044 28364
rect 37324 27858 37380 27870
rect 37324 27806 37326 27858
rect 37378 27806 37380 27858
rect 37100 27748 37156 27758
rect 37100 27186 37156 27692
rect 37100 27134 37102 27186
rect 37154 27134 37156 27186
rect 37100 27122 37156 27134
rect 37212 27636 37268 27646
rect 37212 27076 37268 27580
rect 37212 27010 37268 27020
rect 36988 26852 37156 26908
rect 36540 26348 36820 26404
rect 36540 24388 36596 26348
rect 36988 25508 37044 25518
rect 36988 25414 37044 25452
rect 36540 22596 36596 24332
rect 36652 24724 36708 24734
rect 36652 23380 36708 24668
rect 36988 23716 37044 23726
rect 36988 23622 37044 23660
rect 37100 23604 37156 26852
rect 37324 26852 37380 27806
rect 37324 26786 37380 26796
rect 37436 26292 37492 29932
rect 37772 28754 37828 30828
rect 37996 30212 38052 30222
rect 37996 29986 38052 30156
rect 37996 29934 37998 29986
rect 38050 29934 38052 29986
rect 37996 29652 38052 29934
rect 37996 29586 38052 29596
rect 38108 29538 38164 30940
rect 38444 29650 38500 31052
rect 38780 31042 38836 31052
rect 39340 30324 39396 30334
rect 39564 30324 39620 33740
rect 39676 33346 39732 33358
rect 40124 33348 40180 33358
rect 39676 33294 39678 33346
rect 39730 33294 39732 33346
rect 39676 32676 39732 33294
rect 39788 33346 40180 33348
rect 39788 33294 40126 33346
rect 40178 33294 40180 33346
rect 39788 33292 40180 33294
rect 39788 32788 39844 33292
rect 40124 33282 40180 33292
rect 40348 33236 40404 33852
rect 40572 33570 40628 34748
rect 40796 34356 40852 36764
rect 41020 36754 41076 36764
rect 41020 36484 41076 36494
rect 40908 36372 40964 36382
rect 40908 36278 40964 36316
rect 41020 36036 41076 36428
rect 40572 33518 40574 33570
rect 40626 33518 40628 33570
rect 40572 33506 40628 33518
rect 40684 34300 40852 34356
rect 40908 35698 40964 35710
rect 40908 35646 40910 35698
rect 40962 35646 40964 35698
rect 40684 33348 40740 34300
rect 40908 34244 40964 35646
rect 41020 34914 41076 35980
rect 41020 34862 41022 34914
rect 41074 34862 41076 34914
rect 41020 34850 41076 34862
rect 41132 35810 41188 37100
rect 41244 36596 41300 37996
rect 41692 38050 41748 38062
rect 41692 37998 41694 38050
rect 41746 37998 41748 38050
rect 41468 37492 41524 37502
rect 41524 37436 41636 37492
rect 41468 37426 41524 37436
rect 41356 37378 41412 37390
rect 41356 37326 41358 37378
rect 41410 37326 41412 37378
rect 41356 36820 41412 37326
rect 41356 36754 41412 36764
rect 41244 36540 41412 36596
rect 41132 35758 41134 35810
rect 41186 35758 41188 35810
rect 41132 34692 41188 35758
rect 41132 34626 41188 34636
rect 41244 34468 41300 34478
rect 40908 34178 40964 34188
rect 41020 34242 41076 34254
rect 41020 34190 41022 34242
rect 41074 34190 41076 34242
rect 40796 34132 40852 34142
rect 40796 34038 40852 34076
rect 41020 33572 41076 34190
rect 41132 34130 41188 34142
rect 41132 34078 41134 34130
rect 41186 34078 41188 34130
rect 41132 33908 41188 34078
rect 41132 33842 41188 33852
rect 41020 33506 41076 33516
rect 40348 33170 40404 33180
rect 40460 33292 40740 33348
rect 40236 32788 40292 32798
rect 39788 32694 39844 32732
rect 40012 32786 40292 32788
rect 40012 32734 40238 32786
rect 40290 32734 40292 32786
rect 40012 32732 40292 32734
rect 39676 32340 39732 32620
rect 39676 32284 39844 32340
rect 39676 31892 39732 31902
rect 39676 31778 39732 31836
rect 39676 31726 39678 31778
rect 39730 31726 39732 31778
rect 39676 31218 39732 31726
rect 39676 31166 39678 31218
rect 39730 31166 39732 31218
rect 39676 31154 39732 31166
rect 39788 30884 39844 32284
rect 40012 31220 40068 32732
rect 40236 32722 40292 32732
rect 40460 32786 40516 33292
rect 40460 32734 40462 32786
rect 40514 32734 40516 32786
rect 40460 32722 40516 32734
rect 41132 33124 41188 33134
rect 40012 31154 40068 31164
rect 40124 32564 40180 32574
rect 40124 31108 40180 32508
rect 40684 31780 40740 31818
rect 40684 31714 40740 31724
rect 41132 31666 41188 33068
rect 41132 31614 41134 31666
rect 41186 31614 41188 31666
rect 41132 31602 41188 31614
rect 40124 31042 40180 31052
rect 40124 30884 40180 30894
rect 39788 30882 40180 30884
rect 39788 30830 40126 30882
rect 40178 30830 40180 30882
rect 39788 30828 40180 30830
rect 40124 30818 40180 30828
rect 40908 30884 40964 30894
rect 40908 30790 40964 30828
rect 41244 30772 41300 34412
rect 41356 34356 41412 36540
rect 41468 36484 41524 36494
rect 41580 36484 41636 37436
rect 41692 37156 41748 37998
rect 41692 37090 41748 37100
rect 41916 37378 41972 38220
rect 41916 37326 41918 37378
rect 41970 37326 41972 37378
rect 41468 36482 41636 36484
rect 41468 36430 41470 36482
rect 41522 36430 41636 36482
rect 41468 36428 41636 36430
rect 41692 36932 41748 36942
rect 41468 36418 41524 36428
rect 41468 35588 41524 35598
rect 41468 35494 41524 35532
rect 41580 34916 41636 34926
rect 41468 34356 41524 34366
rect 41356 34354 41524 34356
rect 41356 34302 41470 34354
rect 41522 34302 41524 34354
rect 41356 34300 41524 34302
rect 41468 34290 41524 34300
rect 41356 34020 41412 34030
rect 41356 33346 41412 33964
rect 41580 33908 41636 34860
rect 41580 33842 41636 33852
rect 41692 34354 41748 36876
rect 41916 35140 41972 37326
rect 42028 37042 42084 38332
rect 42140 38052 42196 38062
rect 42140 37378 42196 37996
rect 42140 37326 42142 37378
rect 42194 37326 42196 37378
rect 42140 37314 42196 37326
rect 42028 36990 42030 37042
rect 42082 36990 42084 37042
rect 42028 36978 42084 36990
rect 42028 36484 42084 36494
rect 42028 36390 42084 36428
rect 42028 35698 42084 35710
rect 42028 35646 42030 35698
rect 42082 35646 42084 35698
rect 42028 35364 42084 35646
rect 42252 35588 42308 41692
rect 42364 38668 42420 43932
rect 42924 43540 42980 43550
rect 42924 43446 42980 43484
rect 42588 43426 42644 43438
rect 42588 43374 42590 43426
rect 42642 43374 42644 43426
rect 42588 42980 42644 43374
rect 42588 42924 42980 42980
rect 42812 42756 42868 42766
rect 42588 42754 42868 42756
rect 42588 42702 42814 42754
rect 42866 42702 42868 42754
rect 42588 42700 42868 42702
rect 42476 42530 42532 42542
rect 42476 42478 42478 42530
rect 42530 42478 42532 42530
rect 42476 41524 42532 42478
rect 42588 42194 42644 42700
rect 42812 42690 42868 42700
rect 42588 42142 42590 42194
rect 42642 42142 42644 42194
rect 42588 42130 42644 42142
rect 42924 42196 42980 42924
rect 42924 42082 42980 42140
rect 42924 42030 42926 42082
rect 42978 42030 42980 42082
rect 42924 42018 42980 42030
rect 42700 41972 42756 41982
rect 42700 41878 42756 41916
rect 42476 41468 42756 41524
rect 42588 41074 42644 41086
rect 42588 41022 42590 41074
rect 42642 41022 42644 41074
rect 42476 40852 42532 40862
rect 42476 40514 42532 40796
rect 42476 40462 42478 40514
rect 42530 40462 42532 40514
rect 42476 40450 42532 40462
rect 42588 40292 42644 41022
rect 42700 40514 42756 41468
rect 43036 40852 43092 45054
rect 43148 44996 43204 45006
rect 43148 44902 43204 44940
rect 43372 44546 43428 45164
rect 43708 45106 43764 47740
rect 43820 47684 43876 48748
rect 43820 47458 43876 47628
rect 43820 47406 43822 47458
rect 43874 47406 43876 47458
rect 43820 47394 43876 47406
rect 43820 46900 43876 46910
rect 43932 46900 43988 52108
rect 44604 52052 44660 52062
rect 44604 51490 44660 51996
rect 44716 51602 44772 53116
rect 44716 51550 44718 51602
rect 44770 51550 44772 51602
rect 44716 51538 44772 51550
rect 44828 51938 44884 51950
rect 44828 51886 44830 51938
rect 44882 51886 44884 51938
rect 44604 51438 44606 51490
rect 44658 51438 44660 51490
rect 44268 51268 44324 51278
rect 44268 51266 44436 51268
rect 44268 51214 44270 51266
rect 44322 51214 44436 51266
rect 44268 51212 44436 51214
rect 44268 51202 44324 51212
rect 44268 50594 44324 50606
rect 44268 50542 44270 50594
rect 44322 50542 44324 50594
rect 44268 50372 44324 50542
rect 44268 50306 44324 50316
rect 44380 50484 44436 51212
rect 44156 49586 44212 49598
rect 44156 49534 44158 49586
rect 44210 49534 44212 49586
rect 44044 49140 44100 49150
rect 44044 49046 44100 49084
rect 44156 48354 44212 49534
rect 44156 48302 44158 48354
rect 44210 48302 44212 48354
rect 44156 47460 44212 48302
rect 44380 48244 44436 50428
rect 44492 50932 44548 50942
rect 44492 48468 44548 50876
rect 44604 48580 44660 51438
rect 44828 49810 44884 51886
rect 44940 51602 44996 53564
rect 45052 53526 45108 53564
rect 45276 53058 45332 54460
rect 45388 54450 45444 54460
rect 45612 54404 45668 54572
rect 45724 54516 45780 54526
rect 45724 54422 45780 54460
rect 45612 54338 45668 54348
rect 45388 53844 45444 53854
rect 45388 53750 45444 53788
rect 45612 53732 45668 53742
rect 45500 53730 45668 53732
rect 45500 53678 45614 53730
rect 45666 53678 45668 53730
rect 45500 53676 45668 53678
rect 45500 53170 45556 53676
rect 45612 53666 45668 53676
rect 45836 53732 45892 54908
rect 46284 54852 46340 55806
rect 46396 54964 46452 57484
rect 46508 57474 46564 57484
rect 47068 57538 47124 57550
rect 47068 57486 47070 57538
rect 47122 57486 47124 57538
rect 46620 57428 46676 57438
rect 46508 56756 46564 56766
rect 46508 56662 46564 56700
rect 46620 55636 46676 57372
rect 46732 57426 46788 57438
rect 46732 57374 46734 57426
rect 46786 57374 46788 57426
rect 46732 56306 46788 57374
rect 47068 57316 47124 57486
rect 47068 57250 47124 57260
rect 47628 57540 47684 58158
rect 47628 57204 47684 57484
rect 46732 56254 46734 56306
rect 46786 56254 46788 56306
rect 46732 56242 46788 56254
rect 47516 57148 47684 57204
rect 47068 56196 47124 56206
rect 46956 56194 47124 56196
rect 46956 56142 47070 56194
rect 47122 56142 47124 56194
rect 46956 56140 47124 56142
rect 46844 55972 46900 55982
rect 46620 55570 46676 55580
rect 46732 55916 46844 55972
rect 46508 55188 46564 55198
rect 46508 55094 46564 55132
rect 46396 54898 46452 54908
rect 46284 54786 46340 54796
rect 46284 54514 46340 54526
rect 46284 54462 46286 54514
rect 46338 54462 46340 54514
rect 46284 54404 46340 54462
rect 46620 54516 46676 54526
rect 46732 54516 46788 55916
rect 46844 55906 46900 55916
rect 46676 54460 46788 54516
rect 46956 54514 47012 56140
rect 47068 56130 47124 56140
rect 47180 55076 47236 55086
rect 47180 54982 47236 55020
rect 47404 55076 47460 55086
rect 47404 54982 47460 55020
rect 47516 54852 47572 57148
rect 47628 56756 47684 56766
rect 47740 56756 47796 59948
rect 47964 59938 48020 59948
rect 48412 59444 48468 63200
rect 48972 60228 49028 60238
rect 48972 60134 49028 60172
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 48412 59378 48468 59388
rect 49756 59444 49812 59454
rect 49756 59350 49812 59388
rect 62188 59330 62244 59342
rect 62188 59278 62190 59330
rect 62242 59278 62244 59330
rect 48748 59220 48804 59230
rect 48188 59218 48804 59220
rect 48188 59166 48750 59218
rect 48802 59166 48804 59218
rect 48188 59164 48804 59166
rect 48076 58548 48132 58558
rect 48076 58210 48132 58492
rect 48076 58158 48078 58210
rect 48130 58158 48132 58210
rect 48076 57764 48132 58158
rect 48188 57874 48244 59164
rect 48748 59154 48804 59164
rect 52108 58548 52164 58558
rect 52108 58454 52164 58492
rect 52780 58548 52836 58558
rect 62188 58548 62244 59278
rect 52780 58546 52948 58548
rect 52780 58494 52782 58546
rect 52834 58494 52948 58546
rect 52780 58492 52948 58494
rect 52780 58482 52836 58492
rect 51324 58436 51380 58446
rect 51324 58342 51380 58380
rect 50764 58324 50820 58334
rect 50764 58230 50820 58268
rect 51548 58324 51604 58334
rect 48524 58212 48580 58222
rect 48524 58118 48580 58156
rect 48972 58210 49028 58222
rect 48972 58158 48974 58210
rect 49026 58158 49028 58210
rect 48972 58100 49028 58158
rect 48972 58034 49028 58044
rect 49196 58212 49252 58222
rect 48188 57822 48190 57874
rect 48242 57822 48244 57874
rect 48188 57810 48244 57822
rect 48412 57988 48468 57998
rect 48076 57698 48132 57708
rect 47964 57652 48020 57662
rect 47964 57558 48020 57596
rect 47684 56700 47796 56756
rect 47628 56662 47684 56700
rect 48076 56306 48132 56318
rect 48076 56254 48078 56306
rect 48130 56254 48132 56306
rect 48076 56196 48132 56254
rect 48076 56130 48132 56140
rect 48188 56084 48244 56094
rect 48188 55990 48244 56028
rect 47628 55970 47684 55982
rect 47628 55918 47630 55970
rect 47682 55918 47684 55970
rect 47628 55748 47684 55918
rect 47628 55682 47684 55692
rect 47740 55412 47796 55422
rect 47740 55318 47796 55356
rect 47964 55300 48020 55310
rect 47516 54796 47796 54852
rect 47068 54740 47124 54750
rect 47068 54738 47460 54740
rect 47068 54686 47070 54738
rect 47122 54686 47460 54738
rect 47068 54684 47460 54686
rect 47068 54674 47124 54684
rect 47404 54626 47460 54684
rect 47404 54574 47406 54626
rect 47458 54574 47460 54626
rect 47404 54562 47460 54574
rect 47628 54626 47684 54638
rect 47628 54574 47630 54626
rect 47682 54574 47684 54626
rect 46956 54462 46958 54514
rect 47010 54462 47012 54514
rect 46620 54422 46676 54460
rect 46284 54338 46340 54348
rect 46844 54290 46900 54302
rect 46844 54238 46846 54290
rect 46898 54238 46900 54290
rect 46620 54180 46676 54190
rect 45836 53666 45892 53676
rect 46508 53732 46564 53742
rect 45500 53118 45502 53170
rect 45554 53118 45556 53170
rect 45500 53106 45556 53118
rect 45724 53620 45780 53630
rect 45276 53006 45278 53058
rect 45330 53006 45332 53058
rect 45276 52994 45332 53006
rect 45052 52946 45108 52958
rect 45052 52894 45054 52946
rect 45106 52894 45108 52946
rect 45052 52612 45108 52894
rect 45052 52546 45108 52556
rect 45388 52836 45444 52846
rect 45388 52274 45444 52780
rect 45612 52724 45668 52734
rect 45724 52724 45780 53564
rect 46508 53618 46564 53676
rect 46508 53566 46510 53618
rect 46562 53566 46564 53618
rect 46508 53554 46564 53566
rect 46060 53508 46116 53518
rect 45836 53060 45892 53070
rect 45836 52946 45892 53004
rect 45836 52894 45838 52946
rect 45890 52894 45892 52946
rect 45836 52882 45892 52894
rect 46060 52946 46116 53452
rect 46508 53396 46564 53406
rect 46396 53172 46452 53182
rect 46396 53078 46452 53116
rect 46060 52894 46062 52946
rect 46114 52894 46116 52946
rect 46060 52882 46116 52894
rect 46508 53058 46564 53340
rect 46508 53006 46510 53058
rect 46562 53006 46564 53058
rect 46508 52948 46564 53006
rect 46508 52882 46564 52892
rect 45612 52722 45780 52724
rect 45612 52670 45614 52722
rect 45666 52670 45780 52722
rect 45612 52668 45780 52670
rect 45612 52658 45668 52668
rect 45388 52222 45390 52274
rect 45442 52222 45444 52274
rect 45164 52164 45220 52174
rect 45164 52070 45220 52108
rect 44940 51550 44942 51602
rect 44994 51550 44996 51602
rect 44940 51538 44996 51550
rect 44828 49758 44830 49810
rect 44882 49758 44884 49810
rect 44828 49746 44884 49758
rect 45052 50482 45108 50494
rect 45052 50430 45054 50482
rect 45106 50430 45108 50482
rect 45052 50372 45108 50430
rect 45052 48916 45108 50316
rect 45052 48850 45108 48860
rect 45164 50370 45220 50382
rect 45164 50318 45166 50370
rect 45218 50318 45220 50370
rect 44940 48802 44996 48814
rect 44940 48750 44942 48802
rect 44994 48750 44996 48802
rect 44604 48524 44884 48580
rect 44492 48412 44772 48468
rect 44604 48244 44660 48254
rect 44380 48188 44604 48244
rect 44604 48150 44660 48188
rect 44156 47394 44212 47404
rect 44716 47348 44772 48412
rect 44828 47572 44884 48524
rect 44828 47506 44884 47516
rect 44380 47292 44772 47348
rect 44268 47236 44324 47246
rect 44268 47142 44324 47180
rect 43820 46898 43988 46900
rect 43820 46846 43822 46898
rect 43874 46846 43988 46898
rect 43820 46844 43988 46846
rect 44044 46900 44100 46910
rect 43820 45780 43876 46844
rect 44044 46806 44100 46844
rect 44380 46674 44436 47292
rect 44828 47236 44884 47246
rect 44380 46622 44382 46674
rect 44434 46622 44436 46674
rect 43820 45714 43876 45724
rect 43932 46562 43988 46574
rect 43932 46510 43934 46562
rect 43986 46510 43988 46562
rect 43932 45444 43988 46510
rect 44268 46002 44324 46014
rect 44268 45950 44270 46002
rect 44322 45950 44324 46002
rect 44268 45668 44324 45950
rect 44268 45602 44324 45612
rect 44380 45556 44436 46622
rect 44380 45490 44436 45500
rect 44492 47234 44884 47236
rect 44492 47182 44830 47234
rect 44882 47182 44884 47234
rect 44492 47180 44884 47182
rect 43932 45378 43988 45388
rect 44492 45332 44548 47180
rect 44828 47170 44884 47180
rect 44828 46676 44884 46686
rect 44828 46582 44884 46620
rect 44940 46564 44996 48750
rect 45164 48356 45220 50318
rect 45164 48290 45220 48300
rect 45276 48914 45332 48926
rect 45276 48862 45278 48914
rect 45330 48862 45332 48914
rect 44940 46498 44996 46508
rect 45164 47234 45220 47246
rect 45164 47182 45166 47234
rect 45218 47182 45220 47234
rect 44940 46340 44996 46350
rect 44940 46004 44996 46284
rect 45164 46116 45220 47182
rect 45164 46050 45220 46060
rect 44940 45910 44996 45948
rect 44156 45276 44548 45332
rect 44828 45668 44884 45678
rect 45276 45668 45332 48862
rect 45388 48916 45444 52222
rect 45948 52388 46004 52398
rect 45724 52162 45780 52174
rect 45724 52110 45726 52162
rect 45778 52110 45780 52162
rect 45724 50484 45780 52110
rect 45836 52164 45892 52174
rect 45836 51602 45892 52108
rect 45948 52164 46004 52332
rect 45948 52162 46116 52164
rect 45948 52110 45950 52162
rect 46002 52110 46116 52162
rect 45948 52108 46116 52110
rect 45948 52098 46004 52108
rect 45836 51550 45838 51602
rect 45890 51550 45892 51602
rect 45836 51538 45892 51550
rect 45948 50594 46004 50606
rect 45948 50542 45950 50594
rect 46002 50542 46004 50594
rect 45724 50418 45780 50428
rect 45836 50482 45892 50494
rect 45836 50430 45838 50482
rect 45890 50430 45892 50482
rect 45500 50036 45556 50046
rect 45500 49698 45556 49980
rect 45500 49646 45502 49698
rect 45554 49646 45556 49698
rect 45500 49140 45556 49646
rect 45724 49810 45780 49822
rect 45724 49758 45726 49810
rect 45778 49758 45780 49810
rect 45724 49140 45780 49758
rect 45836 49364 45892 50430
rect 45948 49364 46004 50542
rect 46060 49588 46116 52108
rect 46060 49522 46116 49532
rect 46284 51938 46340 51950
rect 46284 51886 46286 51938
rect 46338 51886 46340 51938
rect 45948 49308 46116 49364
rect 45836 49298 45892 49308
rect 45948 49140 46004 49150
rect 45724 49138 46004 49140
rect 45724 49086 45950 49138
rect 46002 49086 46004 49138
rect 45724 49084 46004 49086
rect 45500 49074 45556 49084
rect 45948 49028 46004 49084
rect 45948 48962 46004 48972
rect 45724 48916 45780 48926
rect 45388 48914 45892 48916
rect 45388 48862 45726 48914
rect 45778 48862 45892 48914
rect 45388 48860 45892 48862
rect 45724 48850 45780 48860
rect 45388 48244 45444 48254
rect 45388 46786 45444 48188
rect 45500 48242 45556 48254
rect 45500 48190 45502 48242
rect 45554 48190 45556 48242
rect 45500 48132 45556 48190
rect 45500 48066 45556 48076
rect 45612 48130 45668 48142
rect 45612 48078 45614 48130
rect 45666 48078 45668 48130
rect 45612 47684 45668 48078
rect 45612 47012 45668 47628
rect 45388 46734 45390 46786
rect 45442 46734 45444 46786
rect 45388 46722 45444 46734
rect 45500 46956 45668 47012
rect 45724 47460 45780 47470
rect 45388 45780 45444 45790
rect 45388 45686 45444 45724
rect 44884 45612 45332 45668
rect 43820 45220 43876 45258
rect 43820 45154 43876 45164
rect 43932 45220 43988 45230
rect 44156 45220 44212 45276
rect 43932 45218 44212 45220
rect 43932 45166 43934 45218
rect 43986 45166 44212 45218
rect 43932 45164 44212 45166
rect 43932 45154 43988 45164
rect 43708 45054 43710 45106
rect 43762 45054 43764 45106
rect 43708 44772 43764 45054
rect 43708 44716 44100 44772
rect 43372 44494 43374 44546
rect 43426 44494 43428 44546
rect 43372 44482 43428 44494
rect 43708 44548 43764 44558
rect 43932 44548 43988 44558
rect 43764 44492 43876 44548
rect 43708 44482 43764 44492
rect 43148 44324 43204 44334
rect 43148 44230 43204 44268
rect 43820 44322 43876 44492
rect 43932 44454 43988 44492
rect 43820 44270 43822 44322
rect 43874 44270 43876 44322
rect 43820 44258 43876 44270
rect 44044 43764 44100 44716
rect 43932 43708 44100 43764
rect 43484 43652 43540 43662
rect 43484 42642 43540 43596
rect 43820 43652 43876 43662
rect 43932 43652 43988 43708
rect 43876 43596 43988 43652
rect 43820 43558 43876 43596
rect 43596 43540 43652 43550
rect 43596 42754 43652 43484
rect 44156 43540 44212 45164
rect 44492 45108 44548 45118
rect 44156 43446 44212 43484
rect 44268 44882 44324 44894
rect 44268 44830 44270 44882
rect 44322 44830 44324 44882
rect 44268 43764 44324 44830
rect 44268 43538 44324 43708
rect 44268 43486 44270 43538
rect 44322 43486 44324 43538
rect 44268 43474 44324 43486
rect 44380 44212 44436 44222
rect 44380 43538 44436 44156
rect 44492 43764 44548 45052
rect 44716 44996 44772 45006
rect 44716 44322 44772 44940
rect 44716 44270 44718 44322
rect 44770 44270 44772 44322
rect 44716 44258 44772 44270
rect 44828 43876 44884 45612
rect 45164 45220 45220 45230
rect 44940 44324 44996 44334
rect 44940 44230 44996 44268
rect 45164 44322 45220 45164
rect 45164 44270 45166 44322
rect 45218 44270 45220 44322
rect 45164 44258 45220 44270
rect 44828 43810 44884 43820
rect 45388 44212 45444 44222
rect 44492 43708 44660 43764
rect 44380 43486 44382 43538
rect 44434 43486 44436 43538
rect 43596 42702 43598 42754
rect 43650 42702 43652 42754
rect 43596 42690 43652 42702
rect 43932 43426 43988 43438
rect 43932 43374 43934 43426
rect 43986 43374 43988 43426
rect 43484 42590 43486 42642
rect 43538 42590 43540 42642
rect 43484 42578 43540 42590
rect 43708 42196 43764 42206
rect 43260 41972 43316 41982
rect 43260 41878 43316 41916
rect 43708 41970 43764 42140
rect 43708 41918 43710 41970
rect 43762 41918 43764 41970
rect 43708 41906 43764 41918
rect 43932 41972 43988 43374
rect 44380 43204 44436 43486
rect 44156 43148 44436 43204
rect 44156 42866 44212 43148
rect 44604 43092 44660 43708
rect 45276 43652 45332 43662
rect 44268 43036 44660 43092
rect 44716 43650 45332 43652
rect 44716 43598 45278 43650
rect 45330 43598 45332 43650
rect 44716 43596 45332 43598
rect 44268 42978 44324 43036
rect 44268 42926 44270 42978
rect 44322 42926 44324 42978
rect 44268 42914 44324 42926
rect 44156 42814 44158 42866
rect 44210 42814 44212 42866
rect 44156 42802 44212 42814
rect 44380 42644 44436 42654
rect 44268 42588 44380 42644
rect 44156 41972 44212 41982
rect 43932 41970 44212 41972
rect 43932 41918 44158 41970
rect 44210 41918 44212 41970
rect 43932 41916 44212 41918
rect 44156 41906 44212 41916
rect 44268 40852 44324 42588
rect 44380 42578 44436 42588
rect 44716 42308 44772 43596
rect 45276 43586 45332 43596
rect 45388 43428 45444 44156
rect 45276 43372 45444 43428
rect 45276 42754 45332 43372
rect 45276 42702 45278 42754
rect 45330 42702 45332 42754
rect 44492 42252 44772 42308
rect 45052 42642 45108 42654
rect 45052 42590 45054 42642
rect 45106 42590 45108 42642
rect 45052 42532 45108 42590
rect 44380 42196 44436 42206
rect 44380 42102 44436 42140
rect 44492 41858 44548 42252
rect 44492 41806 44494 41858
rect 44546 41806 44548 41858
rect 44492 41794 44548 41806
rect 44940 42084 44996 42094
rect 44380 41412 44436 41422
rect 44940 41412 44996 42028
rect 44380 41410 44996 41412
rect 44380 41358 44382 41410
rect 44434 41358 44996 41410
rect 44380 41356 44996 41358
rect 44380 41346 44436 41356
rect 44940 41074 44996 41356
rect 44940 41022 44942 41074
rect 44994 41022 44996 41074
rect 44940 41010 44996 41022
rect 42700 40462 42702 40514
rect 42754 40462 42756 40514
rect 42700 40450 42756 40462
rect 42812 40796 43092 40852
rect 44044 40796 44324 40852
rect 42812 40626 42868 40796
rect 42812 40574 42814 40626
rect 42866 40574 42868 40626
rect 42700 40292 42756 40302
rect 42588 40290 42756 40292
rect 42588 40238 42702 40290
rect 42754 40238 42756 40290
rect 42588 40236 42756 40238
rect 42700 40226 42756 40236
rect 42700 39508 42756 39518
rect 42700 39414 42756 39452
rect 42812 39284 42868 40574
rect 43036 40628 43092 40638
rect 43036 40534 43092 40572
rect 42924 40292 42980 40302
rect 42924 39618 42980 40236
rect 43932 39732 43988 39742
rect 43932 39638 43988 39676
rect 42924 39566 42926 39618
rect 42978 39566 42980 39618
rect 42924 39554 42980 39566
rect 42812 39218 42868 39228
rect 43596 39394 43652 39406
rect 43596 39342 43598 39394
rect 43650 39342 43652 39394
rect 43036 39172 43092 39182
rect 42924 38722 42980 38734
rect 42924 38670 42926 38722
rect 42978 38670 42980 38722
rect 42364 38612 42644 38668
rect 42476 37042 42532 37054
rect 42476 36990 42478 37042
rect 42530 36990 42532 37042
rect 42364 36596 42420 36606
rect 42364 35700 42420 36540
rect 42364 35606 42420 35644
rect 42028 35298 42084 35308
rect 42140 35532 42308 35588
rect 42476 35588 42532 36990
rect 41692 34302 41694 34354
rect 41746 34302 41748 34354
rect 41356 33294 41358 33346
rect 41410 33294 41412 33346
rect 41356 33282 41412 33294
rect 41692 32562 41748 34302
rect 41692 32510 41694 32562
rect 41746 32510 41748 32562
rect 41692 32452 41748 32510
rect 41692 32386 41748 32396
rect 41804 35084 41916 35140
rect 41692 32116 41748 32126
rect 41244 30706 41300 30716
rect 41468 31556 41524 31566
rect 41468 31218 41524 31500
rect 41468 31166 41470 31218
rect 41522 31166 41524 31218
rect 39340 30322 39620 30324
rect 39340 30270 39342 30322
rect 39394 30270 39620 30322
rect 39340 30268 39620 30270
rect 40012 30324 40068 30334
rect 38444 29598 38446 29650
rect 38498 29598 38500 29650
rect 38444 29586 38500 29598
rect 38556 30210 38612 30222
rect 38556 30158 38558 30210
rect 38610 30158 38612 30210
rect 38556 30100 38612 30158
rect 38108 29486 38110 29538
rect 38162 29486 38164 29538
rect 38108 29474 38164 29486
rect 37772 28702 37774 28754
rect 37826 28702 37828 28754
rect 37772 28690 37828 28702
rect 38220 28644 38276 28654
rect 38108 28642 38276 28644
rect 38108 28590 38222 28642
rect 38274 28590 38276 28642
rect 38108 28588 38276 28590
rect 37772 28084 37828 28094
rect 37772 27990 37828 28028
rect 37548 27860 37604 27870
rect 37548 27766 37604 27804
rect 37996 27858 38052 27870
rect 37996 27806 37998 27858
rect 38050 27806 38052 27858
rect 37884 27748 37940 27758
rect 37996 27748 38052 27806
rect 37660 27746 38052 27748
rect 37660 27694 37886 27746
rect 37938 27694 38052 27746
rect 37660 27692 38052 27694
rect 37660 27524 37716 27692
rect 37884 27682 37940 27692
rect 37548 27468 37716 27524
rect 37548 26962 37604 27468
rect 37772 27300 37828 27310
rect 37772 27186 37828 27244
rect 37772 27134 37774 27186
rect 37826 27134 37828 27186
rect 37772 27122 37828 27134
rect 37548 26910 37550 26962
rect 37602 26910 37604 26962
rect 37548 26898 37604 26910
rect 37660 27076 37716 27086
rect 37324 26236 37492 26292
rect 37324 25394 37380 26236
rect 37660 26180 37716 27020
rect 38108 26908 38164 28588
rect 38220 28578 38276 28588
rect 38556 28644 38612 30044
rect 38892 29988 38948 29998
rect 38892 29894 38948 29932
rect 39228 29988 39284 29998
rect 39004 29538 39060 29550
rect 39004 29486 39006 29538
rect 39058 29486 39060 29538
rect 38780 29204 38836 29214
rect 38780 29110 38836 29148
rect 39004 28868 39060 29486
rect 39004 28802 39060 28812
rect 38556 28578 38612 28588
rect 39228 28642 39284 29932
rect 39340 29652 39396 30268
rect 39788 29988 39844 29998
rect 39788 29894 39844 29932
rect 39340 29586 39396 29596
rect 39228 28590 39230 28642
rect 39282 28590 39284 28642
rect 38332 28530 38388 28542
rect 38332 28478 38334 28530
rect 38386 28478 38388 28530
rect 38332 27860 38388 28478
rect 39116 28420 39172 28430
rect 39116 28326 39172 28364
rect 38444 28308 38500 28318
rect 38444 28082 38500 28252
rect 38444 28030 38446 28082
rect 38498 28030 38500 28082
rect 38444 28018 38500 28030
rect 38556 28196 38612 28206
rect 38556 28082 38612 28140
rect 38556 28030 38558 28082
rect 38610 28030 38612 28082
rect 38556 28018 38612 28030
rect 38668 28084 38724 28094
rect 39228 28084 39284 28590
rect 39676 29426 39732 29438
rect 39676 29374 39678 29426
rect 39730 29374 39732 29426
rect 39676 28644 39732 29374
rect 39900 28868 39956 28878
rect 39676 28578 39732 28588
rect 39788 28642 39844 28654
rect 39788 28590 39790 28642
rect 39842 28590 39844 28642
rect 38668 28082 39060 28084
rect 38668 28030 38670 28082
rect 38722 28030 39060 28082
rect 38668 28028 39060 28030
rect 38668 28018 38724 28028
rect 38332 27300 38388 27804
rect 38668 27860 38724 27870
rect 38332 27234 38388 27244
rect 38444 27748 38500 27758
rect 38444 26908 38500 27692
rect 38668 27074 38724 27804
rect 39004 27188 39060 28028
rect 39228 28018 39284 28028
rect 39788 28420 39844 28590
rect 39788 27748 39844 28364
rect 39788 27682 39844 27692
rect 39900 28642 39956 28812
rect 40012 28756 40068 30268
rect 41356 30212 41412 30222
rect 40124 29986 40180 29998
rect 40124 29934 40126 29986
rect 40178 29934 40180 29986
rect 40124 29652 40180 29934
rect 40460 29988 40516 29998
rect 40460 29894 40516 29932
rect 40796 29986 40852 29998
rect 40796 29934 40798 29986
rect 40850 29934 40852 29986
rect 40124 29586 40180 29596
rect 40124 29426 40180 29438
rect 40124 29374 40126 29426
rect 40178 29374 40180 29426
rect 40124 29092 40180 29374
rect 40348 29428 40404 29438
rect 40348 29334 40404 29372
rect 40236 29316 40292 29326
rect 40236 29222 40292 29260
rect 40124 29026 40180 29036
rect 40684 28868 40740 28878
rect 40236 28866 40740 28868
rect 40236 28814 40686 28866
rect 40738 28814 40740 28866
rect 40236 28812 40740 28814
rect 40124 28756 40180 28766
rect 40012 28754 40180 28756
rect 40012 28702 40126 28754
rect 40178 28702 40180 28754
rect 40012 28700 40180 28702
rect 40124 28690 40180 28700
rect 39900 28590 39902 28642
rect 39954 28590 39956 28642
rect 39900 28308 39956 28590
rect 39116 27636 39172 27646
rect 39116 27634 39284 27636
rect 39116 27582 39118 27634
rect 39170 27582 39284 27634
rect 39116 27580 39284 27582
rect 39116 27570 39172 27580
rect 39116 27188 39172 27198
rect 39004 27132 39116 27188
rect 38668 27022 38670 27074
rect 38722 27022 38724 27074
rect 38668 27010 38724 27022
rect 39116 27074 39172 27132
rect 39116 27022 39118 27074
rect 39170 27022 39172 27074
rect 38108 26852 38276 26908
rect 38444 26852 38612 26908
rect 38108 26290 38164 26302
rect 38108 26238 38110 26290
rect 38162 26238 38164 26290
rect 37660 26124 37940 26180
rect 37324 25342 37326 25394
rect 37378 25342 37380 25394
rect 37324 24164 37380 25342
rect 37436 26068 37492 26078
rect 37436 26066 37716 26068
rect 37436 26014 37438 26066
rect 37490 26014 37716 26066
rect 37436 26012 37716 26014
rect 37436 24724 37492 26012
rect 37660 25506 37716 26012
rect 37660 25454 37662 25506
rect 37714 25454 37716 25506
rect 37660 25442 37716 25454
rect 37772 25956 37828 25966
rect 37548 24948 37604 24958
rect 37772 24948 37828 25900
rect 37548 24946 37828 24948
rect 37548 24894 37550 24946
rect 37602 24894 37828 24946
rect 37548 24892 37828 24894
rect 37548 24882 37604 24892
rect 37436 24668 37604 24724
rect 37324 24098 37380 24108
rect 37324 23940 37380 23950
rect 37324 23826 37380 23884
rect 37324 23774 37326 23826
rect 37378 23774 37380 23826
rect 37324 23762 37380 23774
rect 37100 23548 37380 23604
rect 36988 23492 37044 23502
rect 36876 23436 36988 23492
rect 36652 23314 36708 23324
rect 36764 23380 36820 23390
rect 36876 23380 36932 23436
rect 36988 23426 37044 23436
rect 36764 23378 36932 23380
rect 36764 23326 36766 23378
rect 36818 23326 36932 23378
rect 36764 23324 36932 23326
rect 36764 23314 36820 23324
rect 36988 23268 37044 23278
rect 36988 23174 37044 23212
rect 36652 23156 36708 23166
rect 36652 23062 36708 23100
rect 36540 22540 36932 22596
rect 36428 22316 36596 22372
rect 36316 22278 36372 22316
rect 36428 22148 36484 22158
rect 36428 22054 36484 22092
rect 36204 21084 36484 21140
rect 36316 20914 36372 20926
rect 36316 20862 36318 20914
rect 36370 20862 36372 20914
rect 35980 20066 36036 20076
rect 36204 20802 36260 20814
rect 36204 20750 36206 20802
rect 36258 20750 36260 20802
rect 36092 20020 36148 20030
rect 36092 19926 36148 19964
rect 35812 19180 35924 19236
rect 35980 19908 36036 19918
rect 35756 19142 35812 19180
rect 35756 18564 35812 18574
rect 35644 18562 35924 18564
rect 35644 18510 35758 18562
rect 35810 18510 35924 18562
rect 35644 18508 35924 18510
rect 35756 18498 35812 18508
rect 35868 18228 35924 18508
rect 35756 17780 35812 17790
rect 35532 17778 35812 17780
rect 35532 17726 35758 17778
rect 35810 17726 35812 17778
rect 35532 17724 35812 17726
rect 35756 17714 35812 17724
rect 35868 17780 35924 18172
rect 35868 17714 35924 17724
rect 34748 17666 35028 17668
rect 34748 17614 34974 17666
rect 35026 17614 35028 17666
rect 34748 17612 35028 17614
rect 34748 16994 34804 17612
rect 34972 17602 35028 17612
rect 34748 16942 34750 16994
rect 34802 16942 34804 16994
rect 34748 16930 34804 16942
rect 35084 17442 35140 17454
rect 35084 17390 35086 17442
rect 35138 17390 35140 17442
rect 34524 16830 34526 16882
rect 34578 16830 34580 16882
rect 34524 16818 34580 16830
rect 34972 16884 35028 16894
rect 35084 16884 35140 17390
rect 35308 17444 35364 17454
rect 35308 17442 35588 17444
rect 35308 17390 35310 17442
rect 35362 17390 35588 17442
rect 35308 17388 35588 17390
rect 35308 17378 35364 17388
rect 34972 16882 35140 16884
rect 34972 16830 34974 16882
rect 35026 16830 35140 16882
rect 34972 16828 35140 16830
rect 35308 16882 35364 16894
rect 35308 16830 35310 16882
rect 35362 16830 35364 16882
rect 33964 16770 34020 16782
rect 33964 16718 33966 16770
rect 34018 16718 34020 16770
rect 33964 15148 34020 16718
rect 34860 16770 34916 16782
rect 34860 16718 34862 16770
rect 34914 16718 34916 16770
rect 34300 15986 34356 15998
rect 34300 15934 34302 15986
rect 34354 15934 34356 15986
rect 34300 15540 34356 15934
rect 34636 15876 34692 15886
rect 34412 15540 34468 15550
rect 34300 15538 34468 15540
rect 34300 15486 34414 15538
rect 34466 15486 34468 15538
rect 34300 15484 34468 15486
rect 34412 15474 34468 15484
rect 34076 15316 34132 15326
rect 34524 15316 34580 15326
rect 34076 15314 34580 15316
rect 34076 15262 34078 15314
rect 34130 15262 34526 15314
rect 34578 15262 34580 15314
rect 34076 15260 34580 15262
rect 34076 15250 34132 15260
rect 34524 15250 34580 15260
rect 34636 15148 34692 15820
rect 34860 15314 34916 16718
rect 34860 15262 34862 15314
rect 34914 15262 34916 15314
rect 34860 15250 34916 15262
rect 33964 15092 34132 15148
rect 33964 14756 34020 14766
rect 33964 13858 34020 14700
rect 33964 13806 33966 13858
rect 34018 13806 34020 13858
rect 33964 13794 34020 13806
rect 34076 13300 34132 15092
rect 34300 15090 34356 15102
rect 34300 15038 34302 15090
rect 34354 15038 34356 15090
rect 34188 14308 34244 14318
rect 34300 14308 34356 15038
rect 34412 15092 34692 15148
rect 34412 14530 34468 15092
rect 34636 14980 34692 14990
rect 34524 14756 34580 14766
rect 34524 14662 34580 14700
rect 34412 14478 34414 14530
rect 34466 14478 34468 14530
rect 34412 14466 34468 14478
rect 34524 14420 34580 14430
rect 34188 14306 34356 14308
rect 34188 14254 34190 14306
rect 34242 14254 34356 14306
rect 34188 14252 34356 14254
rect 34412 14308 34468 14318
rect 34188 14242 34244 14252
rect 34076 13244 34356 13300
rect 34076 12852 34132 12862
rect 34076 12758 34132 12796
rect 33740 12460 34132 12516
rect 32844 12348 33124 12404
rect 32956 12180 33012 12190
rect 32284 12178 33012 12180
rect 32284 12126 32958 12178
rect 33010 12126 33012 12178
rect 32284 12124 33012 12126
rect 32284 11394 32340 12124
rect 32956 12114 33012 12124
rect 33068 11732 33124 12348
rect 33180 12290 33236 12302
rect 33180 12238 33182 12290
rect 33234 12238 33236 12290
rect 33180 12068 33236 12238
rect 33292 12290 33348 12460
rect 33964 12292 34020 12302
rect 33292 12238 33294 12290
rect 33346 12238 33348 12290
rect 33292 12226 33348 12238
rect 33404 12290 34020 12292
rect 33404 12238 33966 12290
rect 34018 12238 34020 12290
rect 33404 12236 34020 12238
rect 33180 12002 33236 12012
rect 32284 11342 32286 11394
rect 32338 11342 32340 11394
rect 32284 11330 32340 11342
rect 32844 11676 33124 11732
rect 33292 11956 33348 11966
rect 32732 11172 32788 11182
rect 32172 11170 32788 11172
rect 32172 11118 32734 11170
rect 32786 11118 32788 11170
rect 32172 11116 32788 11118
rect 32732 11106 32788 11116
rect 31500 10780 31892 10836
rect 31388 10668 31556 10724
rect 31500 10610 31556 10668
rect 31500 10558 31502 10610
rect 31554 10558 31556 10610
rect 31500 10546 31556 10558
rect 31388 10498 31444 10510
rect 31388 10446 31390 10498
rect 31442 10446 31444 10498
rect 31276 10388 31332 10398
rect 31276 10294 31332 10332
rect 31388 10164 31444 10446
rect 31276 10108 31444 10164
rect 31276 10052 31332 10108
rect 31276 9986 31332 9996
rect 31724 10050 31780 10062
rect 31724 9998 31726 10050
rect 31778 9998 31780 10050
rect 31388 9940 31444 9950
rect 31388 9846 31444 9884
rect 31164 9660 31556 9716
rect 30940 9214 30942 9266
rect 30994 9214 30996 9266
rect 30940 9202 30996 9214
rect 31276 9380 31332 9390
rect 31276 9266 31332 9324
rect 31276 9214 31278 9266
rect 31330 9214 31332 9266
rect 31276 9202 31332 9214
rect 31500 9266 31556 9660
rect 31500 9214 31502 9266
rect 31554 9214 31556 9266
rect 31500 9202 31556 9214
rect 31612 9268 31668 9278
rect 31612 9174 31668 9212
rect 31724 9266 31780 9998
rect 31724 9214 31726 9266
rect 31778 9214 31780 9266
rect 31724 9202 31780 9214
rect 30716 8204 30884 8260
rect 31164 8820 31220 8830
rect 30044 7420 30212 7476
rect 30492 7476 30548 7486
rect 30044 7364 30100 7420
rect 29820 6690 29876 6748
rect 29820 6638 29822 6690
rect 29874 6638 29876 6690
rect 29820 6626 29876 6638
rect 29932 7308 30100 7364
rect 30268 7364 30324 7374
rect 29484 6300 29764 6356
rect 29596 5684 29652 5694
rect 29596 5010 29652 5628
rect 29596 4958 29598 5010
rect 29650 4958 29652 5010
rect 29596 4946 29652 4958
rect 28924 3666 29428 3668
rect 28924 3614 28926 3666
rect 28978 3614 29428 3666
rect 28924 3612 29428 3614
rect 29596 4340 29652 4350
rect 29596 3666 29652 4284
rect 29596 3614 29598 3666
rect 29650 3614 29652 3666
rect 27916 3602 27972 3612
rect 28924 3602 28980 3612
rect 29596 3602 29652 3614
rect 27020 3390 27022 3442
rect 27074 3390 27076 3442
rect 27020 3378 27076 3390
rect 29484 3556 29540 3566
rect 29484 3388 29540 3500
rect 29708 3444 29764 6300
rect 29932 6130 29988 7308
rect 30268 7252 30324 7308
rect 30044 7250 30324 7252
rect 30044 7198 30270 7250
rect 30322 7198 30324 7250
rect 30044 7196 30324 7198
rect 30044 6914 30100 7196
rect 30268 7186 30324 7196
rect 30044 6862 30046 6914
rect 30098 6862 30100 6914
rect 30044 6850 30100 6862
rect 30268 6916 30324 6926
rect 30268 6804 30324 6860
rect 30492 6916 30548 7420
rect 30492 6850 30548 6860
rect 30156 6748 30324 6804
rect 30044 6690 30100 6702
rect 30044 6638 30046 6690
rect 30098 6638 30100 6690
rect 30044 6356 30100 6638
rect 30044 6290 30100 6300
rect 29932 6078 29934 6130
rect 29986 6078 29988 6130
rect 29932 6066 29988 6078
rect 30156 6020 30212 6748
rect 30716 6132 30772 8204
rect 30828 8036 30884 8046
rect 30828 7586 30884 7980
rect 31164 7698 31220 8764
rect 31164 7646 31166 7698
rect 31218 7646 31220 7698
rect 31164 7634 31220 7646
rect 31388 8260 31444 8270
rect 30828 7534 30830 7586
rect 30882 7534 30884 7586
rect 30828 7522 30884 7534
rect 31052 7474 31108 7486
rect 31052 7422 31054 7474
rect 31106 7422 31108 7474
rect 30940 6804 30996 6814
rect 31052 6804 31108 7422
rect 30996 6748 31108 6804
rect 30940 6578 30996 6748
rect 30940 6526 30942 6578
rect 30994 6526 30996 6578
rect 30940 6514 30996 6526
rect 31276 6468 31332 6478
rect 31276 6374 31332 6412
rect 31388 6244 31444 8204
rect 31500 8036 31556 8046
rect 31500 7474 31556 7980
rect 31500 7422 31502 7474
rect 31554 7422 31556 7474
rect 31500 7410 31556 7422
rect 31612 6916 31668 6926
rect 31612 6822 31668 6860
rect 31724 6578 31780 6590
rect 31724 6526 31726 6578
rect 31778 6526 31780 6578
rect 31724 6356 31780 6526
rect 31724 6290 31780 6300
rect 31388 6178 31444 6188
rect 30716 6076 30884 6132
rect 30156 5906 30212 5964
rect 30156 5854 30158 5906
rect 30210 5854 30212 5906
rect 30156 5842 30212 5854
rect 30380 5682 30436 5694
rect 30380 5630 30382 5682
rect 30434 5630 30436 5682
rect 30380 5572 30436 5630
rect 30380 5506 30436 5516
rect 30716 5682 30772 5694
rect 30716 5630 30718 5682
rect 30770 5630 30772 5682
rect 30156 5124 30212 5134
rect 30156 4450 30212 5068
rect 30716 5124 30772 5630
rect 30716 5058 30772 5068
rect 30828 5012 30884 6076
rect 31612 6130 31668 6142
rect 31612 6078 31614 6130
rect 31666 6078 31668 6130
rect 31052 6020 31108 6030
rect 31612 6020 31668 6078
rect 31108 5964 31220 6020
rect 31052 5926 31108 5964
rect 31164 5684 31220 5964
rect 31612 5954 31668 5964
rect 31276 5906 31332 5918
rect 31276 5854 31278 5906
rect 31330 5854 31332 5906
rect 31276 5796 31332 5854
rect 31724 5908 31780 5918
rect 31276 5740 31556 5796
rect 31164 5628 31444 5684
rect 31388 5346 31444 5628
rect 31388 5294 31390 5346
rect 31442 5294 31444 5346
rect 31388 5282 31444 5294
rect 31500 5572 31556 5740
rect 31556 5516 31668 5572
rect 30828 4946 30884 4956
rect 31388 4564 31444 4574
rect 31500 4564 31556 5516
rect 31612 5234 31668 5516
rect 31724 5346 31780 5852
rect 31724 5294 31726 5346
rect 31778 5294 31780 5346
rect 31724 5282 31780 5294
rect 31612 5182 31614 5234
rect 31666 5182 31668 5234
rect 31612 5170 31668 5182
rect 31388 4562 31556 4564
rect 31388 4510 31390 4562
rect 31442 4510 31556 4562
rect 31388 4508 31556 4510
rect 31388 4498 31444 4508
rect 30156 4398 30158 4450
rect 30210 4398 30212 4450
rect 30044 3556 30100 3566
rect 30156 3556 30212 4398
rect 31052 3892 31108 3902
rect 31052 3666 31108 3836
rect 31052 3614 31054 3666
rect 31106 3614 31108 3666
rect 31052 3602 31108 3614
rect 31500 3668 31556 3678
rect 30268 3556 30324 3566
rect 30156 3500 30268 3556
rect 30044 3462 30100 3500
rect 30268 3490 30324 3500
rect 31388 3556 31444 3566
rect 31500 3556 31556 3612
rect 31388 3554 31556 3556
rect 31388 3502 31390 3554
rect 31442 3502 31556 3554
rect 31388 3500 31556 3502
rect 31388 3490 31444 3500
rect 29820 3444 29876 3454
rect 29708 3442 29876 3444
rect 29708 3390 29822 3442
rect 29874 3390 29876 3442
rect 29708 3388 29876 3390
rect 29484 3332 29652 3388
rect 29820 3378 29876 3388
rect 23100 3220 23156 3332
rect 23212 3220 23268 3230
rect 19836 3164 20100 3174
rect 23100 3164 23212 3220
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 23212 3154 23268 3164
rect 19836 3098 20100 3108
rect 13804 2930 13860 2940
rect 29596 800 29652 3332
rect 31500 1764 31556 3500
rect 31612 3444 31668 3454
rect 31836 3444 31892 10780
rect 31948 9828 32004 9838
rect 31948 8820 32004 9772
rect 32508 9604 32564 9614
rect 32508 9510 32564 9548
rect 32396 9156 32452 9166
rect 32284 9044 32340 9054
rect 32284 8950 32340 8988
rect 31948 8754 32004 8764
rect 32172 8484 32228 8494
rect 32060 8372 32116 8382
rect 31948 8370 32116 8372
rect 31948 8318 32062 8370
rect 32114 8318 32116 8370
rect 31948 8316 32116 8318
rect 31948 6804 32004 8316
rect 32060 8306 32116 8316
rect 32060 7364 32116 7374
rect 32172 7364 32228 8428
rect 32396 7924 32452 9100
rect 32508 9044 32564 9054
rect 32508 8484 32564 8988
rect 32508 8418 32564 8428
rect 32620 9042 32676 9054
rect 32620 8990 32622 9042
rect 32674 8990 32676 9042
rect 32620 8146 32676 8990
rect 32620 8094 32622 8146
rect 32674 8094 32676 8146
rect 32620 8082 32676 8094
rect 32732 8372 32788 8382
rect 32396 7868 32676 7924
rect 32060 7362 32228 7364
rect 32060 7310 32062 7362
rect 32114 7310 32228 7362
rect 32060 7308 32228 7310
rect 32508 7474 32564 7486
rect 32508 7422 32510 7474
rect 32562 7422 32564 7474
rect 32060 7298 32116 7308
rect 31948 6738 32004 6748
rect 32172 7028 32228 7038
rect 32172 6802 32228 6972
rect 32508 6916 32564 7422
rect 32620 7028 32676 7868
rect 32620 6962 32676 6972
rect 32508 6850 32564 6860
rect 32172 6750 32174 6802
rect 32226 6750 32228 6802
rect 32172 6738 32228 6750
rect 32060 6692 32116 6702
rect 31948 6468 32004 6478
rect 31948 5460 32004 6412
rect 32060 5794 32116 6636
rect 32620 6692 32676 6702
rect 32732 6692 32788 8316
rect 32620 6690 32788 6692
rect 32620 6638 32622 6690
rect 32674 6638 32788 6690
rect 32620 6636 32788 6638
rect 32620 6626 32676 6636
rect 32620 6244 32676 6254
rect 32508 6188 32620 6244
rect 32676 6188 32788 6244
rect 32060 5742 32062 5794
rect 32114 5742 32116 5794
rect 32060 5730 32116 5742
rect 32396 5908 32452 5918
rect 32060 5460 32116 5470
rect 31948 5404 32060 5460
rect 31948 4338 32004 5404
rect 32060 5394 32116 5404
rect 32060 5124 32116 5134
rect 32060 5030 32116 5068
rect 32172 5012 32228 5022
rect 32172 4918 32228 4956
rect 31948 4286 31950 4338
rect 32002 4286 32004 4338
rect 31948 4274 32004 4286
rect 32396 4338 32452 5852
rect 32508 5906 32564 6188
rect 32620 6178 32676 6188
rect 32508 5854 32510 5906
rect 32562 5854 32564 5906
rect 32508 5842 32564 5854
rect 32620 6020 32676 6030
rect 32396 4286 32398 4338
rect 32450 4286 32452 4338
rect 32396 4274 32452 4286
rect 32508 5684 32564 5694
rect 31612 3442 31892 3444
rect 31612 3390 31614 3442
rect 31666 3390 31892 3442
rect 31612 3388 31892 3390
rect 32284 3444 32340 3454
rect 32396 3444 32452 3454
rect 32340 3442 32452 3444
rect 32340 3390 32398 3442
rect 32450 3390 32452 3442
rect 32340 3388 32452 3390
rect 32508 3444 32564 5628
rect 32620 4004 32676 5964
rect 32732 4564 32788 6188
rect 32844 5684 32900 11676
rect 33292 11394 33348 11900
rect 33404 11506 33460 12236
rect 33964 12226 34020 12236
rect 33404 11454 33406 11506
rect 33458 11454 33460 11506
rect 33404 11442 33460 11454
rect 33516 12068 33572 12078
rect 33292 11342 33294 11394
rect 33346 11342 33348 11394
rect 33292 11330 33348 11342
rect 33516 11394 33572 12012
rect 33516 11342 33518 11394
rect 33570 11342 33572 11394
rect 33516 11330 33572 11342
rect 34076 11396 34132 12460
rect 34300 11618 34356 13244
rect 34412 12962 34468 14252
rect 34524 13746 34580 14364
rect 34524 13694 34526 13746
rect 34578 13694 34580 13746
rect 34524 13682 34580 13694
rect 34412 12910 34414 12962
rect 34466 12910 34468 12962
rect 34412 12898 34468 12910
rect 34524 13074 34580 13086
rect 34524 13022 34526 13074
rect 34578 13022 34580 13074
rect 34524 12964 34580 13022
rect 34524 12740 34580 12908
rect 34524 12674 34580 12684
rect 34300 11566 34302 11618
rect 34354 11566 34356 11618
rect 34300 11554 34356 11566
rect 34076 11340 34356 11396
rect 33068 11172 33124 11182
rect 33068 11078 33124 11116
rect 33964 11172 34020 11182
rect 33964 11078 34020 11116
rect 33516 10836 33572 10846
rect 33516 10742 33572 10780
rect 33180 10722 33236 10734
rect 33180 10670 33182 10722
rect 33234 10670 33236 10722
rect 33180 10612 33236 10670
rect 33404 10724 33460 10734
rect 33404 10612 33460 10668
rect 34188 10724 34244 10734
rect 33180 10546 33236 10556
rect 33292 10610 33460 10612
rect 33292 10558 33406 10610
rect 33458 10558 33460 10610
rect 33292 10556 33460 10558
rect 33292 9828 33348 10556
rect 33404 10546 33460 10556
rect 33628 10612 33684 10622
rect 33964 10612 34020 10622
rect 33628 10610 34020 10612
rect 33628 10558 33630 10610
rect 33682 10558 33966 10610
rect 34018 10558 34020 10610
rect 33628 10556 34020 10558
rect 33628 10546 33684 10556
rect 33292 9762 33348 9772
rect 32956 9714 33012 9726
rect 32956 9662 32958 9714
rect 33010 9662 33012 9714
rect 32956 9156 33012 9662
rect 32956 9090 33012 9100
rect 33404 9714 33460 9726
rect 33404 9662 33406 9714
rect 33458 9662 33460 9714
rect 33404 9604 33460 9662
rect 33404 9042 33460 9548
rect 33404 8990 33406 9042
rect 33458 8990 33460 9042
rect 33404 8428 33460 8990
rect 33628 8932 33684 8942
rect 33628 8838 33684 8876
rect 33740 8596 33796 10556
rect 33964 10546 34020 10556
rect 34076 10612 34132 10622
rect 34076 9938 34132 10556
rect 34188 10610 34244 10668
rect 34188 10558 34190 10610
rect 34242 10558 34244 10610
rect 34188 10546 34244 10558
rect 34300 10388 34356 11340
rect 34636 10722 34692 14924
rect 34972 14980 35028 16828
rect 35308 16660 35364 16830
rect 35532 16882 35588 17388
rect 35644 17442 35700 17454
rect 35644 17390 35646 17442
rect 35698 17390 35700 17442
rect 35644 17220 35700 17390
rect 35868 17444 35924 17454
rect 35868 17350 35924 17388
rect 35980 17220 36036 19852
rect 36204 19572 36260 20750
rect 36316 20580 36372 20862
rect 36316 20514 36372 20524
rect 36204 19516 36372 19572
rect 36204 19346 36260 19358
rect 36204 19294 36206 19346
rect 36258 19294 36260 19346
rect 36092 19234 36148 19246
rect 36092 19182 36094 19234
rect 36146 19182 36148 19234
rect 36092 19012 36148 19182
rect 36092 18946 36148 18956
rect 36204 18788 36260 19294
rect 36204 18722 36260 18732
rect 36204 18450 36260 18462
rect 36204 18398 36206 18450
rect 36258 18398 36260 18450
rect 36092 18340 36148 18350
rect 36092 17780 36148 18284
rect 36092 17554 36148 17724
rect 36092 17502 36094 17554
rect 36146 17502 36148 17554
rect 36092 17490 36148 17502
rect 35644 17164 36036 17220
rect 35532 16830 35534 16882
rect 35586 16830 35588 16882
rect 35532 16818 35588 16830
rect 35644 16940 35924 16996
rect 35644 16660 35700 16940
rect 35868 16882 35924 16940
rect 35868 16830 35870 16882
rect 35922 16830 35924 16882
rect 35308 16604 35700 16660
rect 35756 16770 35812 16782
rect 35756 16718 35758 16770
rect 35810 16718 35812 16770
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34972 14914 35028 14924
rect 35084 15764 35140 15774
rect 34748 14420 34804 14430
rect 34748 14326 34804 14364
rect 34972 14420 35028 14430
rect 34972 14326 35028 14364
rect 34636 10670 34638 10722
rect 34690 10670 34692 10722
rect 34636 10658 34692 10670
rect 34748 14196 34804 14206
rect 34076 9886 34078 9938
rect 34130 9886 34132 9938
rect 34076 9874 34132 9886
rect 34188 10332 34356 10388
rect 33964 9828 34020 9838
rect 33852 9156 33908 9166
rect 33852 9062 33908 9100
rect 33964 9044 34020 9772
rect 33964 8950 34020 8988
rect 33740 8540 33908 8596
rect 33404 8372 33796 8428
rect 33292 8258 33348 8270
rect 33292 8206 33294 8258
rect 33346 8206 33348 8258
rect 32956 8148 33012 8158
rect 32956 7700 33012 8092
rect 32956 7644 33236 7700
rect 32956 6692 33012 7644
rect 33180 7586 33236 7644
rect 33180 7534 33182 7586
rect 33234 7534 33236 7586
rect 33180 7522 33236 7534
rect 33292 7476 33348 8206
rect 33628 8036 33684 8046
rect 33628 7942 33684 7980
rect 33516 7476 33572 7486
rect 33292 7420 33516 7476
rect 33516 7382 33572 7420
rect 33180 7364 33236 7374
rect 33180 7270 33236 7308
rect 33292 6916 33348 6926
rect 33292 6822 33348 6860
rect 33628 6802 33684 6814
rect 33628 6750 33630 6802
rect 33682 6750 33684 6802
rect 32956 6626 33012 6636
rect 33516 6690 33572 6702
rect 33516 6638 33518 6690
rect 33570 6638 33572 6690
rect 33516 6244 33572 6638
rect 33628 6468 33684 6750
rect 33628 6402 33684 6412
rect 32844 5618 32900 5628
rect 33068 5906 33124 5918
rect 33068 5854 33070 5906
rect 33122 5854 33124 5906
rect 33068 5796 33124 5854
rect 33292 5908 33348 5918
rect 33292 5814 33348 5852
rect 33516 5908 33572 6188
rect 33516 5842 33572 5852
rect 33068 5122 33124 5740
rect 33628 5796 33684 5806
rect 33068 5070 33070 5122
rect 33122 5070 33124 5122
rect 33068 5058 33124 5070
rect 33404 5348 33460 5358
rect 33404 4564 33460 5292
rect 32732 4508 33012 4564
rect 32956 4452 33012 4508
rect 33180 4508 33460 4564
rect 33516 5012 33572 5022
rect 33068 4452 33124 4462
rect 32956 4450 33124 4452
rect 32956 4398 33070 4450
rect 33122 4398 33124 4450
rect 32956 4396 33124 4398
rect 33068 4386 33124 4396
rect 32620 3948 33124 4004
rect 32956 3780 33012 3790
rect 32732 3444 32788 3454
rect 32508 3442 32788 3444
rect 32508 3390 32734 3442
rect 32786 3390 32788 3442
rect 32508 3388 32788 3390
rect 31612 3378 31668 3388
rect 31500 1708 31668 1764
rect 31612 800 31668 1708
rect 32284 800 32340 3388
rect 32396 3378 32452 3388
rect 32732 3378 32788 3388
rect 32956 800 33012 3724
rect 33068 3554 33124 3948
rect 33068 3502 33070 3554
rect 33122 3502 33124 3554
rect 33068 3490 33124 3502
rect 33180 3556 33236 4508
rect 33404 4340 33460 4350
rect 33404 4246 33460 4284
rect 33516 3666 33572 4956
rect 33516 3614 33518 3666
rect 33570 3614 33572 3666
rect 33516 3602 33572 3614
rect 33404 3556 33460 3566
rect 33180 3554 33460 3556
rect 33180 3502 33406 3554
rect 33458 3502 33460 3554
rect 33180 3500 33460 3502
rect 33404 3490 33460 3500
rect 33628 3554 33684 5740
rect 33740 4564 33796 8372
rect 33852 7588 33908 8540
rect 33852 7140 33908 7532
rect 33852 7074 33908 7084
rect 33964 8258 34020 8270
rect 33964 8206 33966 8258
rect 34018 8206 34020 8258
rect 33964 6916 34020 8206
rect 33964 6850 34020 6860
rect 34076 7474 34132 7486
rect 34076 7422 34078 7474
rect 34130 7422 34132 7474
rect 34076 6244 34132 7422
rect 34188 7364 34244 10332
rect 34524 9828 34580 9838
rect 34524 9734 34580 9772
rect 34748 9380 34804 14140
rect 34860 13746 34916 13758
rect 34860 13694 34862 13746
rect 34914 13694 34916 13746
rect 34860 13524 34916 13694
rect 34860 13458 34916 13468
rect 35084 12740 35140 15708
rect 35532 15428 35588 15438
rect 35756 15428 35812 16718
rect 35532 15426 35812 15428
rect 35532 15374 35534 15426
rect 35586 15374 35812 15426
rect 35532 15372 35812 15374
rect 35532 15362 35588 15372
rect 35868 15092 35924 16830
rect 36092 16882 36148 16894
rect 36092 16830 36094 16882
rect 36146 16830 36148 16882
rect 36092 15148 36148 16830
rect 35644 15036 35868 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35532 14756 35588 14766
rect 35532 14662 35588 14700
rect 35532 14532 35588 14542
rect 35644 14532 35700 15036
rect 35868 15026 35924 15036
rect 35980 15092 36148 15148
rect 35980 14642 36036 15092
rect 35980 14590 35982 14642
rect 36034 14590 36036 14642
rect 35980 14578 36036 14590
rect 35532 14530 35700 14532
rect 35532 14478 35534 14530
rect 35586 14478 35700 14530
rect 35532 14476 35700 14478
rect 35868 14532 35924 14542
rect 35532 14466 35588 14476
rect 35868 14418 35924 14476
rect 35868 14366 35870 14418
rect 35922 14366 35924 14418
rect 35868 14196 35924 14366
rect 36092 14420 36148 14430
rect 36092 14326 36148 14364
rect 35868 14130 35924 14140
rect 35644 13972 35700 13982
rect 35644 13970 35812 13972
rect 35644 13918 35646 13970
rect 35698 13918 35812 13970
rect 35644 13916 35812 13918
rect 35644 13906 35700 13916
rect 35420 13860 35476 13870
rect 35420 13766 35476 13804
rect 35196 13748 35252 13758
rect 35196 13654 35252 13692
rect 35644 13524 35700 13534
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35532 13188 35588 13198
rect 35644 13188 35700 13468
rect 35532 13186 35700 13188
rect 35532 13134 35534 13186
rect 35586 13134 35700 13186
rect 35532 13132 35700 13134
rect 35532 13122 35588 13132
rect 35308 13074 35364 13086
rect 35308 13022 35310 13074
rect 35362 13022 35364 13074
rect 35196 12964 35252 12974
rect 35196 12870 35252 12908
rect 34972 12684 35140 12740
rect 34860 11282 34916 11294
rect 34860 11230 34862 11282
rect 34914 11230 34916 11282
rect 34860 10836 34916 11230
rect 34972 10948 35028 12684
rect 35308 12404 35364 13022
rect 35532 12962 35588 12974
rect 35532 12910 35534 12962
rect 35586 12910 35588 12962
rect 35532 12852 35588 12910
rect 35532 12786 35588 12796
rect 35308 12338 35364 12348
rect 35756 11956 35812 13916
rect 36204 13860 36260 18398
rect 36316 17444 36372 19516
rect 36316 17378 36372 17388
rect 36428 18452 36484 21084
rect 36540 19348 36596 22316
rect 36540 19282 36596 19292
rect 36876 18676 36932 22540
rect 37324 22036 37380 23548
rect 37436 23492 37492 23502
rect 37436 23378 37492 23436
rect 37436 23326 37438 23378
rect 37490 23326 37492 23378
rect 37436 23314 37492 23326
rect 37548 23266 37604 24668
rect 37548 23214 37550 23266
rect 37602 23214 37604 23266
rect 37548 23202 37604 23214
rect 37884 22708 37940 26124
rect 38108 25956 38164 26238
rect 38108 25890 38164 25900
rect 38108 25732 38164 25742
rect 38108 25396 38164 25676
rect 38220 25620 38276 26796
rect 38556 26178 38612 26852
rect 38556 26126 38558 26178
rect 38610 26126 38612 26178
rect 38556 26114 38612 26126
rect 39004 26292 39060 26302
rect 38220 25554 38276 25564
rect 38556 25508 38612 25518
rect 38332 25506 38612 25508
rect 38332 25454 38558 25506
rect 38610 25454 38612 25506
rect 38332 25452 38612 25454
rect 38220 25396 38276 25406
rect 38108 25394 38276 25396
rect 38108 25342 38222 25394
rect 38274 25342 38276 25394
rect 38108 25340 38276 25342
rect 38108 24836 38164 24846
rect 38220 24836 38276 25340
rect 38332 24946 38388 25452
rect 38556 25442 38612 25452
rect 38332 24894 38334 24946
rect 38386 24894 38388 24946
rect 38332 24882 38388 24894
rect 38892 25284 38948 25294
rect 38108 24834 38276 24836
rect 38108 24782 38110 24834
rect 38162 24782 38276 24834
rect 38108 24780 38276 24782
rect 38108 24770 38164 24780
rect 37996 24722 38052 24734
rect 37996 24670 37998 24722
rect 38050 24670 38052 24722
rect 37996 23156 38052 24670
rect 37996 23090 38052 23100
rect 38108 24164 38164 24174
rect 37996 22932 38052 22942
rect 37996 22838 38052 22876
rect 37884 22652 38052 22708
rect 37548 22372 37604 22382
rect 37548 22260 37604 22316
rect 37548 22258 37940 22260
rect 37548 22206 37550 22258
rect 37602 22206 37940 22258
rect 37548 22204 37940 22206
rect 37548 22194 37604 22204
rect 37324 21980 37604 22036
rect 37100 20802 37156 20814
rect 37100 20750 37102 20802
rect 37154 20750 37156 20802
rect 37100 19012 37156 20750
rect 37436 20692 37492 20702
rect 37212 20578 37268 20590
rect 37212 20526 37214 20578
rect 37266 20526 37268 20578
rect 37212 20020 37268 20526
rect 37212 19954 37268 19964
rect 37324 20018 37380 20030
rect 37324 19966 37326 20018
rect 37378 19966 37380 20018
rect 37324 19908 37380 19966
rect 37324 19842 37380 19852
rect 37100 18918 37156 18956
rect 36428 16436 36484 18396
rect 36764 18674 36932 18676
rect 36764 18622 36878 18674
rect 36930 18622 36932 18674
rect 36764 18620 36932 18622
rect 36316 16380 36484 16436
rect 36652 18004 36708 18014
rect 36316 13972 36372 16380
rect 36428 16210 36484 16222
rect 36428 16158 36430 16210
rect 36482 16158 36484 16210
rect 36428 16100 36484 16158
rect 36428 16034 36484 16044
rect 36540 14420 36596 14430
rect 36316 13916 36484 13972
rect 36092 13804 36260 13860
rect 35980 13748 36036 13758
rect 35980 13654 36036 13692
rect 35868 12404 35924 12414
rect 35868 12310 35924 12348
rect 35756 11890 35812 11900
rect 36092 12178 36148 13804
rect 36428 13748 36484 13916
rect 36092 12126 36094 12178
rect 36146 12126 36148 12178
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34972 10882 35028 10892
rect 35084 11508 35140 11518
rect 35084 11394 35140 11452
rect 35868 11508 35924 11518
rect 35924 11452 36036 11508
rect 35868 11414 35924 11452
rect 35084 11342 35086 11394
rect 35138 11342 35140 11394
rect 34860 10770 34916 10780
rect 34972 10612 35028 10622
rect 35084 10612 35140 11342
rect 35196 10612 35252 10622
rect 35084 10610 35252 10612
rect 35084 10558 35198 10610
rect 35250 10558 35252 10610
rect 35084 10556 35252 10558
rect 34972 10518 35028 10556
rect 35196 10546 35252 10556
rect 35980 10610 36036 11452
rect 35980 10558 35982 10610
rect 36034 10558 36036 10610
rect 35980 10546 36036 10558
rect 36092 10834 36148 12126
rect 36092 10782 36094 10834
rect 36146 10782 36148 10834
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35420 9826 35476 9838
rect 35420 9774 35422 9826
rect 35474 9774 35476 9826
rect 34524 9324 34804 9380
rect 34972 9714 35028 9726
rect 34972 9662 34974 9714
rect 35026 9662 35028 9714
rect 34412 8372 34468 8382
rect 34412 8258 34468 8316
rect 34412 8206 34414 8258
rect 34466 8206 34468 8258
rect 34412 8194 34468 8206
rect 34300 8034 34356 8046
rect 34300 7982 34302 8034
rect 34354 7982 34356 8034
rect 34300 7476 34356 7982
rect 34524 7924 34580 9324
rect 34748 9154 34804 9166
rect 34748 9102 34750 9154
rect 34802 9102 34804 9154
rect 34748 9044 34804 9102
rect 34972 9156 35028 9662
rect 34972 9090 35028 9100
rect 34748 8978 34804 8988
rect 34860 9042 34916 9054
rect 34860 8990 34862 9042
rect 34914 8990 34916 9042
rect 34860 8932 34916 8990
rect 34748 8818 34804 8830
rect 34748 8766 34750 8818
rect 34802 8766 34804 8818
rect 34636 8148 34692 8158
rect 34636 8054 34692 8092
rect 34524 7868 34692 7924
rect 34524 7476 34580 7486
rect 34300 7474 34580 7476
rect 34300 7422 34526 7474
rect 34578 7422 34580 7474
rect 34300 7420 34580 7422
rect 34524 7410 34580 7420
rect 34188 7308 34468 7364
rect 34300 6690 34356 6702
rect 34300 6638 34302 6690
rect 34354 6638 34356 6690
rect 34300 6356 34356 6638
rect 34300 6290 34356 6300
rect 33964 6188 34132 6244
rect 33964 5348 34020 6188
rect 34076 6020 34132 6030
rect 34076 5926 34132 5964
rect 33964 5122 34020 5292
rect 33964 5070 33966 5122
rect 34018 5070 34020 5122
rect 33964 5058 34020 5070
rect 34300 5908 34356 5918
rect 34300 5124 34356 5852
rect 34300 5058 34356 5068
rect 33964 4564 34020 4574
rect 33740 4562 34020 4564
rect 33740 4510 33966 4562
rect 34018 4510 34020 4562
rect 33740 4508 34020 4510
rect 33964 4498 34020 4508
rect 33628 3502 33630 3554
rect 33682 3502 33684 3554
rect 33628 3490 33684 3502
rect 33964 3780 34020 3790
rect 33964 3554 34020 3724
rect 33964 3502 33966 3554
rect 34018 3502 34020 3554
rect 33964 3490 34020 3502
rect 34300 3444 34356 3454
rect 34412 3444 34468 7308
rect 34524 6580 34580 6590
rect 34524 5794 34580 6524
rect 34524 5742 34526 5794
rect 34578 5742 34580 5794
rect 34524 5730 34580 5742
rect 34300 3442 34468 3444
rect 34300 3390 34302 3442
rect 34354 3390 34468 3442
rect 34300 3388 34468 3390
rect 34636 3442 34692 7868
rect 34748 7364 34804 8766
rect 34748 7298 34804 7308
rect 34860 6020 34916 8876
rect 35420 8820 35476 9774
rect 36092 9828 36148 10782
rect 36092 9762 36148 9772
rect 36204 13692 36484 13748
rect 35980 9716 36036 9726
rect 35980 9622 36036 9660
rect 35532 9604 35588 9614
rect 35532 9510 35588 9548
rect 36092 9602 36148 9614
rect 36092 9550 36094 9602
rect 36146 9550 36148 9602
rect 35420 8754 35476 8764
rect 35532 9154 35588 9166
rect 35532 9102 35534 9154
rect 35586 9102 35588 9154
rect 35532 9044 35588 9102
rect 35644 9156 35700 9194
rect 35644 9090 35700 9100
rect 35756 9154 35812 9166
rect 35756 9102 35758 9154
rect 35810 9102 35812 9154
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35420 8484 35476 8494
rect 35420 8146 35476 8428
rect 35420 8094 35422 8146
rect 35474 8094 35476 8146
rect 35420 8082 35476 8094
rect 35532 7812 35588 8988
rect 35756 9044 35812 9102
rect 35756 8146 35812 8988
rect 35980 9042 36036 9054
rect 35980 8990 35982 9042
rect 36034 8990 36036 9042
rect 35756 8094 35758 8146
rect 35810 8094 35812 8146
rect 35756 8082 35812 8094
rect 35868 8930 35924 8942
rect 35868 8878 35870 8930
rect 35922 8878 35924 8930
rect 35868 8036 35924 8878
rect 35980 8260 36036 8990
rect 36092 9044 36148 9550
rect 36092 8978 36148 8988
rect 35980 8166 36036 8204
rect 35868 7970 35924 7980
rect 36092 8148 36148 8158
rect 35532 7756 36036 7812
rect 35420 7588 35476 7598
rect 35420 7362 35476 7532
rect 35756 7588 35812 7598
rect 35420 7310 35422 7362
rect 35474 7310 35476 7362
rect 35420 7298 35476 7310
rect 35532 7474 35588 7486
rect 35532 7422 35534 7474
rect 35586 7422 35588 7474
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 6692 35252 6702
rect 35196 6578 35252 6636
rect 35196 6526 35198 6578
rect 35250 6526 35252 6578
rect 35196 6514 35252 6526
rect 35308 6580 35364 6590
rect 35308 6486 35364 6524
rect 35420 6578 35476 6590
rect 35420 6526 35422 6578
rect 35474 6526 35476 6578
rect 34972 6468 35028 6478
rect 34972 6374 35028 6412
rect 35420 6356 35476 6526
rect 35308 6300 35476 6356
rect 35084 6020 35140 6030
rect 34860 6018 35140 6020
rect 34860 5966 35086 6018
rect 35138 5966 35140 6018
rect 34860 5964 35140 5966
rect 35084 5954 35140 5964
rect 35196 6020 35252 6030
rect 35308 6020 35364 6300
rect 35420 6132 35476 6142
rect 35532 6132 35588 7422
rect 35420 6130 35588 6132
rect 35420 6078 35422 6130
rect 35474 6078 35588 6130
rect 35420 6076 35588 6078
rect 35644 7364 35700 7374
rect 35420 6066 35476 6076
rect 35252 5964 35364 6020
rect 35196 5926 35252 5964
rect 35644 5906 35700 7308
rect 35756 6802 35812 7532
rect 35756 6750 35758 6802
rect 35810 6750 35812 6802
rect 35756 6738 35812 6750
rect 35756 6468 35812 6478
rect 35812 6412 35924 6468
rect 35756 6402 35812 6412
rect 35644 5854 35646 5906
rect 35698 5854 35700 5906
rect 35644 5842 35700 5854
rect 35868 5572 35924 6412
rect 35980 6356 36036 7756
rect 35980 6290 36036 6300
rect 36092 7476 36148 8092
rect 36092 5794 36148 7420
rect 36092 5742 36094 5794
rect 36146 5742 36148 5794
rect 36092 5730 36148 5742
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35644 5516 35924 5572
rect 35644 5346 35700 5516
rect 35644 5294 35646 5346
rect 35698 5294 35700 5346
rect 35644 5282 35700 5294
rect 35980 5348 36036 5358
rect 35980 5254 36036 5292
rect 34972 5124 35028 5134
rect 34972 5030 35028 5068
rect 34860 5012 34916 5022
rect 34860 4918 34916 4956
rect 35980 4900 36036 4910
rect 34636 3390 34638 3442
rect 34690 3390 34692 3442
rect 34300 3378 34356 3388
rect 34636 3378 34692 3390
rect 34972 4676 35028 4686
rect 34972 3554 35028 4620
rect 35980 4450 36036 4844
rect 35980 4398 35982 4450
rect 36034 4398 36036 4450
rect 35980 4386 36036 4398
rect 36092 4564 36148 4574
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 36092 3778 36148 4508
rect 36092 3726 36094 3778
rect 36146 3726 36148 3778
rect 36092 3714 36148 3726
rect 34972 3502 34974 3554
rect 35026 3502 35028 3554
rect 34300 924 34692 980
rect 34300 800 34356 924
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 7392 0 7504 800
rect 29568 0 29680 800
rect 31584 0 31696 800
rect 32256 0 32368 800
rect 32928 0 33040 800
rect 34272 0 34384 800
rect 34636 756 34692 924
rect 34972 756 35028 3502
rect 35532 3442 35588 3454
rect 35532 3390 35534 3442
rect 35586 3390 35588 3442
rect 35532 3332 35588 3390
rect 36204 3388 36260 13692
rect 36316 13522 36372 13534
rect 36316 13470 36318 13522
rect 36370 13470 36372 13522
rect 36316 12068 36372 13470
rect 36540 13524 36596 14364
rect 36652 13748 36708 17948
rect 36764 17106 36820 18620
rect 36876 18610 36932 18620
rect 37436 18450 37492 20636
rect 37436 18398 37438 18450
rect 37490 18398 37492 18450
rect 37436 18386 37492 18398
rect 37548 18228 37604 21980
rect 37884 21474 37940 22204
rect 37884 21422 37886 21474
rect 37938 21422 37940 21474
rect 37884 21410 37940 21422
rect 37996 21140 38052 22652
rect 37996 21074 38052 21084
rect 38108 21700 38164 24108
rect 38220 23380 38276 24780
rect 38892 24834 38948 25228
rect 38892 24782 38894 24834
rect 38946 24782 38948 24834
rect 38668 24724 38724 24762
rect 38668 24658 38724 24668
rect 38220 23314 38276 23324
rect 38556 23772 38836 23828
rect 38332 23156 38388 23166
rect 38556 23156 38612 23772
rect 38332 23154 38612 23156
rect 38332 23102 38334 23154
rect 38386 23102 38612 23154
rect 38332 23100 38612 23102
rect 38668 23604 38724 23614
rect 38332 23044 38388 23100
rect 38332 22978 38388 22988
rect 38668 21812 38724 23548
rect 38780 23492 38836 23772
rect 38892 23492 38948 24782
rect 38780 23436 38948 23492
rect 39004 23938 39060 26236
rect 39116 25618 39172 27022
rect 39116 25566 39118 25618
rect 39170 25566 39172 25618
rect 39116 25554 39172 25566
rect 39228 25508 39284 27580
rect 39452 27634 39508 27646
rect 39452 27582 39454 27634
rect 39506 27582 39508 27634
rect 39452 27412 39508 27582
rect 39452 27346 39508 27356
rect 39900 26514 39956 28252
rect 40012 28084 40068 28094
rect 40012 27970 40068 28028
rect 40012 27918 40014 27970
rect 40066 27918 40068 27970
rect 40012 27906 40068 27918
rect 40124 27972 40180 27982
rect 40124 27858 40180 27916
rect 40124 27806 40126 27858
rect 40178 27806 40180 27858
rect 40124 27794 40180 27806
rect 40236 26964 40292 28812
rect 40684 28802 40740 28812
rect 40796 28868 40852 29934
rect 41356 29876 41412 30156
rect 41468 30212 41524 31166
rect 41692 30772 41748 32060
rect 41804 30994 41860 35084
rect 41916 35074 41972 35084
rect 42028 34804 42084 34814
rect 41916 34690 41972 34702
rect 41916 34638 41918 34690
rect 41970 34638 41972 34690
rect 41916 34130 41972 34638
rect 41916 34078 41918 34130
rect 41970 34078 41972 34130
rect 41916 34066 41972 34078
rect 42028 34356 42084 34748
rect 42140 34356 42196 35532
rect 42476 35522 42532 35532
rect 42252 34916 42308 34926
rect 42252 34914 42420 34916
rect 42252 34862 42254 34914
rect 42306 34862 42420 34914
rect 42252 34860 42420 34862
rect 42252 34850 42308 34860
rect 42364 34580 42420 34860
rect 42476 34804 42532 34814
rect 42588 34804 42644 38612
rect 42924 38612 42980 38670
rect 42924 38546 42980 38556
rect 42812 38500 42868 38510
rect 42700 38276 42756 38286
rect 42700 38182 42756 38220
rect 42700 38052 42756 38062
rect 42700 37958 42756 37996
rect 42700 37042 42756 37054
rect 42700 36990 42702 37042
rect 42754 36990 42756 37042
rect 42700 36596 42756 36990
rect 42700 36530 42756 36540
rect 42812 36372 42868 38444
rect 42700 36316 42868 36372
rect 43036 38164 43092 39116
rect 43484 38836 43540 38846
rect 43036 38108 43428 38164
rect 43036 37938 43092 38108
rect 43036 37886 43038 37938
rect 43090 37886 43092 37938
rect 42700 34916 42756 36316
rect 42924 36260 42980 36270
rect 42812 36148 42868 36158
rect 42812 35698 42868 36092
rect 42924 35922 42980 36204
rect 42924 35870 42926 35922
rect 42978 35870 42980 35922
rect 42924 35858 42980 35870
rect 42812 35646 42814 35698
rect 42866 35646 42868 35698
rect 42812 35634 42868 35646
rect 42924 35476 42980 35486
rect 42700 34850 42756 34860
rect 42812 35364 42868 35374
rect 42812 34914 42868 35308
rect 42812 34862 42814 34914
rect 42866 34862 42868 34914
rect 42812 34850 42868 34862
rect 42532 34748 42644 34804
rect 42924 34802 42980 35420
rect 42924 34750 42926 34802
rect 42978 34750 42980 34802
rect 42476 34738 42532 34748
rect 42924 34738 42980 34750
rect 42812 34692 42868 34702
rect 42364 34524 42756 34580
rect 42140 34300 42420 34356
rect 42028 32564 42084 34300
rect 42140 34132 42196 34170
rect 42140 34066 42196 34076
rect 42252 34018 42308 34030
rect 42252 33966 42254 34018
rect 42306 33966 42308 34018
rect 42028 32498 42084 32508
rect 42140 33908 42196 33918
rect 42140 31668 42196 33852
rect 42252 33234 42308 33966
rect 42252 33182 42254 33234
rect 42306 33182 42308 33234
rect 42252 33170 42308 33182
rect 42364 32674 42420 34300
rect 42700 34354 42756 34524
rect 42700 34302 42702 34354
rect 42754 34302 42756 34354
rect 42700 34290 42756 34302
rect 42588 34244 42644 34254
rect 42588 34150 42644 34188
rect 42812 34130 42868 34636
rect 42812 34078 42814 34130
rect 42866 34078 42868 34130
rect 42812 34066 42868 34078
rect 43036 33236 43092 37886
rect 43260 37938 43316 37950
rect 43260 37886 43262 37938
rect 43314 37886 43316 37938
rect 43148 37828 43204 37838
rect 43148 37734 43204 37772
rect 43260 37380 43316 37886
rect 43148 37324 43316 37380
rect 43372 37378 43428 38108
rect 43484 37490 43540 38780
rect 43596 38500 43652 39342
rect 43596 38434 43652 38444
rect 43484 37438 43486 37490
rect 43538 37438 43540 37490
rect 43484 37426 43540 37438
rect 43596 38276 43652 38286
rect 43372 37326 43374 37378
rect 43426 37326 43428 37378
rect 43148 37266 43204 37324
rect 43372 37314 43428 37326
rect 43148 37214 43150 37266
rect 43202 37214 43204 37266
rect 43148 35924 43204 37214
rect 43596 37266 43652 38220
rect 43932 38162 43988 38174
rect 43932 38110 43934 38162
rect 43986 38110 43988 38162
rect 43820 38050 43876 38062
rect 43820 37998 43822 38050
rect 43874 37998 43876 38050
rect 43596 37214 43598 37266
rect 43650 37214 43652 37266
rect 43596 37202 43652 37214
rect 43708 37940 43764 37950
rect 43708 37266 43764 37884
rect 43820 37828 43876 37998
rect 43820 37762 43876 37772
rect 43708 37214 43710 37266
rect 43762 37214 43764 37266
rect 43708 37202 43764 37214
rect 43708 37044 43764 37054
rect 43596 36484 43652 36494
rect 43484 35924 43540 35934
rect 43148 35868 43316 35924
rect 43148 35700 43204 35710
rect 43148 34242 43204 35644
rect 43148 34190 43150 34242
rect 43202 34190 43204 34242
rect 43148 34178 43204 34190
rect 43148 33236 43204 33246
rect 43036 33180 43148 33236
rect 43148 33170 43204 33180
rect 43260 33012 43316 35868
rect 43484 35698 43540 35868
rect 43484 35646 43486 35698
rect 43538 35646 43540 35698
rect 43484 35634 43540 35646
rect 43596 35140 43652 36428
rect 43708 35810 43764 36988
rect 43932 36370 43988 38110
rect 43932 36318 43934 36370
rect 43986 36318 43988 36370
rect 43932 36306 43988 36318
rect 43708 35758 43710 35810
rect 43762 35758 43764 35810
rect 43708 35746 43764 35758
rect 43932 35924 43988 35934
rect 42364 32622 42366 32674
rect 42418 32622 42420 32674
rect 42364 32610 42420 32622
rect 43036 32956 43316 33012
rect 43372 35084 43652 35140
rect 42252 32562 42308 32574
rect 42700 32564 42756 32574
rect 42252 32510 42254 32562
rect 42306 32510 42308 32562
rect 42252 32004 42308 32510
rect 42252 31938 42308 31948
rect 42588 32562 42756 32564
rect 42588 32510 42702 32562
rect 42754 32510 42756 32562
rect 42588 32508 42756 32510
rect 42140 31602 42196 31612
rect 42252 31780 42308 31790
rect 42252 31666 42308 31724
rect 42252 31614 42254 31666
rect 42306 31614 42308 31666
rect 42252 31602 42308 31614
rect 41804 30942 41806 30994
rect 41858 30942 41860 30994
rect 41804 30930 41860 30942
rect 41916 31444 41972 31454
rect 41692 30716 41860 30772
rect 41468 30210 41636 30212
rect 41468 30158 41470 30210
rect 41522 30158 41636 30210
rect 41468 30156 41636 30158
rect 41468 30146 41524 30156
rect 41356 29820 41524 29876
rect 41356 29652 41412 29662
rect 41244 29428 41300 29438
rect 41020 29316 41076 29326
rect 41020 29314 41188 29316
rect 41020 29262 41022 29314
rect 41074 29262 41188 29314
rect 41020 29260 41188 29262
rect 41020 29250 41076 29260
rect 40852 28812 41076 28868
rect 40796 28802 40852 28812
rect 40348 28642 40404 28654
rect 40348 28590 40350 28642
rect 40402 28590 40404 28642
rect 40348 28532 40404 28590
rect 40348 28476 40852 28532
rect 40460 28196 40516 28206
rect 39900 26462 39902 26514
rect 39954 26462 39956 26514
rect 39900 26450 39956 26462
rect 40012 26962 40292 26964
rect 40012 26910 40238 26962
rect 40290 26910 40292 26962
rect 40012 26908 40292 26910
rect 39676 26404 39732 26414
rect 39452 26292 39508 26302
rect 39452 26198 39508 26236
rect 39676 26290 39732 26348
rect 40012 26404 40068 26908
rect 40236 26898 40292 26908
rect 40348 27412 40404 27422
rect 40348 26740 40404 27356
rect 40124 26684 40404 26740
rect 40124 26514 40180 26684
rect 40460 26628 40516 28140
rect 40796 27748 40852 28476
rect 41020 27970 41076 28812
rect 41132 28420 41188 29260
rect 41244 28756 41300 29372
rect 41356 29204 41412 29596
rect 41468 29650 41524 29820
rect 41468 29598 41470 29650
rect 41522 29598 41524 29650
rect 41468 29586 41524 29598
rect 41356 29148 41524 29204
rect 41244 28690 41300 28700
rect 41356 28644 41412 28654
rect 41356 28530 41412 28588
rect 41356 28478 41358 28530
rect 41410 28478 41412 28530
rect 41356 28466 41412 28478
rect 41468 28642 41524 29148
rect 41468 28590 41470 28642
rect 41522 28590 41524 28642
rect 41244 28420 41300 28430
rect 41132 28364 41244 28420
rect 41020 27918 41022 27970
rect 41074 27918 41076 27970
rect 41020 27906 41076 27918
rect 41132 27858 41188 27870
rect 41132 27806 41134 27858
rect 41186 27806 41188 27858
rect 41132 27748 41188 27806
rect 40796 27692 41188 27748
rect 40908 27300 40964 27310
rect 40460 26562 40516 26572
rect 40684 27074 40740 27086
rect 40684 27022 40686 27074
rect 40738 27022 40740 27074
rect 40124 26462 40126 26514
rect 40178 26462 40180 26514
rect 40124 26450 40180 26462
rect 40012 26338 40068 26348
rect 39676 26238 39678 26290
rect 39730 26238 39732 26290
rect 39676 26226 39732 26238
rect 40124 26292 40180 26302
rect 40180 26236 40292 26292
rect 40124 26226 40180 26236
rect 40012 26178 40068 26190
rect 40012 26126 40014 26178
rect 40066 26126 40068 26178
rect 39564 25508 39620 25518
rect 39228 25506 39620 25508
rect 39228 25454 39566 25506
rect 39618 25454 39620 25506
rect 39228 25452 39620 25454
rect 39116 25396 39172 25406
rect 39116 24164 39172 25340
rect 39340 24722 39396 25452
rect 39564 25442 39620 25452
rect 39340 24670 39342 24722
rect 39394 24670 39396 24722
rect 39340 24658 39396 24670
rect 39676 24276 39732 24286
rect 39228 24164 39284 24174
rect 39116 24162 39284 24164
rect 39116 24110 39230 24162
rect 39282 24110 39284 24162
rect 39116 24108 39284 24110
rect 39004 23886 39006 23938
rect 39058 23886 39060 23938
rect 39004 23492 39060 23886
rect 39004 23426 39060 23436
rect 39116 23266 39172 23278
rect 39116 23214 39118 23266
rect 39170 23214 39172 23266
rect 39004 23154 39060 23166
rect 39004 23102 39006 23154
rect 39058 23102 39060 23154
rect 39004 22596 39060 23102
rect 39116 22820 39172 23214
rect 39116 22754 39172 22764
rect 39228 22708 39284 24108
rect 39340 23938 39396 23950
rect 39340 23886 39342 23938
rect 39394 23886 39396 23938
rect 39340 22932 39396 23886
rect 39564 23156 39620 23166
rect 39564 23062 39620 23100
rect 39340 22866 39396 22876
rect 39228 22652 39620 22708
rect 39004 22594 39508 22596
rect 39004 22542 39006 22594
rect 39058 22542 39508 22594
rect 39004 22540 39508 22542
rect 39004 22530 39060 22540
rect 39452 22370 39508 22540
rect 39452 22318 39454 22370
rect 39506 22318 39508 22370
rect 39452 22306 39508 22318
rect 39564 22372 39620 22652
rect 39564 22306 39620 22316
rect 39340 22148 39396 22158
rect 39228 22092 39340 22148
rect 38668 21756 38948 21812
rect 38108 21644 38612 21700
rect 38108 20802 38164 21644
rect 38556 21588 38612 21644
rect 38668 21588 38724 21598
rect 38556 21586 38724 21588
rect 38556 21534 38670 21586
rect 38722 21534 38724 21586
rect 38556 21532 38724 21534
rect 38668 21522 38724 21532
rect 38108 20750 38110 20802
rect 38162 20750 38164 20802
rect 38108 20738 38164 20750
rect 38220 21474 38276 21486
rect 38220 21422 38222 21474
rect 38274 21422 38276 21474
rect 37772 20132 37828 20142
rect 37436 18172 37604 18228
rect 37660 20020 37716 20030
rect 36988 18116 37044 18126
rect 36988 17666 37044 18060
rect 36988 17614 36990 17666
rect 37042 17614 37044 17666
rect 36988 17444 37044 17614
rect 36988 17378 37044 17388
rect 36764 17054 36766 17106
rect 36818 17054 36820 17106
rect 36764 17042 36820 17054
rect 37212 16994 37268 17006
rect 37212 16942 37214 16994
rect 37266 16942 37268 16994
rect 37212 16212 37268 16942
rect 37436 16436 37492 18172
rect 37548 17668 37604 17678
rect 37660 17668 37716 19964
rect 37548 17666 37716 17668
rect 37548 17614 37550 17666
rect 37602 17614 37716 17666
rect 37548 17612 37716 17614
rect 37548 17602 37604 17612
rect 37548 16884 37604 16894
rect 37548 16882 37716 16884
rect 37548 16830 37550 16882
rect 37602 16830 37716 16882
rect 37548 16828 37716 16830
rect 37548 16818 37604 16828
rect 37548 16436 37604 16446
rect 37436 16380 37548 16436
rect 37548 16370 37604 16380
rect 36988 16156 37268 16212
rect 36988 16100 37044 16156
rect 36876 16044 37044 16100
rect 37548 16100 37604 16110
rect 36876 15148 36932 16044
rect 37100 15986 37156 15998
rect 37100 15934 37102 15986
rect 37154 15934 37156 15986
rect 36988 15876 37044 15886
rect 36988 15782 37044 15820
rect 36764 15092 36932 15148
rect 37100 15148 37156 15934
rect 37548 15316 37604 16044
rect 37660 15540 37716 16828
rect 37772 16212 37828 20076
rect 38220 19236 38276 21422
rect 37996 19180 38276 19236
rect 38444 20914 38500 20926
rect 38444 20862 38446 20914
rect 38498 20862 38500 20914
rect 37996 17892 38052 19180
rect 37996 17826 38052 17836
rect 38108 19012 38164 19022
rect 37884 17780 37940 17790
rect 37884 17686 37940 17724
rect 38108 17668 38164 18956
rect 38332 18676 38388 18686
rect 38220 18340 38276 18350
rect 38220 18246 38276 18284
rect 38220 17668 38276 17678
rect 38108 17666 38276 17668
rect 38108 17614 38222 17666
rect 38274 17614 38276 17666
rect 38108 17612 38276 17614
rect 37884 16884 37940 16894
rect 37884 16790 37940 16828
rect 38108 16660 38164 16670
rect 38220 16660 38276 17612
rect 38108 16658 38276 16660
rect 38108 16606 38110 16658
rect 38162 16606 38276 16658
rect 38108 16604 38276 16606
rect 38332 16660 38388 18620
rect 38444 18004 38500 20862
rect 38556 20244 38612 20254
rect 38556 19122 38612 20188
rect 38892 19684 38948 21756
rect 39116 21700 39172 21710
rect 39116 21586 39172 21644
rect 39116 21534 39118 21586
rect 39170 21534 39172 21586
rect 39004 20804 39060 20814
rect 39116 20804 39172 21534
rect 39004 20802 39172 20804
rect 39004 20750 39006 20802
rect 39058 20750 39172 20802
rect 39004 20748 39172 20750
rect 39004 20468 39060 20748
rect 39004 20402 39060 20412
rect 39116 20018 39172 20030
rect 39116 19966 39118 20018
rect 39170 19966 39172 20018
rect 39116 19908 39172 19966
rect 38892 19628 39060 19684
rect 38556 19070 38558 19122
rect 38610 19070 38612 19122
rect 38556 19058 38612 19070
rect 38444 17948 38612 18004
rect 38444 17780 38500 17790
rect 38444 17554 38500 17724
rect 38444 17502 38446 17554
rect 38498 17502 38500 17554
rect 38444 16884 38500 17502
rect 38444 16818 38500 16828
rect 38444 16660 38500 16670
rect 38332 16658 38500 16660
rect 38332 16606 38446 16658
rect 38498 16606 38500 16658
rect 38332 16604 38500 16606
rect 38108 16594 38164 16604
rect 38444 16594 38500 16604
rect 38332 16436 38388 16446
rect 38556 16436 38612 17948
rect 39004 17668 39060 19628
rect 39116 19236 39172 19852
rect 39116 19170 39172 19180
rect 37772 16156 37940 16212
rect 37772 15988 37828 15998
rect 37772 15894 37828 15932
rect 37660 15446 37716 15484
rect 37548 15250 37604 15260
rect 37100 15092 37268 15148
rect 36764 14196 36820 15092
rect 37100 15026 37156 15036
rect 37100 14756 37156 14766
rect 37100 14644 37156 14700
rect 36764 14130 36820 14140
rect 36876 14642 37156 14644
rect 36876 14590 37102 14642
rect 37154 14590 37156 14642
rect 36876 14588 37156 14590
rect 36876 13748 36932 14588
rect 37100 14578 37156 14588
rect 37212 13970 37268 15092
rect 37212 13918 37214 13970
rect 37266 13918 37268 13970
rect 37212 13906 37268 13918
rect 37324 15090 37380 15102
rect 37324 15038 37326 15090
rect 37378 15038 37380 15090
rect 37324 13972 37380 15038
rect 37548 14532 37604 14542
rect 37548 14438 37604 14476
rect 37324 13916 37716 13972
rect 36652 13692 36820 13748
rect 36652 13524 36708 13534
rect 36540 13522 36708 13524
rect 36540 13470 36654 13522
rect 36706 13470 36708 13522
rect 36540 13468 36708 13470
rect 36764 13524 36820 13692
rect 36876 13654 36932 13692
rect 37548 13746 37604 13758
rect 37548 13694 37550 13746
rect 37602 13694 37604 13746
rect 36764 13468 36932 13524
rect 36652 13412 36708 13468
rect 36652 13346 36708 13356
rect 36316 12002 36372 12012
rect 36428 11172 36484 11182
rect 36428 11170 36820 11172
rect 36428 11118 36430 11170
rect 36482 11118 36820 11170
rect 36428 11116 36820 11118
rect 36428 11106 36484 11116
rect 36764 10836 36820 11116
rect 36764 10742 36820 10780
rect 36876 10164 36932 13468
rect 37436 12962 37492 12974
rect 37436 12910 37438 12962
rect 37490 12910 37492 12962
rect 37100 12738 37156 12750
rect 37100 12686 37102 12738
rect 37154 12686 37156 12738
rect 36988 12292 37044 12302
rect 36988 11506 37044 12236
rect 37100 12180 37156 12686
rect 37436 12516 37492 12910
rect 37548 12852 37604 13694
rect 37660 13636 37716 13916
rect 37884 13860 37940 16156
rect 38108 15986 38164 15998
rect 38108 15934 38110 15986
rect 38162 15934 38164 15986
rect 38108 15540 38164 15934
rect 37996 14308 38052 14318
rect 37996 14214 38052 14252
rect 37884 13804 38052 13860
rect 37884 13636 37940 13646
rect 37660 13634 37940 13636
rect 37660 13582 37886 13634
rect 37938 13582 37940 13634
rect 37660 13580 37940 13582
rect 37884 13076 37940 13580
rect 37996 13076 38052 13804
rect 38108 13746 38164 15484
rect 38220 15874 38276 15886
rect 38220 15822 38222 15874
rect 38274 15822 38276 15874
rect 38220 14532 38276 15822
rect 38220 14466 38276 14476
rect 38108 13694 38110 13746
rect 38162 13694 38164 13746
rect 38108 13682 38164 13694
rect 37996 13020 38276 13076
rect 37884 13010 37940 13020
rect 37660 12852 37716 12862
rect 37548 12850 37716 12852
rect 37548 12798 37662 12850
rect 37714 12798 37716 12850
rect 37548 12796 37716 12798
rect 37436 12450 37492 12460
rect 37324 12180 37380 12190
rect 37100 12178 37380 12180
rect 37100 12126 37326 12178
rect 37378 12126 37380 12178
rect 37100 12124 37380 12126
rect 36988 11454 36990 11506
rect 37042 11454 37044 11506
rect 36988 11442 37044 11454
rect 37212 11508 37268 11518
rect 37212 11414 37268 11452
rect 37324 10948 37380 12124
rect 37660 11844 37716 12796
rect 37996 12850 38052 12862
rect 37996 12798 37998 12850
rect 38050 12798 38052 12850
rect 37996 12404 38052 12798
rect 37996 12338 38052 12348
rect 38108 12516 38164 12526
rect 37884 12180 37940 12190
rect 37660 11778 37716 11788
rect 37772 12178 37940 12180
rect 37772 12126 37886 12178
rect 37938 12126 37940 12178
rect 37772 12124 37940 12126
rect 37548 11620 37604 11630
rect 37772 11620 37828 12124
rect 37884 12114 37940 12124
rect 38108 12068 38164 12460
rect 37548 11618 37828 11620
rect 37548 11566 37550 11618
rect 37602 11566 37828 11618
rect 37548 11564 37828 11566
rect 37996 12012 38164 12068
rect 37548 11554 37604 11564
rect 36876 10098 36932 10108
rect 36988 10892 37380 10948
rect 36540 9828 36596 9838
rect 36540 9042 36596 9772
rect 36988 9604 37044 10892
rect 37996 10722 38052 12012
rect 38108 11844 38164 11854
rect 38108 11618 38164 11788
rect 38220 11788 38276 13020
rect 38332 12402 38388 16380
rect 38444 16380 38612 16436
rect 38668 17612 39060 17668
rect 38444 15148 38500 16380
rect 38556 16100 38612 16110
rect 38556 16006 38612 16044
rect 38668 15316 38724 17612
rect 38892 17442 38948 17454
rect 38892 17390 38894 17442
rect 38946 17390 38948 17442
rect 38892 17220 38948 17390
rect 38892 17154 38948 17164
rect 38892 16996 38948 17006
rect 38780 16994 38948 16996
rect 38780 16942 38894 16994
rect 38946 16942 38948 16994
rect 38780 16940 38948 16942
rect 38780 15988 38836 16940
rect 38892 16930 38948 16940
rect 39004 16994 39060 17612
rect 39228 17108 39284 22092
rect 39340 22082 39396 22092
rect 39452 21700 39508 21710
rect 39452 20916 39508 21644
rect 39676 21700 39732 24220
rect 39788 23938 39844 23950
rect 39788 23886 39790 23938
rect 39842 23886 39844 23938
rect 39788 23492 39844 23886
rect 40012 23940 40068 26126
rect 40124 25508 40180 25518
rect 40124 24498 40180 25452
rect 40236 24834 40292 26236
rect 40684 25620 40740 27022
rect 40684 25554 40740 25564
rect 40908 26964 40964 27244
rect 41132 27188 41188 27692
rect 41132 27122 41188 27132
rect 41020 26964 41076 26974
rect 40908 26962 41076 26964
rect 40908 26910 41022 26962
rect 41074 26910 41076 26962
rect 40908 26908 41076 26910
rect 40236 24782 40238 24834
rect 40290 24782 40292 24834
rect 40236 24770 40292 24782
rect 40124 24446 40126 24498
rect 40178 24446 40180 24498
rect 40124 24434 40180 24446
rect 40348 24164 40404 24174
rect 40124 24052 40180 24062
rect 40348 24052 40404 24108
rect 40124 24050 40404 24052
rect 40124 23998 40126 24050
rect 40178 23998 40404 24050
rect 40124 23996 40404 23998
rect 40124 23986 40180 23996
rect 40012 23874 40068 23884
rect 39788 22484 39844 23436
rect 39900 23716 39956 23726
rect 39900 22708 39956 23660
rect 40236 23716 40292 23726
rect 40124 23380 40180 23390
rect 40012 23266 40068 23278
rect 40012 23214 40014 23266
rect 40066 23214 40068 23266
rect 40012 22932 40068 23214
rect 40012 22866 40068 22876
rect 39900 22652 40068 22708
rect 39788 22482 39956 22484
rect 39788 22430 39790 22482
rect 39842 22430 39956 22482
rect 39788 22428 39956 22430
rect 39788 22418 39844 22428
rect 39676 21698 39844 21700
rect 39676 21646 39678 21698
rect 39730 21646 39844 21698
rect 39676 21644 39844 21646
rect 39676 21634 39732 21644
rect 39004 16942 39006 16994
rect 39058 16942 39060 16994
rect 39004 16930 39060 16942
rect 39116 17052 39284 17108
rect 39340 20914 39508 20916
rect 39340 20862 39454 20914
rect 39506 20862 39508 20914
rect 39340 20860 39508 20862
rect 38892 16772 38948 16782
rect 39116 16772 39172 17052
rect 38892 16658 38948 16716
rect 38892 16606 38894 16658
rect 38946 16606 38948 16658
rect 38892 16594 38948 16606
rect 39004 16716 39172 16772
rect 39228 16882 39284 16894
rect 39228 16830 39230 16882
rect 39282 16830 39284 16882
rect 39228 16772 39284 16830
rect 38780 15538 38836 15932
rect 39004 15540 39060 16716
rect 39228 16706 39284 16716
rect 39340 16548 39396 20860
rect 39452 20850 39508 20860
rect 39452 20018 39508 20030
rect 39452 19966 39454 20018
rect 39506 19966 39508 20018
rect 39452 18676 39508 19966
rect 39452 18610 39508 18620
rect 39564 18340 39620 18350
rect 39564 17890 39620 18284
rect 39564 17838 39566 17890
rect 39618 17838 39620 17890
rect 39564 17826 39620 17838
rect 39452 17556 39508 17566
rect 39452 17462 39508 17500
rect 39676 17554 39732 17566
rect 39676 17502 39678 17554
rect 39730 17502 39732 17554
rect 39676 17220 39732 17502
rect 39452 17164 39732 17220
rect 39452 16660 39508 17164
rect 39788 16996 39844 21644
rect 39900 21588 39956 22428
rect 40012 22148 40068 22652
rect 40012 22082 40068 22092
rect 40012 21812 40068 21822
rect 40124 21812 40180 23324
rect 40236 23378 40292 23660
rect 40236 23326 40238 23378
rect 40290 23326 40292 23378
rect 40236 23314 40292 23326
rect 40348 23156 40404 23996
rect 40348 23154 40516 23156
rect 40348 23102 40350 23154
rect 40402 23102 40516 23154
rect 40348 23100 40516 23102
rect 40348 23090 40404 23100
rect 40012 21810 40124 21812
rect 40012 21758 40014 21810
rect 40066 21758 40124 21810
rect 40012 21756 40124 21758
rect 40012 21746 40068 21756
rect 40124 21718 40180 21756
rect 40236 21588 40292 21598
rect 39900 21586 40292 21588
rect 39900 21534 40238 21586
rect 40290 21534 40292 21586
rect 39900 21532 40292 21534
rect 40236 21522 40292 21532
rect 39900 21140 39956 21150
rect 39956 21084 40068 21140
rect 39900 21074 39956 21084
rect 39900 20130 39956 20142
rect 39900 20078 39902 20130
rect 39954 20078 39956 20130
rect 39900 19460 39956 20078
rect 39900 19394 39956 19404
rect 40012 18788 40068 21084
rect 40124 20802 40180 20814
rect 40124 20750 40126 20802
rect 40178 20750 40180 20802
rect 40124 20244 40180 20750
rect 40348 20578 40404 20590
rect 40348 20526 40350 20578
rect 40402 20526 40404 20578
rect 40348 20356 40404 20526
rect 40348 20290 40404 20300
rect 40124 20178 40180 20188
rect 40348 19572 40404 19582
rect 40236 19348 40292 19358
rect 40236 19122 40292 19292
rect 40236 19070 40238 19122
rect 40290 19070 40292 19122
rect 40236 19058 40292 19070
rect 40012 18732 40292 18788
rect 40012 18340 40068 18350
rect 40012 17890 40068 18284
rect 40236 18116 40292 18732
rect 40348 18338 40404 19516
rect 40348 18286 40350 18338
rect 40402 18286 40404 18338
rect 40348 18274 40404 18286
rect 40236 18060 40404 18116
rect 40012 17838 40014 17890
rect 40066 17838 40068 17890
rect 40012 17826 40068 17838
rect 40236 17668 40292 17678
rect 40124 17666 40292 17668
rect 40124 17614 40238 17666
rect 40290 17614 40292 17666
rect 40124 17612 40292 17614
rect 39900 17556 39956 17566
rect 39956 17500 40068 17556
rect 39900 17490 39956 17500
rect 39676 16940 39844 16996
rect 39676 16882 39732 16940
rect 39676 16830 39678 16882
rect 39730 16830 39732 16882
rect 39676 16772 39732 16830
rect 39900 16884 39956 16894
rect 39900 16790 39956 16828
rect 39676 16706 39732 16716
rect 39788 16770 39844 16782
rect 39788 16718 39790 16770
rect 39842 16718 39844 16770
rect 39452 16594 39508 16604
rect 38780 15486 38782 15538
rect 38834 15486 38836 15538
rect 38780 15474 38836 15486
rect 38892 15484 39060 15540
rect 39116 16492 39396 16548
rect 38668 15260 38836 15316
rect 38444 15092 38612 15148
rect 38444 14530 38500 14542
rect 38444 14478 38446 14530
rect 38498 14478 38500 14530
rect 38444 13970 38500 14478
rect 38444 13918 38446 13970
rect 38498 13918 38500 13970
rect 38444 13906 38500 13918
rect 38332 12350 38334 12402
rect 38386 12350 38388 12402
rect 38332 12338 38388 12350
rect 38444 13076 38500 13086
rect 38444 12292 38500 13020
rect 38220 11732 38388 11788
rect 38108 11566 38110 11618
rect 38162 11566 38164 11618
rect 38108 11554 38164 11566
rect 37996 10670 37998 10722
rect 38050 10670 38052 10722
rect 37996 10658 38052 10670
rect 38220 10836 38276 10846
rect 38220 10050 38276 10780
rect 38220 9998 38222 10050
rect 38274 9998 38276 10050
rect 38220 9986 38276 9998
rect 37884 9940 37940 9950
rect 37660 9938 37940 9940
rect 37660 9886 37886 9938
rect 37938 9886 37940 9938
rect 37660 9884 37940 9886
rect 37212 9828 37268 9838
rect 37212 9734 37268 9772
rect 37660 9826 37716 9884
rect 37660 9774 37662 9826
rect 37714 9774 37716 9826
rect 37660 9762 37716 9774
rect 36540 8990 36542 9042
rect 36594 8990 36596 9042
rect 36540 8978 36596 8990
rect 36876 9602 37044 9604
rect 36876 9550 36990 9602
rect 37042 9550 37044 9602
rect 36876 9548 37044 9550
rect 36876 8930 36932 9548
rect 36988 9538 37044 9548
rect 37100 9602 37156 9614
rect 37100 9550 37102 9602
rect 37154 9550 37156 9602
rect 36876 8878 36878 8930
rect 36930 8878 36932 8930
rect 36876 8866 36932 8878
rect 36988 9156 37044 9166
rect 36988 8818 37044 9100
rect 36988 8766 36990 8818
rect 37042 8766 37044 8818
rect 36988 8258 37044 8766
rect 37100 8484 37156 9550
rect 37100 8418 37156 8428
rect 37548 9156 37604 9166
rect 37548 8820 37604 9100
rect 37884 9154 37940 9884
rect 37884 9102 37886 9154
rect 37938 9102 37940 9154
rect 37884 9090 37940 9102
rect 37772 9044 37828 9054
rect 37772 8820 37828 8988
rect 37772 8764 38164 8820
rect 37212 8372 37268 8382
rect 37212 8278 37268 8316
rect 36988 8206 36990 8258
rect 37042 8206 37044 8258
rect 36988 8194 37044 8206
rect 37324 8258 37380 8270
rect 37324 8206 37326 8258
rect 37378 8206 37380 8258
rect 36316 8034 36372 8046
rect 36316 7982 36318 8034
rect 36370 7982 36372 8034
rect 36316 7476 36372 7982
rect 36316 7382 36372 7420
rect 36428 6580 36484 6590
rect 36988 6580 37044 6590
rect 36428 6578 36932 6580
rect 36428 6526 36430 6578
rect 36482 6526 36932 6578
rect 36428 6524 36932 6526
rect 36428 6514 36484 6524
rect 36316 6466 36372 6478
rect 36316 6414 36318 6466
rect 36370 6414 36372 6466
rect 36316 6356 36372 6414
rect 36316 5908 36372 6300
rect 36316 5842 36372 5852
rect 36876 4564 36932 6524
rect 36988 5234 37044 6524
rect 36988 5182 36990 5234
rect 37042 5182 37044 5234
rect 36988 4900 37044 5182
rect 37324 6020 37380 8206
rect 37044 4844 37268 4900
rect 36988 4834 37044 4844
rect 36876 4470 36932 4508
rect 37212 3442 37268 4844
rect 37324 4226 37380 5964
rect 37436 7252 37492 7262
rect 37436 4452 37492 7196
rect 37436 4386 37492 4396
rect 37548 6690 37604 8764
rect 37996 8370 38052 8382
rect 37996 8318 37998 8370
rect 38050 8318 38052 8370
rect 37996 8260 38052 8318
rect 37884 8204 37996 8260
rect 37884 6804 37940 8204
rect 37996 8194 38052 8204
rect 38108 8258 38164 8764
rect 38108 8206 38110 8258
rect 38162 8206 38164 8258
rect 38108 8194 38164 8206
rect 37884 6738 37940 6748
rect 38108 7474 38164 7486
rect 38108 7422 38110 7474
rect 38162 7422 38164 7474
rect 37548 6638 37550 6690
rect 37602 6638 37604 6690
rect 37548 4340 37604 6638
rect 38108 6020 38164 7422
rect 38108 5954 38164 5964
rect 38220 7476 38276 7486
rect 38220 5794 38276 7420
rect 38220 5742 38222 5794
rect 38274 5742 38276 5794
rect 38220 5730 38276 5742
rect 38332 5572 38388 11732
rect 38444 9938 38500 12236
rect 38444 9886 38446 9938
rect 38498 9886 38500 9938
rect 38444 9874 38500 9886
rect 38556 9604 38612 15092
rect 38668 13076 38724 13086
rect 38668 12982 38724 13020
rect 38780 12852 38836 15260
rect 38892 14420 38948 15484
rect 38892 14354 38948 14364
rect 39004 15316 39060 15326
rect 38892 14196 38948 14206
rect 38892 13186 38948 14140
rect 38892 13134 38894 13186
rect 38946 13134 38948 13186
rect 38892 13122 38948 13134
rect 38668 12796 38836 12852
rect 38668 11732 38724 12796
rect 39004 12516 39060 15260
rect 39116 14980 39172 16492
rect 39788 16324 39844 16718
rect 39340 16268 39844 16324
rect 39340 16210 39396 16268
rect 39340 16158 39342 16210
rect 39394 16158 39396 16210
rect 39340 16146 39396 16158
rect 39116 14914 39172 14924
rect 39228 16100 39284 16110
rect 39228 14756 39284 16044
rect 40012 15652 40068 17500
rect 40124 15876 40180 17612
rect 40236 17602 40292 17612
rect 40348 17106 40404 18060
rect 40348 17054 40350 17106
rect 40402 17054 40404 17106
rect 40348 17042 40404 17054
rect 40460 16884 40516 23100
rect 40572 22820 40628 22830
rect 40572 20802 40628 22764
rect 40684 22372 40740 22382
rect 40684 22278 40740 22316
rect 40908 22260 40964 26908
rect 41020 26898 41076 26908
rect 41132 26402 41188 26414
rect 41132 26350 41134 26402
rect 41186 26350 41188 26402
rect 41020 26290 41076 26302
rect 41020 26238 41022 26290
rect 41074 26238 41076 26290
rect 41020 25284 41076 26238
rect 41020 25218 41076 25228
rect 41020 24948 41076 24958
rect 41020 24854 41076 24892
rect 41132 23380 41188 26350
rect 41132 23314 41188 23324
rect 41020 22932 41076 22942
rect 41020 22838 41076 22876
rect 40572 20750 40574 20802
rect 40626 20750 40628 20802
rect 40572 20738 40628 20750
rect 40796 22258 40964 22260
rect 40796 22206 40910 22258
rect 40962 22206 40964 22258
rect 40796 22204 40964 22206
rect 40796 20690 40852 22204
rect 40908 22194 40964 22204
rect 41020 22372 41076 22382
rect 41020 22036 41076 22316
rect 40908 21980 41076 22036
rect 40908 20802 40964 21980
rect 41020 21812 41076 21822
rect 41020 21586 41076 21756
rect 41244 21588 41300 28364
rect 41468 27972 41524 28590
rect 41580 28084 41636 30156
rect 41580 28018 41636 28028
rect 41468 27074 41524 27916
rect 41580 27746 41636 27758
rect 41580 27694 41582 27746
rect 41634 27694 41636 27746
rect 41580 27636 41636 27694
rect 41692 27748 41748 27758
rect 41692 27654 41748 27692
rect 41580 27570 41636 27580
rect 41692 27412 41748 27422
rect 41692 27186 41748 27356
rect 41692 27134 41694 27186
rect 41746 27134 41748 27186
rect 41692 27122 41748 27134
rect 41468 27022 41470 27074
rect 41522 27022 41524 27074
rect 41468 27010 41524 27022
rect 41692 26180 41748 26190
rect 41692 26086 41748 26124
rect 41356 25620 41412 25630
rect 41356 25506 41412 25564
rect 41356 25454 41358 25506
rect 41410 25454 41412 25506
rect 41356 25442 41412 25454
rect 41692 25508 41748 25518
rect 41692 25414 41748 25452
rect 41580 23940 41636 23950
rect 41580 23846 41636 23884
rect 41804 23828 41860 30716
rect 41916 30100 41972 31388
rect 41916 30006 41972 30044
rect 42252 30994 42308 31006
rect 42252 30942 42254 30994
rect 42306 30942 42308 30994
rect 42252 30212 42308 30942
rect 42588 30772 42644 32508
rect 42700 32498 42756 32508
rect 43036 32116 43092 32956
rect 43148 32452 43204 32462
rect 43204 32396 43316 32452
rect 43148 32386 43204 32396
rect 43148 32116 43204 32126
rect 43036 32060 43148 32116
rect 43148 32050 43204 32060
rect 41916 29426 41972 29438
rect 41916 29374 41918 29426
rect 41970 29374 41972 29426
rect 41916 28308 41972 29374
rect 42028 29204 42084 29214
rect 42028 29110 42084 29148
rect 41916 25060 41972 28252
rect 42028 28532 42084 28542
rect 42028 27858 42084 28476
rect 42252 28196 42308 30156
rect 42364 30716 42644 30772
rect 43260 30884 43316 32396
rect 42364 29650 42420 30716
rect 43036 30436 43092 30446
rect 43036 30212 43092 30380
rect 43260 30434 43316 30828
rect 43260 30382 43262 30434
rect 43314 30382 43316 30434
rect 43260 30370 43316 30382
rect 43372 30212 43428 35084
rect 43708 35026 43764 35038
rect 43708 34974 43710 35026
rect 43762 34974 43764 35026
rect 43596 34914 43652 34926
rect 43596 34862 43598 34914
rect 43650 34862 43652 34914
rect 43596 34692 43652 34862
rect 43596 34626 43652 34636
rect 43484 34580 43540 34590
rect 43484 34356 43540 34524
rect 43596 34356 43652 34366
rect 43484 34354 43652 34356
rect 43484 34302 43598 34354
rect 43650 34302 43652 34354
rect 43484 34300 43652 34302
rect 43596 34290 43652 34300
rect 43484 34132 43540 34142
rect 43484 32788 43540 34076
rect 43708 34020 43764 34974
rect 43708 33954 43764 33964
rect 43932 32900 43988 35868
rect 44044 33124 44100 40796
rect 44268 40628 44324 40638
rect 45052 40628 45108 42476
rect 45164 42196 45220 42206
rect 45276 42196 45332 42702
rect 45164 42194 45332 42196
rect 45164 42142 45166 42194
rect 45218 42142 45332 42194
rect 45164 42140 45332 42142
rect 45164 42130 45220 42140
rect 45388 41970 45444 41982
rect 45388 41918 45390 41970
rect 45442 41918 45444 41970
rect 45388 41074 45444 41918
rect 45388 41022 45390 41074
rect 45442 41022 45444 41074
rect 45164 40628 45220 40638
rect 45052 40572 45164 40628
rect 44268 40534 44324 40572
rect 45164 40562 45220 40572
rect 45388 40626 45444 41022
rect 45388 40574 45390 40626
rect 45442 40574 45444 40626
rect 45388 40562 45444 40574
rect 45500 40292 45556 46956
rect 45724 46898 45780 47404
rect 45836 47458 45892 48860
rect 46060 48804 46116 49308
rect 46284 49028 46340 51886
rect 46396 50932 46452 50942
rect 46396 50706 46452 50876
rect 46396 50654 46398 50706
rect 46450 50654 46452 50706
rect 46396 50642 46452 50654
rect 46620 49476 46676 54124
rect 46844 53620 46900 54238
rect 46956 53844 47012 54462
rect 46956 53778 47012 53788
rect 47516 54402 47572 54414
rect 47516 54350 47518 54402
rect 47570 54350 47572 54402
rect 47516 53732 47572 54350
rect 47516 53666 47572 53676
rect 46844 53554 46900 53564
rect 47516 53508 47572 53518
rect 46732 53060 46788 53070
rect 46732 52966 46788 53004
rect 47516 52946 47572 53452
rect 47628 53172 47684 54574
rect 47740 53732 47796 54796
rect 47964 54628 48020 55244
rect 48412 55186 48468 57932
rect 49196 57874 49252 58156
rect 49196 57822 49198 57874
rect 49250 57822 49252 57874
rect 49196 57810 49252 57822
rect 49420 58212 49476 58222
rect 49868 58212 49924 58222
rect 49420 58210 49924 58212
rect 49420 58158 49422 58210
rect 49474 58158 49870 58210
rect 49922 58158 49924 58210
rect 49420 58156 49924 58158
rect 48860 57652 48916 57662
rect 48860 56306 48916 57596
rect 48860 56254 48862 56306
rect 48914 56254 48916 56306
rect 48860 56242 48916 56254
rect 48972 56642 49028 56654
rect 48972 56590 48974 56642
rect 49026 56590 49028 56642
rect 48972 56084 49028 56590
rect 48412 55134 48414 55186
rect 48466 55134 48468 55186
rect 48412 55122 48468 55134
rect 48636 55748 48692 55758
rect 47964 54572 48356 54628
rect 48188 54402 48244 54414
rect 48188 54350 48190 54402
rect 48242 54350 48244 54402
rect 48076 54290 48132 54302
rect 48076 54238 48078 54290
rect 48130 54238 48132 54290
rect 47740 53284 47796 53676
rect 47740 53218 47796 53228
rect 47852 54068 47908 54078
rect 47628 53106 47684 53116
rect 47516 52894 47518 52946
rect 47570 52894 47572 52946
rect 47516 52882 47572 52894
rect 47740 52948 47796 52958
rect 47740 52854 47796 52892
rect 47852 52834 47908 54012
rect 47852 52782 47854 52834
rect 47906 52782 47908 52834
rect 47852 52770 47908 52782
rect 47964 53058 48020 53070
rect 47964 53006 47966 53058
rect 48018 53006 48020 53058
rect 47964 52836 48020 53006
rect 48076 53060 48132 54238
rect 48188 53844 48244 54350
rect 48188 53778 48244 53788
rect 48300 53506 48356 54572
rect 48300 53454 48302 53506
rect 48354 53454 48356 53506
rect 48300 53172 48356 53454
rect 48300 53106 48356 53116
rect 48076 52994 48132 53004
rect 47292 52500 47348 52510
rect 47292 52276 47348 52444
rect 47180 52274 47348 52276
rect 47180 52222 47294 52274
rect 47346 52222 47348 52274
rect 47180 52220 47348 52222
rect 46732 52162 46788 52174
rect 46732 52110 46734 52162
rect 46786 52110 46788 52162
rect 46732 52052 46788 52110
rect 46732 51986 46788 51996
rect 47180 50594 47236 52220
rect 47292 52210 47348 52220
rect 47740 51938 47796 51950
rect 47740 51886 47742 51938
rect 47794 51886 47796 51938
rect 47740 51604 47796 51886
rect 47180 50542 47182 50594
rect 47234 50542 47236 50594
rect 46620 49410 46676 49420
rect 46956 49812 47012 49822
rect 46956 49028 47012 49756
rect 47068 49700 47124 49710
rect 47068 49138 47124 49644
rect 47180 49252 47236 50542
rect 47180 49186 47236 49196
rect 47292 51602 47796 51604
rect 47292 51550 47742 51602
rect 47794 51550 47796 51602
rect 47292 51548 47796 51550
rect 47292 50372 47348 51548
rect 47740 51538 47796 51548
rect 47964 51044 48020 52780
rect 48188 52946 48244 52958
rect 48188 52894 48190 52946
rect 48242 52894 48244 52946
rect 48188 52724 48244 52894
rect 48636 52948 48692 55692
rect 48748 55298 48804 55310
rect 48748 55246 48750 55298
rect 48802 55246 48804 55298
rect 48748 54738 48804 55246
rect 48972 55076 49028 56028
rect 48748 54686 48750 54738
rect 48802 54686 48804 54738
rect 48748 54674 48804 54686
rect 48860 55020 49028 55076
rect 49084 56308 49140 56318
rect 48860 54292 48916 55020
rect 48860 54226 48916 54236
rect 48972 54852 49028 54862
rect 48860 53732 48916 53742
rect 48972 53732 49028 54796
rect 49084 54516 49140 56252
rect 49196 55858 49252 55870
rect 49196 55806 49198 55858
rect 49250 55806 49252 55858
rect 49196 55188 49252 55806
rect 49420 55748 49476 58156
rect 49868 58146 49924 58156
rect 50204 58210 50260 58222
rect 50204 58158 50206 58210
rect 50258 58158 50260 58210
rect 49756 57762 49812 57774
rect 49756 57710 49758 57762
rect 49810 57710 49812 57762
rect 49756 56308 49812 57710
rect 49980 57650 50036 57662
rect 49980 57598 49982 57650
rect 50034 57598 50036 57650
rect 49980 56308 50036 57598
rect 50092 56642 50148 56654
rect 50092 56590 50094 56642
rect 50146 56590 50148 56642
rect 50092 56532 50148 56590
rect 50092 56466 50148 56476
rect 50092 56308 50148 56318
rect 49980 56252 50092 56308
rect 49756 56242 49812 56252
rect 50092 56242 50148 56252
rect 49868 56194 49924 56206
rect 49868 56142 49870 56194
rect 49922 56142 49924 56194
rect 49756 56084 49812 56094
rect 49756 55990 49812 56028
rect 49420 55682 49476 55692
rect 49196 54628 49252 55132
rect 49308 55298 49364 55310
rect 49308 55246 49310 55298
rect 49362 55246 49364 55298
rect 49308 54852 49364 55246
rect 49868 55300 49924 56142
rect 50204 55300 50260 58158
rect 51324 58212 51380 58222
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50652 57540 50708 57550
rect 50652 57538 50932 57540
rect 50652 57486 50654 57538
rect 50706 57486 50932 57538
rect 50652 57484 50932 57486
rect 50652 57474 50708 57484
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 49868 55234 49924 55244
rect 49980 55244 50260 55300
rect 50316 56308 50372 56318
rect 50316 55298 50372 56252
rect 50540 56082 50596 56094
rect 50540 56030 50542 56082
rect 50594 56030 50596 56082
rect 50316 55246 50318 55298
rect 50370 55246 50372 55298
rect 49308 54786 49364 54796
rect 49868 54628 49924 54638
rect 49196 54626 49924 54628
rect 49196 54574 49870 54626
rect 49922 54574 49924 54626
rect 49196 54572 49924 54574
rect 49868 54562 49924 54572
rect 49980 54628 50036 55244
rect 49084 54460 49252 54516
rect 49084 54292 49140 54302
rect 49084 54198 49140 54236
rect 48860 53730 49028 53732
rect 48860 53678 48862 53730
rect 48914 53678 49028 53730
rect 48860 53676 49028 53678
rect 49084 53732 49140 53742
rect 49196 53732 49252 54460
rect 49308 54404 49364 54414
rect 49308 54402 49476 54404
rect 49308 54350 49310 54402
rect 49362 54350 49476 54402
rect 49308 54348 49476 54350
rect 49308 54338 49364 54348
rect 49084 53730 49252 53732
rect 49084 53678 49086 53730
rect 49138 53678 49252 53730
rect 49084 53676 49252 53678
rect 49308 54180 49364 54190
rect 48636 52892 48804 52948
rect 48188 52658 48244 52668
rect 48300 52276 48356 52286
rect 48076 52164 48132 52174
rect 48076 52050 48132 52108
rect 48300 52162 48356 52220
rect 48300 52110 48302 52162
rect 48354 52110 48356 52162
rect 48300 52098 48356 52110
rect 48076 51998 48078 52050
rect 48130 51998 48132 52050
rect 48076 51986 48132 51998
rect 47964 50978 48020 50988
rect 48636 50932 48692 50942
rect 47628 50818 47684 50830
rect 47628 50766 47630 50818
rect 47682 50766 47684 50818
rect 47516 50706 47572 50718
rect 47516 50654 47518 50706
rect 47570 50654 47572 50706
rect 47068 49086 47070 49138
rect 47122 49086 47124 49138
rect 47068 49074 47124 49086
rect 46284 48962 46340 48972
rect 46396 49026 47012 49028
rect 46396 48974 46958 49026
rect 47010 48974 47012 49026
rect 46396 48972 47012 48974
rect 46060 47682 46116 48748
rect 46284 48020 46340 48030
rect 46284 47926 46340 47964
rect 46060 47630 46062 47682
rect 46114 47630 46116 47682
rect 46060 47618 46116 47630
rect 45836 47406 45838 47458
rect 45890 47406 45892 47458
rect 45836 47348 45892 47406
rect 45836 47282 45892 47292
rect 46172 47346 46228 47358
rect 46172 47294 46174 47346
rect 46226 47294 46228 47346
rect 45724 46846 45726 46898
rect 45778 46846 45780 46898
rect 45724 46834 45780 46846
rect 45836 47124 45892 47134
rect 45836 46898 45892 47068
rect 45836 46846 45838 46898
rect 45890 46846 45892 46898
rect 45836 46834 45892 46846
rect 45948 47012 46004 47022
rect 45948 46898 46004 46956
rect 45948 46846 45950 46898
rect 46002 46846 46004 46898
rect 45948 46834 46004 46846
rect 45612 46788 45668 46826
rect 45612 46722 45668 46732
rect 46060 46788 46116 46798
rect 46172 46788 46228 47294
rect 46396 46898 46452 48972
rect 46956 48962 47012 48972
rect 47180 49028 47236 49038
rect 47180 48934 47236 48972
rect 47068 48916 47124 48926
rect 46396 46846 46398 46898
rect 46450 46846 46452 46898
rect 46396 46834 46452 46846
rect 46620 48244 46676 48254
rect 46116 46732 46228 46788
rect 45724 46564 45780 46574
rect 45724 45330 45780 46508
rect 46060 46114 46116 46732
rect 46060 46062 46062 46114
rect 46114 46062 46116 46114
rect 46060 46050 46116 46062
rect 46620 45780 46676 48188
rect 47068 48242 47124 48860
rect 47068 48190 47070 48242
rect 47122 48190 47124 48242
rect 46732 48132 46788 48142
rect 46732 46674 46788 48076
rect 46732 46622 46734 46674
rect 46786 46622 46788 46674
rect 46732 46610 46788 46622
rect 46844 47460 46900 47470
rect 45724 45278 45726 45330
rect 45778 45278 45780 45330
rect 45724 45266 45780 45278
rect 46396 45778 46676 45780
rect 46396 45726 46622 45778
rect 46674 45726 46676 45778
rect 46396 45724 46676 45726
rect 46060 44772 46116 44782
rect 46060 42978 46116 44716
rect 46172 44436 46228 44446
rect 46172 44342 46228 44380
rect 46060 42926 46062 42978
rect 46114 42926 46116 42978
rect 46060 42914 46116 42926
rect 45724 42754 45780 42766
rect 45724 42702 45726 42754
rect 45778 42702 45780 42754
rect 45724 42084 45780 42702
rect 46396 42194 46452 45724
rect 46620 45714 46676 45724
rect 46732 46116 46788 46126
rect 46732 45332 46788 46060
rect 46844 45890 46900 47404
rect 46844 45838 46846 45890
rect 46898 45838 46900 45890
rect 46844 45826 46900 45838
rect 46956 45892 47012 45902
rect 46844 45332 46900 45342
rect 46620 45330 46900 45332
rect 46620 45278 46846 45330
rect 46898 45278 46900 45330
rect 46620 45276 46900 45278
rect 46508 42532 46564 42542
rect 46508 42438 46564 42476
rect 46396 42142 46398 42194
rect 46450 42142 46452 42194
rect 46396 42130 46452 42142
rect 46060 42084 46116 42094
rect 45724 42018 45780 42028
rect 45836 42028 46060 42084
rect 45836 41970 45892 42028
rect 46060 42018 46116 42028
rect 46620 41972 46676 45276
rect 46844 45266 46900 45276
rect 46956 44322 47012 45836
rect 47068 45780 47124 48190
rect 47292 46674 47348 50316
rect 47404 50484 47460 50494
rect 47404 49810 47460 50428
rect 47404 49758 47406 49810
rect 47458 49758 47460 49810
rect 47404 49746 47460 49758
rect 47516 49700 47572 50654
rect 47516 49634 47572 49644
rect 47628 49028 47684 50766
rect 48076 50594 48132 50606
rect 48076 50542 48078 50594
rect 48130 50542 48132 50594
rect 47740 49812 47796 49822
rect 47740 49718 47796 49756
rect 47964 49364 48020 49374
rect 47516 48972 47684 49028
rect 47740 49252 47796 49262
rect 47516 47796 47572 48972
rect 47740 48916 47796 49196
rect 47740 48822 47796 48860
rect 47628 48804 47684 48814
rect 47628 48242 47684 48748
rect 47964 48802 48020 49308
rect 48076 49250 48132 50542
rect 48524 50594 48580 50606
rect 48524 50542 48526 50594
rect 48578 50542 48580 50594
rect 48412 50482 48468 50494
rect 48412 50430 48414 50482
rect 48466 50430 48468 50482
rect 48412 50428 48468 50430
rect 48076 49198 48078 49250
rect 48130 49198 48132 49250
rect 48076 49186 48132 49198
rect 48300 50372 48468 50428
rect 48524 50372 48580 50542
rect 47964 48750 47966 48802
rect 48018 48750 48020 48802
rect 47628 48190 47630 48242
rect 47682 48190 47684 48242
rect 47628 48178 47684 48190
rect 47740 48356 47796 48366
rect 47964 48356 48020 48750
rect 48188 48914 48244 48926
rect 48188 48862 48190 48914
rect 48242 48862 48244 48914
rect 48188 48804 48244 48862
rect 48188 48738 48244 48748
rect 47740 48354 48020 48356
rect 47740 48302 47742 48354
rect 47794 48302 48020 48354
rect 47740 48300 48020 48302
rect 47740 48020 47796 48300
rect 48076 48132 48132 48142
rect 48076 48130 48244 48132
rect 48076 48078 48078 48130
rect 48130 48078 48244 48130
rect 48076 48076 48244 48078
rect 48076 48066 48132 48076
rect 47740 47954 47796 47964
rect 47516 47730 47572 47740
rect 48076 47684 48132 47694
rect 47964 47628 48076 47684
rect 47516 47460 47572 47470
rect 47516 47366 47572 47404
rect 47516 47012 47572 47022
rect 47516 46786 47572 46956
rect 47516 46734 47518 46786
rect 47570 46734 47572 46786
rect 47516 46722 47572 46734
rect 47292 46622 47294 46674
rect 47346 46622 47348 46674
rect 47292 46610 47348 46622
rect 47068 45714 47124 45724
rect 47516 46004 47572 46014
rect 47180 45106 47236 45118
rect 47180 45054 47182 45106
rect 47234 45054 47236 45106
rect 47180 44996 47236 45054
rect 47404 44996 47460 45006
rect 47180 44930 47236 44940
rect 47292 44994 47460 44996
rect 47292 44942 47406 44994
rect 47458 44942 47460 44994
rect 47292 44940 47460 44942
rect 47516 44996 47572 45948
rect 47964 46002 48020 47628
rect 48076 47618 48132 47628
rect 48188 47012 48244 48076
rect 48300 47460 48356 50372
rect 48524 50306 48580 50316
rect 48636 49252 48692 50876
rect 48524 49196 48692 49252
rect 48524 47796 48580 49196
rect 48748 49140 48804 52892
rect 48860 52162 48916 53676
rect 48972 53506 49028 53518
rect 48972 53454 48974 53506
rect 49026 53454 49028 53506
rect 48972 53284 49028 53454
rect 49084 53508 49140 53676
rect 49308 53620 49364 54124
rect 49084 53442 49140 53452
rect 49196 53564 49364 53620
rect 48972 53218 49028 53228
rect 49196 52946 49252 53564
rect 49420 53172 49476 54348
rect 49980 54180 50036 54572
rect 49644 54124 50036 54180
rect 50092 55076 50148 55086
rect 49532 53730 49588 53742
rect 49532 53678 49534 53730
rect 49586 53678 49588 53730
rect 49532 53508 49588 53678
rect 49532 53442 49588 53452
rect 49420 53106 49476 53116
rect 49196 52894 49198 52946
rect 49250 52894 49252 52946
rect 49196 52882 49252 52894
rect 49308 52948 49364 52958
rect 49420 52948 49476 52958
rect 49364 52946 49476 52948
rect 49364 52894 49422 52946
rect 49474 52894 49476 52946
rect 49364 52892 49476 52894
rect 48860 52110 48862 52162
rect 48914 52110 48916 52162
rect 48860 52098 48916 52110
rect 49196 52612 49252 52622
rect 49196 51380 49252 52556
rect 49196 51286 49252 51324
rect 48972 51268 49028 51278
rect 48972 51174 49028 51212
rect 49196 50594 49252 50606
rect 49196 50542 49198 50594
rect 49250 50542 49252 50594
rect 49196 50372 49252 50542
rect 49196 50306 49252 50316
rect 48860 49922 48916 49934
rect 48860 49870 48862 49922
rect 48914 49870 48916 49922
rect 48860 49364 48916 49870
rect 49196 49810 49252 49822
rect 49196 49758 49198 49810
rect 49250 49758 49252 49810
rect 48860 49298 48916 49308
rect 48972 49700 49028 49710
rect 48748 49084 48916 49140
rect 48748 48916 48804 48926
rect 48748 48822 48804 48860
rect 48748 48468 48804 48478
rect 48748 48132 48804 48412
rect 48860 48356 48916 49084
rect 48972 49026 49028 49644
rect 48972 48974 48974 49026
rect 49026 48974 49028 49026
rect 48972 48962 49028 48974
rect 49196 48804 49252 49758
rect 49308 49364 49364 52892
rect 49420 52882 49476 52892
rect 49532 51380 49588 51390
rect 49420 50820 49476 50830
rect 49420 50726 49476 50764
rect 49532 49588 49588 51324
rect 49644 50428 49700 54124
rect 49756 53732 49812 53742
rect 49756 53638 49812 53676
rect 50092 53618 50148 55020
rect 50092 53566 50094 53618
rect 50146 53566 50148 53618
rect 49980 53396 50036 53406
rect 49980 53058 50036 53340
rect 49980 53006 49982 53058
rect 50034 53006 50036 53058
rect 49980 52994 50036 53006
rect 49868 52946 49924 52958
rect 49868 52894 49870 52946
rect 49922 52894 49924 52946
rect 49868 52836 49924 52894
rect 49868 52770 49924 52780
rect 50092 52612 50148 53566
rect 50092 52546 50148 52556
rect 50204 52834 50260 52846
rect 50204 52782 50206 52834
rect 50258 52782 50260 52834
rect 50204 52724 50260 52782
rect 50092 52386 50148 52398
rect 50092 52334 50094 52386
rect 50146 52334 50148 52386
rect 49980 52164 50036 52174
rect 49980 52070 50036 52108
rect 49980 51266 50036 51278
rect 49980 51214 49982 51266
rect 50034 51214 50036 51266
rect 49756 50708 49812 50746
rect 49756 50642 49812 50652
rect 49980 50708 50036 51214
rect 49980 50642 50036 50652
rect 49756 50482 49812 50494
rect 49756 50430 49758 50482
rect 49810 50430 49812 50482
rect 49756 50428 49812 50430
rect 49644 50372 49812 50428
rect 49980 50484 50036 50522
rect 49980 50418 50036 50428
rect 49644 50260 49700 50270
rect 49644 49810 49700 50204
rect 49980 50260 50036 50270
rect 49756 50034 49812 50046
rect 49756 49982 49758 50034
rect 49810 49982 49812 50034
rect 49756 49924 49812 49982
rect 49756 49858 49812 49868
rect 49644 49758 49646 49810
rect 49698 49758 49700 49810
rect 49644 49746 49700 49758
rect 49532 49532 49812 49588
rect 49308 49308 49476 49364
rect 49308 49140 49364 49150
rect 49308 49046 49364 49084
rect 49196 48738 49252 48748
rect 49196 48580 49252 48590
rect 48860 48300 49028 48356
rect 48860 48132 48916 48142
rect 48748 48130 48916 48132
rect 48748 48078 48862 48130
rect 48914 48078 48916 48130
rect 48748 48076 48916 48078
rect 48860 48066 48916 48076
rect 48524 47740 48692 47796
rect 48300 47394 48356 47404
rect 48636 47460 48692 47740
rect 48860 47460 48916 47470
rect 48636 47458 48916 47460
rect 48636 47406 48862 47458
rect 48914 47406 48916 47458
rect 48636 47404 48916 47406
rect 48636 47012 48692 47404
rect 48860 47394 48916 47404
rect 48188 46956 48468 47012
rect 48076 46786 48132 46798
rect 48076 46734 48078 46786
rect 48130 46734 48132 46786
rect 48076 46676 48132 46734
rect 48188 46788 48244 46798
rect 48188 46694 48244 46732
rect 48076 46610 48132 46620
rect 47964 45950 47966 46002
rect 48018 45950 48020 46002
rect 47852 45892 47908 45902
rect 47852 45798 47908 45836
rect 47628 45220 47684 45230
rect 47628 45126 47684 45164
rect 47740 45108 47796 45118
rect 47740 45014 47796 45052
rect 47516 44940 47684 44996
rect 46956 44270 46958 44322
rect 47010 44270 47012 44322
rect 46956 44258 47012 44270
rect 46732 43652 46788 43662
rect 47292 43652 47348 44940
rect 47404 44930 47460 44940
rect 47404 44772 47460 44782
rect 47404 44322 47460 44716
rect 47628 44660 47684 44940
rect 47964 44772 48020 45950
rect 47964 44706 48020 44716
rect 48076 46450 48132 46462
rect 48076 46398 48078 46450
rect 48130 46398 48132 46450
rect 47628 44604 47796 44660
rect 47404 44270 47406 44322
rect 47458 44270 47460 44322
rect 47404 44258 47460 44270
rect 46732 42754 46788 43596
rect 47068 43596 47348 43652
rect 46956 43428 47012 43438
rect 46732 42702 46734 42754
rect 46786 42702 46788 42754
rect 46732 42690 46788 42702
rect 46844 43372 46956 43428
rect 46844 42084 46900 43372
rect 46956 43362 47012 43372
rect 47068 42196 47124 43596
rect 47516 43540 47572 43550
rect 47292 43538 47572 43540
rect 47292 43486 47518 43538
rect 47570 43486 47572 43538
rect 47292 43484 47572 43486
rect 47180 43428 47236 43438
rect 47180 43334 47236 43372
rect 47068 42130 47124 42140
rect 45836 41918 45838 41970
rect 45890 41918 45892 41970
rect 45836 41906 45892 41918
rect 46172 41916 46676 41972
rect 46732 41972 46788 41982
rect 46844 41972 46900 42028
rect 47292 41972 47348 43484
rect 47516 43474 47572 43484
rect 46732 41970 46900 41972
rect 46732 41918 46734 41970
rect 46786 41918 46900 41970
rect 46732 41916 46900 41918
rect 47180 41916 47348 41972
rect 46060 41860 46116 41870
rect 46172 41860 46228 41916
rect 46732 41906 46788 41916
rect 46060 41858 46228 41860
rect 46060 41806 46062 41858
rect 46114 41806 46228 41858
rect 46060 41804 46228 41806
rect 46060 41794 46116 41804
rect 46508 41748 46564 41758
rect 45500 40226 45556 40236
rect 45724 41186 45780 41198
rect 45724 41134 45726 41186
rect 45778 41134 45780 41186
rect 45724 40628 45780 41134
rect 46060 40964 46116 40974
rect 46060 40870 46116 40908
rect 44268 40068 44324 40078
rect 44268 39730 44324 40012
rect 44940 40068 44996 40078
rect 44940 39842 44996 40012
rect 44940 39790 44942 39842
rect 44994 39790 44996 39842
rect 44940 39778 44996 39790
rect 44268 39678 44270 39730
rect 44322 39678 44324 39730
rect 44268 39666 44324 39678
rect 45724 39508 45780 40572
rect 46060 40404 46116 40414
rect 46060 40290 46116 40348
rect 46060 40238 46062 40290
rect 46114 40238 46116 40290
rect 46060 40226 46116 40238
rect 46284 39508 46340 39518
rect 45724 39506 46340 39508
rect 45724 39454 46286 39506
rect 46338 39454 46340 39506
rect 45724 39452 46340 39454
rect 46284 39442 46340 39452
rect 46508 39060 46564 41692
rect 46956 41746 47012 41758
rect 46956 41694 46958 41746
rect 47010 41694 47012 41746
rect 46956 40852 47012 41694
rect 46732 40796 47012 40852
rect 47180 41186 47236 41916
rect 47628 41860 47684 41870
rect 47628 41766 47684 41804
rect 47292 41746 47348 41758
rect 47292 41694 47294 41746
rect 47346 41694 47348 41746
rect 47292 41636 47348 41694
rect 47292 41580 47572 41636
rect 47180 41134 47182 41186
rect 47234 41134 47236 41186
rect 46732 40068 46788 40796
rect 47068 40740 47124 40750
rect 46844 40684 47068 40740
rect 46844 40402 46900 40684
rect 47068 40674 47124 40684
rect 46844 40350 46846 40402
rect 46898 40350 46900 40402
rect 46844 40338 46900 40350
rect 46844 40068 46900 40078
rect 46732 40012 46844 40068
rect 46844 40002 46900 40012
rect 47180 39172 47236 41134
rect 47292 40964 47348 40974
rect 47292 40402 47348 40908
rect 47292 40350 47294 40402
rect 47346 40350 47348 40402
rect 47292 39508 47348 40350
rect 47404 40740 47460 40750
rect 47404 39732 47460 40684
rect 47516 40404 47572 41580
rect 47740 41188 47796 44604
rect 48076 44324 48132 46398
rect 48300 45668 48356 45678
rect 48076 44258 48132 44268
rect 48188 45220 48244 45230
rect 47964 44100 48020 44110
rect 47852 43652 47908 43662
rect 47852 42754 47908 43596
rect 47964 43650 48020 44044
rect 48188 43764 48244 45164
rect 48300 44322 48356 45612
rect 48300 44270 48302 44322
rect 48354 44270 48356 44322
rect 48300 44258 48356 44270
rect 48188 43698 48244 43708
rect 47964 43598 47966 43650
rect 48018 43598 48020 43650
rect 47964 43586 48020 43598
rect 48188 43538 48244 43550
rect 48188 43486 48190 43538
rect 48242 43486 48244 43538
rect 47852 42702 47854 42754
rect 47906 42702 47908 42754
rect 47852 42690 47908 42702
rect 48076 43426 48132 43438
rect 48076 43374 48078 43426
rect 48130 43374 48132 43426
rect 47852 41972 47908 41982
rect 47852 41878 47908 41916
rect 47740 41122 47796 41132
rect 47852 40852 47908 40862
rect 47628 40404 47684 40414
rect 47516 40402 47684 40404
rect 47516 40350 47630 40402
rect 47682 40350 47684 40402
rect 47516 40348 47684 40350
rect 47628 40338 47684 40348
rect 47404 39620 47460 39676
rect 47516 39620 47572 39630
rect 47404 39618 47572 39620
rect 47404 39566 47518 39618
rect 47570 39566 47572 39618
rect 47404 39564 47572 39566
rect 47516 39554 47572 39564
rect 47292 39414 47348 39452
rect 47404 39396 47460 39406
rect 47404 39302 47460 39340
rect 47516 39284 47572 39294
rect 47180 39116 47460 39172
rect 46508 38966 46564 39004
rect 45500 38946 45556 38958
rect 45500 38894 45502 38946
rect 45554 38894 45556 38946
rect 45052 38836 45108 38846
rect 45052 38722 45108 38780
rect 45052 38670 45054 38722
rect 45106 38670 45108 38722
rect 45052 38658 45108 38670
rect 44940 38164 44996 38174
rect 44156 37938 44212 37950
rect 44156 37886 44158 37938
rect 44210 37886 44212 37938
rect 44156 37828 44212 37886
rect 44716 37940 44772 37950
rect 44156 37772 44660 37828
rect 44268 37492 44324 37502
rect 44268 37266 44324 37436
rect 44268 37214 44270 37266
rect 44322 37214 44324 37266
rect 44268 37202 44324 37214
rect 44380 37154 44436 37166
rect 44380 37102 44382 37154
rect 44434 37102 44436 37154
rect 44380 36036 44436 37102
rect 44380 35970 44436 35980
rect 44268 35810 44324 35822
rect 44268 35758 44270 35810
rect 44322 35758 44324 35810
rect 44268 35700 44324 35758
rect 44268 35364 44324 35644
rect 44268 35298 44324 35308
rect 44492 35698 44548 35710
rect 44492 35646 44494 35698
rect 44546 35646 44548 35698
rect 44156 34132 44212 34142
rect 44156 34038 44212 34076
rect 44492 34132 44548 35646
rect 44604 35140 44660 37772
rect 44716 35476 44772 37884
rect 44940 37268 44996 38108
rect 45500 38164 45556 38894
rect 45836 38836 45892 38846
rect 45836 38742 45892 38780
rect 46060 38834 46116 38846
rect 46060 38782 46062 38834
rect 46114 38782 46116 38834
rect 45500 38108 45892 38164
rect 45276 38052 45332 38062
rect 44940 37202 44996 37212
rect 45164 38050 45332 38052
rect 45164 37998 45278 38050
rect 45330 37998 45332 38050
rect 45164 37996 45332 37998
rect 44828 36484 44884 36494
rect 45052 36484 45108 36494
rect 44828 36390 44884 36428
rect 44940 36482 45108 36484
rect 44940 36430 45054 36482
rect 45106 36430 45108 36482
rect 44940 36428 45108 36430
rect 44940 35700 44996 36428
rect 45052 36418 45108 36428
rect 45164 35924 45220 37996
rect 45276 37986 45332 37996
rect 45164 35858 45220 35868
rect 45276 36596 45332 36606
rect 45052 35812 45108 35822
rect 45052 35718 45108 35756
rect 44940 35634 44996 35644
rect 45164 35588 45220 35598
rect 44716 35420 44996 35476
rect 44828 35140 44884 35150
rect 44604 35138 44884 35140
rect 44604 35086 44830 35138
rect 44882 35086 44884 35138
rect 44604 35084 44884 35086
rect 44828 35074 44884 35084
rect 44940 35138 44996 35420
rect 44940 35086 44942 35138
rect 44994 35086 44996 35138
rect 44492 34066 44548 34076
rect 44940 33908 44996 35086
rect 45164 35138 45220 35532
rect 45164 35086 45166 35138
rect 45218 35086 45220 35138
rect 45164 35074 45220 35086
rect 45276 35138 45332 36540
rect 45388 36258 45444 36270
rect 45388 36206 45390 36258
rect 45442 36206 45444 36258
rect 45388 35698 45444 36206
rect 45388 35646 45390 35698
rect 45442 35646 45444 35698
rect 45388 35634 45444 35646
rect 45276 35086 45278 35138
rect 45330 35086 45332 35138
rect 45276 35074 45332 35086
rect 45388 34244 45444 34254
rect 45500 34244 45556 38108
rect 45724 37938 45780 37950
rect 45724 37886 45726 37938
rect 45778 37886 45780 37938
rect 45724 37828 45780 37886
rect 45836 37938 45892 38108
rect 46060 38050 46116 38782
rect 46732 38834 46788 38846
rect 46732 38782 46734 38834
rect 46786 38782 46788 38834
rect 46620 38722 46676 38734
rect 46620 38670 46622 38722
rect 46674 38670 46676 38722
rect 46620 38668 46676 38670
rect 46508 38612 46676 38668
rect 46732 38612 46788 38782
rect 46396 38164 46452 38174
rect 46060 37998 46062 38050
rect 46114 37998 46116 38050
rect 46060 37986 46116 37998
rect 46172 38162 46452 38164
rect 46172 38110 46398 38162
rect 46450 38110 46452 38162
rect 46172 38108 46452 38110
rect 45836 37886 45838 37938
rect 45890 37886 45892 37938
rect 45836 37874 45892 37886
rect 45724 36820 45780 37772
rect 46172 37716 46228 38108
rect 46396 38098 46452 38108
rect 45948 37660 46228 37716
rect 46284 37938 46340 37950
rect 46284 37886 46286 37938
rect 46338 37886 46340 37938
rect 45836 37380 45892 37390
rect 45836 37286 45892 37324
rect 45724 36754 45780 36764
rect 45612 36484 45668 36494
rect 45668 36428 45780 36484
rect 45612 36418 45668 36428
rect 45612 35700 45668 35710
rect 45612 34692 45668 35644
rect 45612 34626 45668 34636
rect 45388 34242 45556 34244
rect 45388 34190 45390 34242
rect 45442 34190 45556 34242
rect 45388 34188 45556 34190
rect 45388 34178 45444 34188
rect 45724 34020 45780 36428
rect 45948 35588 46004 37660
rect 46284 37492 46340 37886
rect 46060 37436 46340 37492
rect 46060 36260 46116 37436
rect 46396 37378 46452 37390
rect 46396 37326 46398 37378
rect 46450 37326 46452 37378
rect 46172 37268 46228 37278
rect 46396 37268 46452 37326
rect 46228 37212 46340 37268
rect 46172 37202 46228 37212
rect 46172 36596 46228 36634
rect 46172 36530 46228 36540
rect 46284 36370 46340 37212
rect 46396 37202 46452 37212
rect 46284 36318 46286 36370
rect 46338 36318 46340 36370
rect 46284 36306 46340 36318
rect 46396 36482 46452 36494
rect 46396 36430 46398 36482
rect 46450 36430 46452 36482
rect 46060 36194 46116 36204
rect 46396 36260 46452 36430
rect 46396 36194 46452 36204
rect 45836 35532 46004 35588
rect 45836 35476 45892 35532
rect 46508 35476 46564 38612
rect 46732 38546 46788 38556
rect 46956 38836 47012 38846
rect 46732 38388 46788 38398
rect 46620 38164 46676 38174
rect 46620 38050 46676 38108
rect 46620 37998 46622 38050
rect 46674 37998 46676 38050
rect 46620 37986 46676 37998
rect 46732 37378 46788 38332
rect 46732 37326 46734 37378
rect 46786 37326 46788 37378
rect 46732 37314 46788 37326
rect 46844 37938 46900 37950
rect 46844 37886 46846 37938
rect 46898 37886 46900 37938
rect 46844 37492 46900 37886
rect 46620 37266 46676 37278
rect 46620 37214 46622 37266
rect 46674 37214 46676 37266
rect 46620 37044 46676 37214
rect 46620 36978 46676 36988
rect 46844 36594 46900 37436
rect 46844 36542 46846 36594
rect 46898 36542 46900 36594
rect 46844 36530 46900 36542
rect 45836 35410 45892 35420
rect 45948 35420 46564 35476
rect 46844 35812 46900 35822
rect 45836 34690 45892 34702
rect 45836 34638 45838 34690
rect 45890 34638 45892 34690
rect 45836 34356 45892 34638
rect 45836 34290 45892 34300
rect 45724 33954 45780 33964
rect 44940 33852 45108 33908
rect 44156 33348 44212 33358
rect 44156 33254 44212 33292
rect 45052 33346 45108 33852
rect 45836 33796 45892 33806
rect 45836 33460 45892 33740
rect 45724 33348 45780 33358
rect 45052 33294 45054 33346
rect 45106 33294 45108 33346
rect 44044 33058 44100 33068
rect 44268 33236 44324 33246
rect 43932 32844 44100 32900
rect 43596 32788 43652 32798
rect 43484 32786 43652 32788
rect 43484 32734 43598 32786
rect 43650 32734 43652 32786
rect 43484 32732 43652 32734
rect 43596 32722 43652 32732
rect 43932 32338 43988 32350
rect 43932 32286 43934 32338
rect 43986 32286 43988 32338
rect 43820 32228 43876 32238
rect 43596 31892 43652 31902
rect 43596 31798 43652 31836
rect 43708 31780 43764 31790
rect 43708 31218 43764 31724
rect 43708 31166 43710 31218
rect 43762 31166 43764 31218
rect 43708 31154 43764 31166
rect 42700 30210 43092 30212
rect 42700 30158 43038 30210
rect 43090 30158 43092 30210
rect 42700 30156 43092 30158
rect 42364 29598 42366 29650
rect 42418 29598 42420 29650
rect 42364 29586 42420 29598
rect 42476 29986 42532 29998
rect 42476 29934 42478 29986
rect 42530 29934 42532 29986
rect 42476 29540 42532 29934
rect 42476 29474 42532 29484
rect 42700 29426 42756 30156
rect 43036 30146 43092 30156
rect 43148 30156 43372 30212
rect 42700 29374 42702 29426
rect 42754 29374 42756 29426
rect 42700 29362 42756 29374
rect 42924 29428 42980 29438
rect 43148 29428 43204 30156
rect 43372 30146 43428 30156
rect 43820 30100 43876 32172
rect 43932 32116 43988 32286
rect 43932 32050 43988 32060
rect 43932 31892 43988 31902
rect 43932 30436 43988 31836
rect 43932 30342 43988 30380
rect 42924 29426 43204 29428
rect 42924 29374 42926 29426
rect 42978 29374 43204 29426
rect 42924 29372 43204 29374
rect 43372 29988 43428 29998
rect 42924 29362 42980 29372
rect 43260 29316 43316 29326
rect 43036 29314 43316 29316
rect 43036 29262 43262 29314
rect 43314 29262 43316 29314
rect 43036 29260 43316 29262
rect 42700 29092 42756 29102
rect 42700 28642 42756 29036
rect 42700 28590 42702 28642
rect 42754 28590 42756 28642
rect 42700 28532 42756 28590
rect 42700 28466 42756 28476
rect 42252 28140 42532 28196
rect 42028 27806 42030 27858
rect 42082 27806 42084 27858
rect 42028 27794 42084 27806
rect 42476 27860 42532 28140
rect 43036 27972 43092 29260
rect 43260 29250 43316 29260
rect 43148 28084 43204 28094
rect 43148 27990 43204 28028
rect 42924 27916 43092 27972
rect 42812 27860 42868 27870
rect 42476 27858 42868 27860
rect 42476 27806 42814 27858
rect 42866 27806 42868 27858
rect 42476 27804 42868 27806
rect 42812 27794 42868 27804
rect 42924 27636 42980 27916
rect 42588 27580 42980 27636
rect 42252 26292 42308 26302
rect 42252 26198 42308 26236
rect 42476 26290 42532 26302
rect 42476 26238 42478 26290
rect 42530 26238 42532 26290
rect 41916 24994 41972 25004
rect 41916 24834 41972 24846
rect 41916 24782 41918 24834
rect 41970 24782 41972 24834
rect 41916 23940 41972 24782
rect 41916 23884 42084 23940
rect 41804 23762 41860 23772
rect 41692 23716 41748 23726
rect 41692 23622 41748 23660
rect 41916 23714 41972 23726
rect 41916 23662 41918 23714
rect 41970 23662 41972 23714
rect 41580 23604 41636 23614
rect 41020 21534 41022 21586
rect 41074 21534 41076 21586
rect 41020 21522 41076 21534
rect 41132 21532 41300 21588
rect 41356 23044 41412 23054
rect 40908 20750 40910 20802
rect 40962 20750 40964 20802
rect 40908 20738 40964 20750
rect 40796 20638 40798 20690
rect 40850 20638 40852 20690
rect 40796 20626 40852 20638
rect 40684 20468 40740 20478
rect 40684 19796 40740 20412
rect 40684 19730 40740 19740
rect 41132 19572 41188 21532
rect 41244 21364 41300 21374
rect 41356 21364 41412 22988
rect 41580 22146 41636 23548
rect 41804 23492 41860 23502
rect 41692 23380 41748 23390
rect 41692 22370 41748 23324
rect 41804 23154 41860 23436
rect 41804 23102 41806 23154
rect 41858 23102 41860 23154
rect 41804 23090 41860 23102
rect 41692 22318 41694 22370
rect 41746 22318 41748 22370
rect 41692 22306 41748 22318
rect 41804 22596 41860 22606
rect 41580 22094 41582 22146
rect 41634 22094 41636 22146
rect 41580 22082 41636 22094
rect 41580 21812 41636 21822
rect 41804 21812 41860 22540
rect 41580 21810 41860 21812
rect 41580 21758 41582 21810
rect 41634 21758 41860 21810
rect 41580 21756 41860 21758
rect 41916 21810 41972 23662
rect 42028 23268 42084 23884
rect 42476 23604 42532 26238
rect 42588 25732 42644 27580
rect 43372 27412 43428 29932
rect 43596 29986 43652 29998
rect 43596 29934 43598 29986
rect 43650 29934 43652 29986
rect 43596 29316 43652 29934
rect 43820 29650 43876 30044
rect 43820 29598 43822 29650
rect 43874 29598 43876 29650
rect 43820 29586 43876 29598
rect 43596 29250 43652 29260
rect 43932 28756 43988 28766
rect 43932 28642 43988 28700
rect 43932 28590 43934 28642
rect 43986 28590 43988 28642
rect 43932 28578 43988 28590
rect 44044 28420 44100 32844
rect 44156 32676 44212 32686
rect 44268 32676 44324 33180
rect 45052 33236 45108 33294
rect 45612 33292 45724 33348
rect 45052 33170 45108 33180
rect 45164 33234 45220 33246
rect 45164 33182 45166 33234
rect 45218 33182 45220 33234
rect 44492 32676 44548 32686
rect 44156 32674 44548 32676
rect 44156 32622 44158 32674
rect 44210 32622 44494 32674
rect 44546 32622 44548 32674
rect 44156 32620 44548 32622
rect 44156 32610 44212 32620
rect 44492 32610 44548 32620
rect 44716 32562 44772 32574
rect 44716 32510 44718 32562
rect 44770 32510 44772 32562
rect 44716 31892 44772 32510
rect 44716 31826 44772 31836
rect 45164 31892 45220 33182
rect 45388 32564 45444 32574
rect 45388 32470 45444 32508
rect 45164 31826 45220 31836
rect 45276 31778 45332 31790
rect 45276 31726 45278 31778
rect 45330 31726 45332 31778
rect 44156 31668 44212 31678
rect 44156 31574 44212 31612
rect 45276 31556 45332 31726
rect 45276 31490 45332 31500
rect 44828 31220 44884 31230
rect 44828 31126 44884 31164
rect 45612 31106 45668 33292
rect 45724 33254 45780 33292
rect 45724 31892 45780 31902
rect 45836 31892 45892 33404
rect 45948 32676 46004 35420
rect 46284 34916 46340 34926
rect 46844 34916 46900 35756
rect 46172 34914 46900 34916
rect 46172 34862 46286 34914
rect 46338 34862 46900 34914
rect 46172 34860 46900 34862
rect 46060 33572 46116 33582
rect 46172 33572 46228 34860
rect 46284 34850 46340 34860
rect 46508 34692 46564 34702
rect 46508 34130 46564 34636
rect 46844 34356 46900 34366
rect 46844 34262 46900 34300
rect 46956 34244 47012 38780
rect 47180 38052 47236 38062
rect 47180 37958 47236 37996
rect 47292 37940 47348 37950
rect 47292 37846 47348 37884
rect 47404 37492 47460 39116
rect 47516 38946 47572 39228
rect 47852 39058 47908 40796
rect 47964 39620 48020 39630
rect 47964 39526 48020 39564
rect 47852 39006 47854 39058
rect 47906 39006 47908 39058
rect 47852 38994 47908 39006
rect 47964 39060 48020 39070
rect 47964 38966 48020 39004
rect 47516 38894 47518 38946
rect 47570 38894 47572 38946
rect 47516 38882 47572 38894
rect 47628 38948 47684 38958
rect 47628 38854 47684 38892
rect 47740 38946 47796 38958
rect 47740 38894 47742 38946
rect 47794 38894 47796 38946
rect 47740 38836 47796 38894
rect 47740 38770 47796 38780
rect 47516 38612 47572 38622
rect 47572 38556 47684 38612
rect 47516 38546 47572 38556
rect 47292 37436 47460 37492
rect 47516 37716 47572 37726
rect 47180 37154 47236 37166
rect 47180 37102 47182 37154
rect 47234 37102 47236 37154
rect 47180 36932 47236 37102
rect 47180 36866 47236 36876
rect 47180 36482 47236 36494
rect 47180 36430 47182 36482
rect 47234 36430 47236 36482
rect 47180 35700 47236 36430
rect 47180 35606 47236 35644
rect 46956 34178 47012 34188
rect 46508 34078 46510 34130
rect 46562 34078 46564 34130
rect 46508 34066 46564 34078
rect 47180 34132 47236 34142
rect 47180 34038 47236 34076
rect 46284 34020 46340 34030
rect 46284 33926 46340 33964
rect 46060 33570 46228 33572
rect 46060 33518 46062 33570
rect 46114 33518 46228 33570
rect 46060 33516 46228 33518
rect 47068 33572 47124 33582
rect 46060 33506 46116 33516
rect 46844 33236 46900 33246
rect 46844 33142 46900 33180
rect 46508 33124 46564 33134
rect 46172 33122 46564 33124
rect 46172 33070 46510 33122
rect 46562 33070 46564 33122
rect 46172 33068 46564 33070
rect 46060 32676 46116 32686
rect 45948 32674 46116 32676
rect 45948 32622 46062 32674
rect 46114 32622 46116 32674
rect 45948 32620 46116 32622
rect 46060 32610 46116 32620
rect 45724 31890 45892 31892
rect 45724 31838 45726 31890
rect 45778 31838 45892 31890
rect 45724 31836 45892 31838
rect 45724 31826 45780 31836
rect 46172 31780 46228 33068
rect 46508 33058 46564 33068
rect 46508 32004 46564 32014
rect 45612 31054 45614 31106
rect 45666 31054 45668 31106
rect 45612 31042 45668 31054
rect 45948 31724 46228 31780
rect 46284 31892 46340 31902
rect 45948 31220 46004 31724
rect 46284 31668 46340 31836
rect 46172 31612 46340 31668
rect 46060 31556 46116 31566
rect 46060 31462 46116 31500
rect 45948 31106 46004 31164
rect 45948 31054 45950 31106
rect 46002 31054 46004 31106
rect 45948 31042 46004 31054
rect 46172 30994 46228 31612
rect 46172 30942 46174 30994
rect 46226 30942 46228 30994
rect 46172 30930 46228 30942
rect 46284 31220 46340 31230
rect 46508 31220 46564 31948
rect 44380 30884 44436 30894
rect 44156 30212 44212 30222
rect 44156 30118 44212 30156
rect 43932 28364 44100 28420
rect 44156 29426 44212 29438
rect 44156 29374 44158 29426
rect 44210 29374 44212 29426
rect 44156 29204 44212 29374
rect 43932 27746 43988 28364
rect 43932 27694 43934 27746
rect 43986 27694 43988 27746
rect 43932 27682 43988 27694
rect 44044 27970 44100 27982
rect 44044 27918 44046 27970
rect 44098 27918 44100 27970
rect 42812 27356 43428 27412
rect 43820 27636 43876 27646
rect 42588 25666 42644 25676
rect 42700 27188 42756 27198
rect 42588 25508 42644 25518
rect 42588 25414 42644 25452
rect 42588 23828 42644 23838
rect 42700 23828 42756 27132
rect 42588 23826 42756 23828
rect 42588 23774 42590 23826
rect 42642 23774 42756 23826
rect 42588 23772 42756 23774
rect 42812 26964 42868 27356
rect 43148 27188 43204 27198
rect 43148 27094 43204 27132
rect 42588 23762 42644 23772
rect 42476 23538 42532 23548
rect 42028 22260 42084 23212
rect 42364 23156 42420 23166
rect 42364 23062 42420 23100
rect 42700 22260 42756 22270
rect 42028 22258 42756 22260
rect 42028 22206 42702 22258
rect 42754 22206 42756 22258
rect 42028 22204 42756 22206
rect 41916 21758 41918 21810
rect 41970 21758 41972 21810
rect 41580 21746 41636 21756
rect 41916 21746 41972 21758
rect 42140 21812 42196 21822
rect 42140 21718 42196 21756
rect 41244 21362 41412 21364
rect 41244 21310 41246 21362
rect 41298 21310 41412 21362
rect 41244 21308 41412 21310
rect 41468 21700 41524 21710
rect 41244 21298 41300 21308
rect 41356 20692 41412 20702
rect 40124 15810 40180 15820
rect 40348 16828 40516 16884
rect 40572 19516 41188 19572
rect 41244 20690 41412 20692
rect 41244 20638 41358 20690
rect 41410 20638 41412 20690
rect 41244 20636 41412 20638
rect 41244 19572 41300 20636
rect 41356 20626 41412 20636
rect 40012 15596 40292 15652
rect 39788 15484 40180 15540
rect 39788 15314 39844 15484
rect 39788 15262 39790 15314
rect 39842 15262 39844 15314
rect 39788 15250 39844 15262
rect 40012 15314 40068 15326
rect 40012 15262 40014 15314
rect 40066 15262 40068 15314
rect 39900 15202 39956 15214
rect 39900 15150 39902 15202
rect 39954 15150 39956 15202
rect 39900 15148 39956 15150
rect 39116 14700 39284 14756
rect 39340 15092 39956 15148
rect 39116 12740 39172 14700
rect 39228 14532 39284 14542
rect 39228 14438 39284 14476
rect 39340 13858 39396 15092
rect 39452 14980 39508 14990
rect 39508 14924 39844 14980
rect 39452 14914 39508 14924
rect 39452 14420 39508 14430
rect 39508 14364 39732 14420
rect 39452 14354 39508 14364
rect 39340 13806 39342 13858
rect 39394 13806 39396 13858
rect 39340 13794 39396 13806
rect 39564 14196 39620 14206
rect 39564 13858 39620 14140
rect 39564 13806 39566 13858
rect 39618 13806 39620 13858
rect 39564 13794 39620 13806
rect 39564 13524 39620 13534
rect 39228 13074 39284 13086
rect 39228 13022 39230 13074
rect 39282 13022 39284 13074
rect 39228 12964 39284 13022
rect 39228 12898 39284 12908
rect 39228 12740 39284 12750
rect 39116 12684 39228 12740
rect 39228 12674 39284 12684
rect 38668 11666 38724 11676
rect 38780 12460 39060 12516
rect 39116 12516 39172 12526
rect 38780 9826 38836 12460
rect 39116 12292 39172 12460
rect 39116 12290 39508 12292
rect 39116 12238 39118 12290
rect 39170 12238 39508 12290
rect 39116 12236 39508 12238
rect 38892 12180 38948 12190
rect 38892 12086 38948 12124
rect 38780 9774 38782 9826
rect 38834 9774 38836 9826
rect 38780 9762 38836 9774
rect 39116 9714 39172 12236
rect 39452 11282 39508 12236
rect 39452 11230 39454 11282
rect 39506 11230 39508 11282
rect 39452 11218 39508 11230
rect 39116 9662 39118 9714
rect 39170 9662 39172 9714
rect 39116 9650 39172 9662
rect 39228 10498 39284 10510
rect 39228 10446 39230 10498
rect 39282 10446 39284 10498
rect 38444 9548 38612 9604
rect 38668 9604 38724 9614
rect 38444 8820 38500 9548
rect 38668 9156 38724 9548
rect 38892 9380 38948 9390
rect 38556 9100 38724 9156
rect 38780 9156 38836 9166
rect 38556 9044 38612 9100
rect 38556 9042 38724 9044
rect 38556 8990 38558 9042
rect 38610 8990 38724 9042
rect 38556 8988 38724 8990
rect 38556 8978 38612 8988
rect 38668 8820 38724 8988
rect 38444 8764 38612 8820
rect 38444 5908 38500 5918
rect 38444 5814 38500 5852
rect 38332 5506 38388 5516
rect 37548 4274 37604 4284
rect 38332 5124 38388 5134
rect 37324 4174 37326 4226
rect 37378 4174 37380 4226
rect 37324 4162 37380 4174
rect 38220 4226 38276 4238
rect 38220 4174 38222 4226
rect 38274 4174 38276 4226
rect 37212 3390 37214 3442
rect 37266 3390 37268 3442
rect 36204 3332 36372 3388
rect 37212 3378 37268 3390
rect 35532 3266 35588 3276
rect 36316 3266 36372 3276
rect 38220 1764 38276 4174
rect 38332 3778 38388 5068
rect 38444 4900 38500 4910
rect 38556 4900 38612 8764
rect 38668 8754 38724 8764
rect 38780 7812 38836 9100
rect 38892 9042 38948 9324
rect 38892 8990 38894 9042
rect 38946 8990 38948 9042
rect 38892 7924 38948 8990
rect 39116 9042 39172 9054
rect 39116 8990 39118 9042
rect 39170 8990 39172 9042
rect 39004 8930 39060 8942
rect 39004 8878 39006 8930
rect 39058 8878 39060 8930
rect 39004 8708 39060 8878
rect 39004 8642 39060 8652
rect 39116 8484 39172 8990
rect 39004 8428 39172 8484
rect 39004 8258 39060 8428
rect 39004 8206 39006 8258
rect 39058 8206 39060 8258
rect 39004 8148 39060 8206
rect 39228 8260 39284 10446
rect 39340 10386 39396 10398
rect 39340 10334 39342 10386
rect 39394 10334 39396 10386
rect 39340 9044 39396 10334
rect 39564 9156 39620 13468
rect 39676 12852 39732 14364
rect 39788 12964 39844 14924
rect 40012 14756 40068 15262
rect 39900 14644 39956 14654
rect 39900 13746 39956 14588
rect 39900 13694 39902 13746
rect 39954 13694 39956 13746
rect 39900 13682 39956 13694
rect 40012 13636 40068 14700
rect 40012 13570 40068 13580
rect 40124 14418 40180 15484
rect 40124 14366 40126 14418
rect 40178 14366 40180 14418
rect 40124 13076 40180 14366
rect 40236 13748 40292 15596
rect 40348 14868 40404 16828
rect 40348 13972 40404 14812
rect 40348 13906 40404 13916
rect 40460 15314 40516 15326
rect 40460 15262 40462 15314
rect 40514 15262 40516 15314
rect 40236 13692 40404 13748
rect 40236 13524 40292 13534
rect 40236 13430 40292 13468
rect 39788 12908 39956 12964
rect 39676 12796 39844 12852
rect 39676 12404 39732 12414
rect 39676 12178 39732 12348
rect 39676 12126 39678 12178
rect 39730 12126 39732 12178
rect 39676 12114 39732 12126
rect 39788 10834 39844 12796
rect 39788 10782 39790 10834
rect 39842 10782 39844 10834
rect 39788 10770 39844 10782
rect 39900 9940 39956 12908
rect 40012 12404 40068 12414
rect 40124 12404 40180 13020
rect 40012 12402 40180 12404
rect 40012 12350 40014 12402
rect 40066 12350 40180 12402
rect 40012 12348 40180 12350
rect 40012 12338 40068 12348
rect 40348 11394 40404 13692
rect 40460 12964 40516 15262
rect 40460 12898 40516 12908
rect 40572 11396 40628 19516
rect 41244 19506 41300 19516
rect 41356 20356 41412 20366
rect 41020 19236 41076 19246
rect 41020 18674 41076 19180
rect 41020 18622 41022 18674
rect 41074 18622 41076 18674
rect 41020 18610 41076 18622
rect 41356 18228 41412 20300
rect 41020 18226 41412 18228
rect 41020 18174 41358 18226
rect 41410 18174 41412 18226
rect 41020 18172 41412 18174
rect 40796 18004 40852 18014
rect 40796 17556 40852 17948
rect 40796 17462 40852 17500
rect 40908 17556 40964 17566
rect 41020 17556 41076 18172
rect 41356 18162 41412 18172
rect 41468 17890 41524 21644
rect 42028 21588 42084 21598
rect 42028 21494 42084 21532
rect 42252 21364 42308 22204
rect 42700 22194 42756 22204
rect 42364 21700 42420 21710
rect 42364 21606 42420 21644
rect 42812 21476 42868 26908
rect 43484 26964 43540 27002
rect 43484 26898 43540 26908
rect 43596 26962 43652 26974
rect 43596 26910 43598 26962
rect 43650 26910 43652 26962
rect 43820 26964 43876 27580
rect 43372 26852 43428 26862
rect 42924 26628 42980 26638
rect 42924 26514 42980 26572
rect 42924 26462 42926 26514
rect 42978 26462 42980 26514
rect 42924 26450 42980 26462
rect 42924 25506 42980 25518
rect 42924 25454 42926 25506
rect 42978 25454 42980 25506
rect 42924 24164 42980 25454
rect 43148 25396 43204 25406
rect 42924 24098 42980 24108
rect 43036 25394 43204 25396
rect 43036 25342 43150 25394
rect 43202 25342 43204 25394
rect 43036 25340 43204 25342
rect 43036 23492 43092 25340
rect 43148 25330 43204 25340
rect 43148 25060 43204 25070
rect 43148 24946 43204 25004
rect 43148 24894 43150 24946
rect 43202 24894 43204 24946
rect 43148 24882 43204 24894
rect 43036 23426 43092 23436
rect 43036 23154 43092 23166
rect 43036 23102 43038 23154
rect 43090 23102 43092 23154
rect 43036 21924 43092 23102
rect 43036 21858 43092 21868
rect 43260 23156 43316 23166
rect 43260 22372 43316 23100
rect 43148 21812 43204 21822
rect 42924 21476 42980 21486
rect 42812 21474 42980 21476
rect 42812 21422 42926 21474
rect 42978 21422 42980 21474
rect 42812 21420 42980 21422
rect 41916 21308 42308 21364
rect 41692 20578 41748 20590
rect 41692 20526 41694 20578
rect 41746 20526 41748 20578
rect 41692 20244 41748 20526
rect 41692 20178 41748 20188
rect 41804 20356 41860 20366
rect 41804 20130 41860 20300
rect 41804 20078 41806 20130
rect 41858 20078 41860 20130
rect 41804 20066 41860 20078
rect 41468 17838 41470 17890
rect 41522 17838 41524 17890
rect 41468 17826 41524 17838
rect 41580 19684 41636 19694
rect 41132 17668 41188 17678
rect 41132 17574 41188 17612
rect 41356 17668 41412 17678
rect 41580 17668 41636 19628
rect 41356 17666 41636 17668
rect 41356 17614 41358 17666
rect 41410 17614 41636 17666
rect 41356 17612 41636 17614
rect 40908 17554 41076 17556
rect 40908 17502 40910 17554
rect 40962 17502 41076 17554
rect 40908 17500 41076 17502
rect 41356 17556 41412 17612
rect 40908 17490 40964 17500
rect 41356 17490 41412 17500
rect 41468 17444 41524 17454
rect 41916 17444 41972 21308
rect 42924 20916 42980 21420
rect 42700 20860 42980 20916
rect 42140 20804 42196 20814
rect 42700 20804 42756 20860
rect 42028 20748 42140 20804
rect 42028 19458 42084 20748
rect 42140 20738 42196 20748
rect 42476 20748 42756 20804
rect 43036 20804 43092 20814
rect 42252 20690 42308 20702
rect 42252 20638 42254 20690
rect 42306 20638 42308 20690
rect 42252 20356 42308 20638
rect 42252 20290 42308 20300
rect 42364 20580 42420 20590
rect 42028 19406 42030 19458
rect 42082 19406 42084 19458
rect 42028 18562 42084 19406
rect 42252 19348 42308 19358
rect 42252 19254 42308 19292
rect 42364 19234 42420 20524
rect 42364 19182 42366 19234
rect 42418 19182 42420 19234
rect 42364 19170 42420 19182
rect 42028 18510 42030 18562
rect 42082 18510 42084 18562
rect 42028 18498 42084 18510
rect 42140 18452 42196 18462
rect 42140 18358 42196 18396
rect 42252 17556 42308 17566
rect 42252 17462 42308 17500
rect 41468 17442 41972 17444
rect 41468 17390 41470 17442
rect 41522 17390 41972 17442
rect 41468 17388 41972 17390
rect 41468 17378 41524 17388
rect 41356 16996 41412 17006
rect 41244 16994 41412 16996
rect 41244 16942 41358 16994
rect 41410 16942 41412 16994
rect 41244 16940 41412 16942
rect 41132 16884 41188 16894
rect 41132 16790 41188 16828
rect 40684 16772 40740 16782
rect 40684 13300 40740 16716
rect 41244 16100 41300 16940
rect 41356 16930 41412 16940
rect 41916 16994 41972 17006
rect 41916 16942 41918 16994
rect 41970 16942 41972 16994
rect 41468 16884 41524 16894
rect 41468 16882 41636 16884
rect 41468 16830 41470 16882
rect 41522 16830 41636 16882
rect 41468 16828 41636 16830
rect 41468 16818 41524 16828
rect 41468 16212 41524 16222
rect 41468 16118 41524 16156
rect 41244 16044 41412 16100
rect 40796 14980 40852 14990
rect 40796 14308 40852 14924
rect 40908 14644 40964 14654
rect 40908 14530 40964 14588
rect 41244 14644 41300 14654
rect 41356 14644 41412 16044
rect 41468 15426 41524 15438
rect 41468 15374 41470 15426
rect 41522 15374 41524 15426
rect 41468 15204 41524 15374
rect 41580 15204 41636 16828
rect 41804 16882 41860 16894
rect 41804 16830 41806 16882
rect 41858 16830 41860 16882
rect 41804 15764 41860 16830
rect 41916 16212 41972 16942
rect 42140 16884 42196 16894
rect 42140 16882 42308 16884
rect 42140 16830 42142 16882
rect 42194 16830 42308 16882
rect 42140 16828 42308 16830
rect 42140 16818 42196 16828
rect 41916 16210 42084 16212
rect 41916 16158 41918 16210
rect 41970 16158 42084 16210
rect 41916 16156 42084 16158
rect 41916 16146 41972 16156
rect 42028 16100 42084 16156
rect 42252 16100 42308 16828
rect 42476 16772 42532 20748
rect 43036 20710 43092 20748
rect 42812 20692 42868 20702
rect 42812 20690 42980 20692
rect 42812 20638 42814 20690
rect 42866 20638 42980 20690
rect 42812 20636 42980 20638
rect 42812 20626 42868 20636
rect 42924 20580 42980 20636
rect 42924 20244 42980 20524
rect 43148 20356 43204 21756
rect 43260 21810 43316 22316
rect 43260 21758 43262 21810
rect 43314 21758 43316 21810
rect 43260 21746 43316 21758
rect 43372 20804 43428 26796
rect 43484 25394 43540 25406
rect 43484 25342 43486 25394
rect 43538 25342 43540 25394
rect 43484 22484 43540 25342
rect 43596 25284 43652 26910
rect 43708 26906 43764 26918
rect 43708 26854 43710 26906
rect 43762 26854 43764 26906
rect 43820 26898 43876 26908
rect 43708 26292 43764 26854
rect 43932 26850 43988 26862
rect 43932 26798 43934 26850
rect 43986 26798 43988 26850
rect 43708 26226 43764 26236
rect 43820 26628 43876 26638
rect 43596 25218 43652 25228
rect 43484 22418 43540 22428
rect 43596 23828 43652 23838
rect 43596 22036 43652 23772
rect 43596 21970 43652 21980
rect 43820 21700 43876 26572
rect 43932 23380 43988 26798
rect 44044 26068 44100 27918
rect 44156 27858 44212 29148
rect 44156 27806 44158 27858
rect 44210 27806 44212 27858
rect 44156 27794 44212 27806
rect 44380 26908 44436 30828
rect 45052 29988 45108 29998
rect 45052 29894 45108 29932
rect 46060 29988 46116 29998
rect 46060 29428 46116 29932
rect 46060 29362 46116 29372
rect 46284 29426 46340 31164
rect 46284 29374 46286 29426
rect 46338 29374 46340 29426
rect 46284 29362 46340 29374
rect 46396 31218 46564 31220
rect 46396 31166 46510 31218
rect 46562 31166 46564 31218
rect 46396 31164 46564 31166
rect 46396 29988 46452 31164
rect 46508 31154 46564 31164
rect 46620 31778 46676 31790
rect 46620 31726 46622 31778
rect 46674 31726 46676 31778
rect 46620 30436 46676 31726
rect 47068 31218 47124 33516
rect 47292 33460 47348 37436
rect 47516 37266 47572 37660
rect 47516 37214 47518 37266
rect 47570 37214 47572 37266
rect 47516 37202 47572 37214
rect 47628 36484 47684 38556
rect 48076 38276 48132 43374
rect 48188 42194 48244 43486
rect 48188 42142 48190 42194
rect 48242 42142 48244 42194
rect 48188 42130 48244 42142
rect 48412 42196 48468 46956
rect 48636 46946 48692 46956
rect 48748 47124 48804 47134
rect 48636 44324 48692 44334
rect 48524 44322 48692 44324
rect 48524 44270 48638 44322
rect 48690 44270 48692 44322
rect 48524 44268 48692 44270
rect 48748 44324 48804 47068
rect 48972 47012 49028 48300
rect 48972 46946 49028 46956
rect 48972 46674 49028 46686
rect 48972 46622 48974 46674
rect 49026 46622 49028 46674
rect 48972 45332 49028 46622
rect 49196 46004 49252 48524
rect 49420 48468 49476 49308
rect 49308 48412 49476 48468
rect 49308 46898 49364 48412
rect 49420 48242 49476 48254
rect 49420 48190 49422 48242
rect 49474 48190 49476 48242
rect 49420 48020 49476 48190
rect 49420 47236 49476 47964
rect 49420 47170 49476 47180
rect 49532 47458 49588 47470
rect 49532 47406 49534 47458
rect 49586 47406 49588 47458
rect 49308 46846 49310 46898
rect 49362 46846 49364 46898
rect 49308 46834 49364 46846
rect 49420 46900 49476 46910
rect 49420 46786 49476 46844
rect 49420 46734 49422 46786
rect 49474 46734 49476 46786
rect 49420 46722 49476 46734
rect 49532 46788 49588 47406
rect 49532 46722 49588 46732
rect 49756 46228 49812 49532
rect 49868 49028 49924 49038
rect 49868 48934 49924 48972
rect 49868 48356 49924 48366
rect 49868 48130 49924 48300
rect 49980 48354 50036 50204
rect 49980 48302 49982 48354
rect 50034 48302 50036 48354
rect 49980 48290 50036 48302
rect 49868 48078 49870 48130
rect 49922 48078 49924 48130
rect 49868 48066 49924 48078
rect 50092 47684 50148 52334
rect 50204 50148 50260 52668
rect 50316 52164 50372 55246
rect 50428 55858 50484 55870
rect 50428 55806 50430 55858
rect 50482 55806 50484 55858
rect 50428 54514 50484 55806
rect 50540 55412 50596 56030
rect 50540 55346 50596 55356
rect 50876 55076 50932 57484
rect 50988 57538 51044 57550
rect 50988 57486 50990 57538
rect 51042 57486 51044 57538
rect 50988 56084 51044 57486
rect 50988 56018 51044 56028
rect 51100 57316 51156 57326
rect 50876 55010 50932 55020
rect 50988 55412 51044 55422
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50428 54462 50430 54514
rect 50482 54462 50484 54514
rect 50428 54450 50484 54462
rect 50876 54740 50932 54750
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50316 52098 50372 52108
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50876 51604 50932 54684
rect 50988 53730 51044 55356
rect 51100 53842 51156 57260
rect 51212 55076 51268 55086
rect 51212 54982 51268 55020
rect 51100 53790 51102 53842
rect 51154 53790 51156 53842
rect 51100 53778 51156 53790
rect 50988 53678 50990 53730
rect 51042 53678 51044 53730
rect 50988 53666 51044 53678
rect 51212 53620 51268 53630
rect 51212 53526 51268 53564
rect 51324 53172 51380 58156
rect 51436 57650 51492 57662
rect 51436 57598 51438 57650
rect 51490 57598 51492 57650
rect 51436 57090 51492 57598
rect 51436 57038 51438 57090
rect 51490 57038 51492 57090
rect 51436 55412 51492 57038
rect 51436 55346 51492 55356
rect 51212 53116 51380 53172
rect 51436 53508 51492 53518
rect 50988 52948 51044 52958
rect 50988 52854 51044 52892
rect 50652 51548 50932 51604
rect 51100 52834 51156 52846
rect 51100 52782 51102 52834
rect 51154 52782 51156 52834
rect 50316 51492 50372 51502
rect 50316 50594 50372 51436
rect 50316 50542 50318 50594
rect 50370 50542 50372 50594
rect 50316 50148 50372 50542
rect 50652 50594 50708 51548
rect 51100 51156 51156 52782
rect 50764 51100 51156 51156
rect 50764 50820 50820 51100
rect 50764 50754 50820 50764
rect 50876 50820 50932 50830
rect 50876 50818 51156 50820
rect 50876 50766 50878 50818
rect 50930 50766 51156 50818
rect 50876 50764 51156 50766
rect 50876 50754 50932 50764
rect 50652 50542 50654 50594
rect 50706 50542 50708 50594
rect 50652 50428 50708 50542
rect 50988 50596 51044 50606
rect 50988 50502 51044 50540
rect 50428 50372 50484 50382
rect 50652 50372 50932 50428
rect 50428 50278 50484 50316
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50316 50092 50484 50148
rect 50556 50138 50820 50148
rect 50204 50082 50260 50092
rect 50204 49924 50260 49934
rect 50204 49026 50260 49868
rect 50428 49812 50484 50092
rect 50764 49812 50820 49822
rect 50876 49812 50932 50372
rect 50428 49810 50596 49812
rect 50428 49758 50430 49810
rect 50482 49758 50596 49810
rect 50428 49756 50596 49758
rect 50428 49746 50484 49756
rect 50428 49252 50484 49262
rect 50204 48974 50206 49026
rect 50258 48974 50260 49026
rect 50204 48962 50260 48974
rect 50316 49196 50428 49252
rect 49980 47628 50148 47684
rect 49980 47346 50036 47628
rect 50316 47572 50372 49196
rect 50428 49186 50484 49196
rect 50540 48916 50596 49756
rect 50764 49810 50932 49812
rect 50764 49758 50766 49810
rect 50818 49758 50932 49810
rect 50764 49756 50932 49758
rect 50988 50148 51044 50158
rect 50988 49810 51044 50092
rect 50988 49758 50990 49810
rect 51042 49758 51044 49810
rect 50764 49028 50820 49756
rect 50988 49746 51044 49758
rect 50876 49588 50932 49598
rect 51100 49588 51156 50764
rect 51212 50708 51268 53116
rect 51324 52946 51380 52958
rect 51324 52894 51326 52946
rect 51378 52894 51380 52946
rect 51324 52388 51380 52894
rect 51436 52724 51492 53452
rect 51548 53172 51604 58268
rect 51660 58212 51716 58222
rect 51660 58118 51716 58156
rect 51884 57762 51940 57774
rect 51884 57710 51886 57762
rect 51938 57710 51940 57762
rect 51884 57652 51940 57710
rect 52108 57764 52164 57774
rect 52108 57670 52164 57708
rect 51884 57586 51940 57596
rect 52332 57650 52388 57662
rect 52556 57652 52612 57662
rect 52332 57598 52334 57650
rect 52386 57598 52388 57650
rect 51772 57426 51828 57438
rect 51772 57374 51774 57426
rect 51826 57374 51828 57426
rect 51660 56308 51716 56318
rect 51660 56214 51716 56252
rect 51660 55074 51716 55086
rect 51660 55022 51662 55074
rect 51714 55022 51716 55074
rect 51660 54964 51716 55022
rect 51660 54898 51716 54908
rect 51660 54516 51716 54526
rect 51660 54422 51716 54460
rect 51660 53620 51716 53630
rect 51660 53526 51716 53564
rect 51772 53508 51828 57374
rect 52332 57428 52388 57598
rect 52332 57362 52388 57372
rect 52444 57650 52612 57652
rect 52444 57598 52558 57650
rect 52610 57598 52612 57650
rect 52444 57596 52612 57598
rect 52220 56642 52276 56654
rect 52220 56590 52222 56642
rect 52274 56590 52276 56642
rect 52220 55636 52276 56590
rect 52220 55570 52276 55580
rect 51884 55074 51940 55086
rect 51884 55022 51886 55074
rect 51938 55022 51940 55074
rect 51884 53844 51940 55022
rect 51996 55076 52052 55086
rect 51996 54982 52052 55020
rect 52108 55076 52164 55086
rect 52108 55074 52276 55076
rect 52108 55022 52110 55074
rect 52162 55022 52276 55074
rect 52108 55020 52276 55022
rect 52108 55010 52164 55020
rect 52108 54628 52164 54638
rect 52108 54534 52164 54572
rect 51884 53778 51940 53788
rect 52108 54404 52164 54414
rect 51996 53732 52052 53742
rect 52108 53732 52164 54348
rect 51996 53730 52164 53732
rect 51996 53678 51998 53730
rect 52050 53678 52164 53730
rect 51996 53676 52164 53678
rect 51996 53666 52052 53676
rect 51772 53452 52052 53508
rect 51548 53116 51828 53172
rect 51548 52948 51604 52958
rect 51548 52946 51716 52948
rect 51548 52894 51550 52946
rect 51602 52894 51716 52946
rect 51548 52892 51716 52894
rect 51548 52882 51604 52892
rect 51548 52724 51604 52734
rect 51436 52668 51548 52724
rect 51324 52322 51380 52332
rect 51212 50642 51268 50652
rect 51324 52164 51380 52174
rect 50876 49586 51156 49588
rect 50876 49534 50878 49586
rect 50930 49534 51156 49586
rect 50876 49532 51156 49534
rect 51212 50034 51268 50046
rect 51212 49982 51214 50034
rect 51266 49982 51268 50034
rect 50876 49140 50932 49532
rect 50876 49074 50932 49084
rect 50764 48934 50820 48972
rect 50652 48916 50708 48926
rect 50540 48914 50708 48916
rect 50540 48862 50654 48914
rect 50706 48862 50708 48914
rect 50540 48860 50708 48862
rect 50652 48850 50708 48860
rect 51100 48804 51156 48814
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50876 48356 50932 48366
rect 50652 48244 50708 48254
rect 50652 48242 50820 48244
rect 50652 48190 50654 48242
rect 50706 48190 50820 48242
rect 50652 48188 50820 48190
rect 50652 48178 50708 48188
rect 50652 47796 50708 47806
rect 49980 47294 49982 47346
rect 50034 47294 50036 47346
rect 49196 45938 49252 45948
rect 49420 46172 49812 46228
rect 49868 46786 49924 46798
rect 49868 46734 49870 46786
rect 49922 46734 49924 46786
rect 48972 45276 49252 45332
rect 48860 45220 48916 45230
rect 48860 45126 48916 45164
rect 48972 45108 49028 45118
rect 48972 45014 49028 45052
rect 48860 44882 48916 44894
rect 48860 44830 48862 44882
rect 48914 44830 48916 44882
rect 48860 44548 48916 44830
rect 48860 44482 48916 44492
rect 48748 44268 48916 44324
rect 48524 43652 48580 44268
rect 48636 44258 48692 44268
rect 48748 44100 48804 44110
rect 48524 43586 48580 43596
rect 48636 44044 48748 44100
rect 48412 42130 48468 42140
rect 48636 41186 48692 44044
rect 48748 44006 48804 44044
rect 48748 43876 48804 43886
rect 48748 42308 48804 43820
rect 48860 43428 48916 44268
rect 49196 44322 49252 45276
rect 49420 44884 49476 46172
rect 49756 46004 49812 46014
rect 49756 45778 49812 45948
rect 49756 45726 49758 45778
rect 49810 45726 49812 45778
rect 49756 45714 49812 45726
rect 49532 45220 49588 45230
rect 49532 44996 49588 45164
rect 49868 45220 49924 46734
rect 49868 45154 49924 45164
rect 49980 45218 50036 47294
rect 50092 47516 50372 47572
rect 50428 47740 50652 47796
rect 50092 47346 50148 47516
rect 50092 47294 50094 47346
rect 50146 47294 50148 47346
rect 50092 45892 50148 47294
rect 50204 47348 50260 47358
rect 50204 47254 50260 47292
rect 50316 47234 50372 47246
rect 50316 47182 50318 47234
rect 50370 47182 50372 47234
rect 50316 47012 50372 47182
rect 50092 45798 50148 45836
rect 50204 46900 50260 46910
rect 49980 45166 49982 45218
rect 50034 45166 50036 45218
rect 49980 45154 50036 45166
rect 50092 45556 50148 45566
rect 49532 44940 49700 44996
rect 49420 44828 49588 44884
rect 49196 44270 49198 44322
rect 49250 44270 49252 44322
rect 49196 44212 49252 44270
rect 49084 44156 49252 44212
rect 48860 43426 49028 43428
rect 48860 43374 48862 43426
rect 48914 43374 49028 43426
rect 48860 43372 49028 43374
rect 48860 43362 48916 43372
rect 48860 42308 48916 42318
rect 48748 42252 48860 42308
rect 48636 41134 48638 41186
rect 48690 41134 48692 41186
rect 48636 41122 48692 41134
rect 48860 40292 48916 42252
rect 48972 41860 49028 43372
rect 49084 43092 49140 44156
rect 49084 43026 49140 43036
rect 49196 43764 49252 43774
rect 48972 41076 49028 41804
rect 48972 41010 49028 41020
rect 48860 40226 48916 40236
rect 48748 40178 48804 40190
rect 48748 40126 48750 40178
rect 48802 40126 48804 40178
rect 48748 39620 48804 40126
rect 48748 39508 48804 39564
rect 49084 40178 49140 40190
rect 49084 40126 49086 40178
rect 49138 40126 49140 40178
rect 49084 40068 49140 40126
rect 48860 39508 48916 39518
rect 48748 39506 48916 39508
rect 48748 39454 48862 39506
rect 48914 39454 48916 39506
rect 48748 39452 48916 39454
rect 48860 39442 48916 39452
rect 48748 38948 48804 38958
rect 48748 38854 48804 38892
rect 49084 38834 49140 40012
rect 49084 38782 49086 38834
rect 49138 38782 49140 38834
rect 49084 38770 49140 38782
rect 49196 38722 49252 43708
rect 49308 43652 49364 43662
rect 49308 43558 49364 43596
rect 49308 43428 49364 43438
rect 49308 40514 49364 43372
rect 49420 42530 49476 42542
rect 49420 42478 49422 42530
rect 49474 42478 49476 42530
rect 49420 42084 49476 42478
rect 49420 41990 49476 42028
rect 49308 40462 49310 40514
rect 49362 40462 49364 40514
rect 49308 40450 49364 40462
rect 49532 40404 49588 44828
rect 49644 44212 49700 44940
rect 49644 44146 49700 44156
rect 49756 44548 49812 44558
rect 49756 43538 49812 44492
rect 49756 43486 49758 43538
rect 49810 43486 49812 43538
rect 49756 43474 49812 43486
rect 50092 43426 50148 45500
rect 50204 43652 50260 46844
rect 50316 46116 50372 46956
rect 50428 46898 50484 47740
rect 50652 47730 50708 47740
rect 50764 47684 50820 48188
rect 50876 47908 50932 48300
rect 50876 47842 50932 47852
rect 50764 47628 51044 47684
rect 50876 47346 50932 47358
rect 50876 47294 50878 47346
rect 50930 47294 50932 47346
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50428 46846 50430 46898
rect 50482 46846 50484 46898
rect 50428 46452 50484 46846
rect 50428 46386 50484 46396
rect 50540 46674 50596 46686
rect 50540 46622 50542 46674
rect 50594 46622 50596 46674
rect 50540 46228 50596 46622
rect 50316 46050 50372 46060
rect 50428 46172 50596 46228
rect 50428 46004 50484 46172
rect 50428 45938 50484 45948
rect 50764 46116 50820 46126
rect 50540 45892 50596 45902
rect 50764 45892 50820 46060
rect 50540 45890 50820 45892
rect 50540 45838 50542 45890
rect 50594 45838 50820 45890
rect 50540 45836 50820 45838
rect 50876 45892 50932 47294
rect 50988 47124 51044 47628
rect 51100 47346 51156 48748
rect 51212 48468 51268 49982
rect 51324 49252 51380 52108
rect 51548 52050 51604 52668
rect 51548 51998 51550 52050
rect 51602 51998 51604 52050
rect 51548 51986 51604 51998
rect 51548 50820 51604 50830
rect 51660 50820 51716 52892
rect 51772 51940 51828 53116
rect 51996 52946 52052 53452
rect 51996 52894 51998 52946
rect 52050 52894 52052 52946
rect 51996 52882 52052 52894
rect 52108 52834 52164 52846
rect 52108 52782 52110 52834
rect 52162 52782 52164 52834
rect 51884 52164 51940 52174
rect 51884 52162 52052 52164
rect 51884 52110 51886 52162
rect 51938 52110 52052 52162
rect 51884 52108 52052 52110
rect 51884 52098 51940 52108
rect 51772 51884 51940 51940
rect 51660 50764 51828 50820
rect 51436 50708 51492 50718
rect 51436 50594 51492 50652
rect 51436 50542 51438 50594
rect 51490 50542 51492 50594
rect 51436 50530 51492 50542
rect 51548 50596 51604 50764
rect 51660 50596 51716 50606
rect 51548 50594 51716 50596
rect 51548 50542 51662 50594
rect 51714 50542 51716 50594
rect 51548 50540 51716 50542
rect 51660 50530 51716 50540
rect 51772 50428 51828 50764
rect 51436 50372 51492 50382
rect 51436 50034 51492 50316
rect 51436 49982 51438 50034
rect 51490 49982 51492 50034
rect 51436 49970 51492 49982
rect 51548 50370 51604 50382
rect 51548 50318 51550 50370
rect 51602 50318 51604 50370
rect 51436 49252 51492 49262
rect 51324 49250 51492 49252
rect 51324 49198 51438 49250
rect 51490 49198 51492 49250
rect 51324 49196 51492 49198
rect 51436 49186 51492 49196
rect 51548 49028 51604 50318
rect 51660 50372 51828 50428
rect 51884 50484 51940 51884
rect 51884 50418 51940 50428
rect 51660 50148 51716 50372
rect 51660 50082 51716 50092
rect 51772 50260 51828 50270
rect 51660 49922 51716 49934
rect 51660 49870 51662 49922
rect 51714 49870 51716 49922
rect 51660 49588 51716 49870
rect 51772 49922 51828 50204
rect 51772 49870 51774 49922
rect 51826 49870 51828 49922
rect 51772 49858 51828 49870
rect 51660 49522 51716 49532
rect 51996 49140 52052 52108
rect 52108 51492 52164 52782
rect 52220 52276 52276 55020
rect 52444 54404 52500 57596
rect 52556 57586 52612 57596
rect 52892 57652 52948 58492
rect 62188 58482 62244 58492
rect 53228 58210 53284 58222
rect 54460 58212 54516 58222
rect 53228 58158 53230 58210
rect 53282 58158 53284 58210
rect 52780 57540 52836 57550
rect 52780 57446 52836 57484
rect 52892 56868 52948 57596
rect 53116 57650 53172 57662
rect 53116 57598 53118 57650
rect 53170 57598 53172 57650
rect 53116 57316 53172 57598
rect 53116 57250 53172 57260
rect 53228 57652 53284 58158
rect 54348 58210 54516 58212
rect 54348 58158 54462 58210
rect 54514 58158 54516 58210
rect 54348 58156 54516 58158
rect 53788 57764 53844 57774
rect 52444 54180 52500 54348
rect 52444 52834 52500 54124
rect 52556 56812 52948 56868
rect 52556 53620 52612 56812
rect 52892 56644 52948 56654
rect 52892 56550 52948 56588
rect 53116 55860 53172 55870
rect 53228 55860 53284 57596
rect 53116 55858 53284 55860
rect 53116 55806 53118 55858
rect 53170 55806 53284 55858
rect 53116 55804 53284 55806
rect 53564 57650 53620 57662
rect 53564 57598 53566 57650
rect 53618 57598 53620 57650
rect 53564 57428 53620 57598
rect 53788 57650 53844 57708
rect 53788 57598 53790 57650
rect 53842 57598 53844 57650
rect 53788 57586 53844 57598
rect 54012 57652 54068 57662
rect 54012 57558 54068 57596
rect 52668 55298 52724 55310
rect 52668 55246 52670 55298
rect 52722 55246 52724 55298
rect 52668 54740 52724 55246
rect 52668 54674 52724 54684
rect 52780 54628 52836 54638
rect 53116 54628 53172 55804
rect 53564 55412 53620 57372
rect 53676 57538 53732 57550
rect 53676 57486 53678 57538
rect 53730 57486 53732 57538
rect 53676 57316 53732 57486
rect 53676 57250 53732 57260
rect 53788 56754 53844 56766
rect 53788 56702 53790 56754
rect 53842 56702 53844 56754
rect 53788 56308 53844 56702
rect 53788 56242 53844 56252
rect 54236 55972 54292 55982
rect 54348 55972 54404 58156
rect 54460 58146 54516 58156
rect 55356 57876 55412 57886
rect 55020 57540 55076 57550
rect 55020 57446 55076 57484
rect 54236 55970 54404 55972
rect 54236 55918 54238 55970
rect 54290 55918 54404 55970
rect 54236 55916 54404 55918
rect 54460 57426 54516 57438
rect 54460 57374 54462 57426
rect 54514 57374 54516 57426
rect 53564 55356 53732 55412
rect 53228 55300 53284 55310
rect 53228 55206 53284 55244
rect 53452 55076 53508 55086
rect 53228 54628 53284 54638
rect 53116 54626 53284 54628
rect 53116 54574 53230 54626
rect 53282 54574 53284 54626
rect 53116 54572 53284 54574
rect 52780 54534 52836 54572
rect 53228 54404 53284 54572
rect 53452 54514 53508 55020
rect 53452 54462 53454 54514
rect 53506 54462 53508 54514
rect 53452 54450 53508 54462
rect 53564 55074 53620 55086
rect 53564 55022 53566 55074
rect 53618 55022 53620 55074
rect 53564 54964 53620 55022
rect 53676 55076 53732 55356
rect 53900 55300 53956 55310
rect 53956 55244 54068 55300
rect 53900 55206 53956 55244
rect 53676 55010 53732 55020
rect 53228 54338 53284 54348
rect 52892 54292 52948 54302
rect 52892 53954 52948 54236
rect 52892 53902 52894 53954
rect 52946 53902 52948 53954
rect 52892 53890 52948 53902
rect 53564 53844 53620 54908
rect 53340 53788 53620 53844
rect 53676 54628 53732 54638
rect 52892 53732 52948 53742
rect 52948 53676 53060 53732
rect 52892 53666 52948 53676
rect 52556 52946 52612 53564
rect 52668 53618 52724 53630
rect 52668 53566 52670 53618
rect 52722 53566 52724 53618
rect 52668 53172 52724 53566
rect 52668 53106 52724 53116
rect 52556 52894 52558 52946
rect 52610 52894 52612 52946
rect 52556 52882 52612 52894
rect 52444 52782 52446 52834
rect 52498 52782 52500 52834
rect 52444 52770 52500 52782
rect 52220 52210 52276 52220
rect 52892 52500 52948 52510
rect 52556 52162 52612 52174
rect 52556 52110 52558 52162
rect 52610 52110 52612 52162
rect 52108 51426 52164 51436
rect 52444 51940 52500 51950
rect 52108 51266 52164 51278
rect 52108 51214 52110 51266
rect 52162 51214 52164 51266
rect 52108 51156 52164 51214
rect 52108 51090 52164 51100
rect 52444 50428 52500 51884
rect 51996 49074 52052 49084
rect 52108 50372 52500 50428
rect 51548 48972 51940 49028
rect 51772 48804 51828 48814
rect 51772 48710 51828 48748
rect 51212 48412 51716 48468
rect 51212 48242 51268 48254
rect 51212 48190 51214 48242
rect 51266 48190 51268 48242
rect 51212 47684 51268 48190
rect 51436 48242 51492 48254
rect 51436 48190 51438 48242
rect 51490 48190 51492 48242
rect 51324 48132 51380 48142
rect 51324 48038 51380 48076
rect 51436 47796 51492 48190
rect 51436 47730 51492 47740
rect 51660 47684 51716 48412
rect 51772 48244 51828 48254
rect 51772 48150 51828 48188
rect 51772 47684 51828 47694
rect 51660 47682 51828 47684
rect 51660 47630 51774 47682
rect 51826 47630 51828 47682
rect 51660 47628 51828 47630
rect 51212 47618 51268 47628
rect 51772 47618 51828 47628
rect 51324 47572 51380 47582
rect 51324 47478 51380 47516
rect 51436 47460 51492 47470
rect 51884 47460 51940 48972
rect 51436 47458 51940 47460
rect 51436 47406 51438 47458
rect 51490 47406 51940 47458
rect 51436 47404 51940 47406
rect 52108 47458 52164 50372
rect 52556 49700 52612 52110
rect 52780 52164 52836 52174
rect 52780 52070 52836 52108
rect 52892 52162 52948 52444
rect 52892 52110 52894 52162
rect 52946 52110 52948 52162
rect 52892 52098 52948 52110
rect 53004 51380 53060 53676
rect 53228 53506 53284 53518
rect 53228 53454 53230 53506
rect 53282 53454 53284 53506
rect 53228 52724 53284 53454
rect 53228 52658 53284 52668
rect 53228 52500 53284 52510
rect 53004 50594 53060 51324
rect 53004 50542 53006 50594
rect 53058 50542 53060 50594
rect 53004 50530 53060 50542
rect 53116 52162 53172 52174
rect 53116 52110 53118 52162
rect 53170 52110 53172 52162
rect 52556 49634 52612 49644
rect 52892 49922 52948 49934
rect 52892 49870 52894 49922
rect 52946 49870 52948 49922
rect 52892 49252 52948 49870
rect 53116 49924 53172 52110
rect 53228 51268 53284 52444
rect 53340 51490 53396 53788
rect 53676 53732 53732 54572
rect 53788 54516 53844 54526
rect 53788 54422 53844 54460
rect 53564 53730 53732 53732
rect 53564 53678 53678 53730
rect 53730 53678 53732 53730
rect 53564 53676 53732 53678
rect 53564 53170 53620 53676
rect 53676 53666 53732 53676
rect 53788 53732 53844 53742
rect 53788 53172 53844 53676
rect 53564 53118 53566 53170
rect 53618 53118 53620 53170
rect 53564 53106 53620 53118
rect 53676 53170 53844 53172
rect 53676 53118 53790 53170
rect 53842 53118 53844 53170
rect 53676 53116 53844 53118
rect 53452 52948 53508 52958
rect 53676 52948 53732 53116
rect 53788 53106 53844 53116
rect 53900 53172 53956 53182
rect 53900 53058 53956 53116
rect 53900 53006 53902 53058
rect 53954 53006 53956 53058
rect 53900 52994 53956 53006
rect 53452 52162 53508 52892
rect 53452 52110 53454 52162
rect 53506 52110 53508 52162
rect 53452 52098 53508 52110
rect 53564 52892 53732 52948
rect 53340 51438 53342 51490
rect 53394 51438 53396 51490
rect 53340 51426 53396 51438
rect 53564 51378 53620 52892
rect 54012 52612 54068 55244
rect 53788 52556 54068 52612
rect 54124 55186 54180 55198
rect 54124 55134 54126 55186
rect 54178 55134 54180 55186
rect 53676 51940 53732 51950
rect 53676 51846 53732 51884
rect 53564 51326 53566 51378
rect 53618 51326 53620 51378
rect 53564 51314 53620 51326
rect 53228 51212 53396 51268
rect 53228 50708 53284 50718
rect 53228 50614 53284 50652
rect 53340 50428 53396 51212
rect 53564 51044 53620 51054
rect 53564 50596 53620 50988
rect 53340 50372 53508 50428
rect 53116 49858 53172 49868
rect 53228 50036 53284 50046
rect 53228 49700 53284 49980
rect 52892 49186 52948 49196
rect 53116 49644 53284 49700
rect 52780 49140 52836 49150
rect 52780 49046 52836 49084
rect 52892 49026 52948 49038
rect 52892 48974 52894 49026
rect 52946 48974 52948 49026
rect 52556 48916 52612 48926
rect 52444 48354 52500 48366
rect 52444 48302 52446 48354
rect 52498 48302 52500 48354
rect 52444 47572 52500 48302
rect 52444 47506 52500 47516
rect 52108 47406 52110 47458
rect 52162 47406 52164 47458
rect 51436 47394 51492 47404
rect 52108 47394 52164 47406
rect 51100 47294 51102 47346
rect 51154 47294 51156 47346
rect 51100 47282 51156 47294
rect 51212 47234 51268 47246
rect 51212 47182 51214 47234
rect 51266 47182 51268 47234
rect 51212 47124 51268 47182
rect 50988 47068 51268 47124
rect 51212 46228 51268 47068
rect 51884 47234 51940 47246
rect 52556 47236 52612 48860
rect 51884 47182 51886 47234
rect 51938 47182 51940 47234
rect 51436 46788 51492 46798
rect 51436 46340 51492 46732
rect 51548 46788 51604 46798
rect 51884 46788 51940 47182
rect 51548 46786 51940 46788
rect 51548 46734 51550 46786
rect 51602 46734 51940 46786
rect 51548 46732 51940 46734
rect 52444 47180 52612 47236
rect 52668 47234 52724 47246
rect 52668 47182 52670 47234
rect 52722 47182 52724 47234
rect 51548 46722 51604 46732
rect 51884 46340 51940 46350
rect 51436 46284 51716 46340
rect 51212 46162 51268 46172
rect 51436 46116 51492 46126
rect 51212 45892 51268 45902
rect 50876 45836 51156 45892
rect 50540 45780 50596 45836
rect 50428 45724 50596 45780
rect 50428 45332 50484 45724
rect 50876 45668 50932 45678
rect 50876 45666 51044 45668
rect 50876 45614 50878 45666
rect 50930 45614 51044 45666
rect 50876 45612 51044 45614
rect 50876 45602 50932 45612
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50428 45276 50596 45332
rect 50316 45108 50372 45118
rect 50316 45014 50372 45052
rect 50428 44324 50484 44334
rect 50428 44230 50484 44268
rect 50540 44100 50596 45276
rect 50652 44882 50708 44894
rect 50652 44830 50654 44882
rect 50706 44830 50708 44882
rect 50652 44436 50708 44830
rect 50652 44370 50708 44380
rect 50988 44322 51044 45612
rect 51100 45108 51156 45836
rect 51100 45042 51156 45052
rect 51212 45106 51268 45836
rect 51212 45054 51214 45106
rect 51266 45054 51268 45106
rect 51212 45042 51268 45054
rect 51324 45890 51380 45902
rect 51324 45838 51326 45890
rect 51378 45838 51380 45890
rect 50988 44270 50990 44322
rect 51042 44270 51044 44322
rect 50204 43586 50260 43596
rect 50428 44044 50596 44100
rect 50652 44210 50708 44222
rect 50652 44158 50654 44210
rect 50706 44158 50708 44210
rect 50652 44100 50708 44158
rect 50092 43374 50094 43426
rect 50146 43374 50148 43426
rect 50092 41972 50148 43374
rect 50092 41186 50148 41916
rect 50092 41134 50094 41186
rect 50146 41134 50148 41186
rect 50092 41122 50148 41134
rect 50316 42084 50372 42094
rect 49868 41076 49924 41086
rect 49868 40982 49924 41020
rect 50092 40964 50148 40974
rect 50092 40962 50260 40964
rect 50092 40910 50094 40962
rect 50146 40910 50260 40962
rect 50092 40908 50260 40910
rect 50092 40898 50148 40908
rect 49980 40516 50036 40526
rect 50036 40460 50148 40516
rect 49980 40422 50036 40460
rect 49644 40404 49700 40414
rect 49532 40402 49700 40404
rect 49532 40350 49646 40402
rect 49698 40350 49700 40402
rect 49532 40348 49700 40350
rect 49644 40180 49700 40348
rect 49644 40114 49700 40124
rect 49756 40404 49812 40414
rect 49196 38670 49198 38722
rect 49250 38670 49252 38722
rect 49196 38658 49252 38670
rect 49308 39842 49364 39854
rect 49308 39790 49310 39842
rect 49362 39790 49364 39842
rect 48076 38210 48132 38220
rect 48188 38612 48244 38622
rect 47964 38164 48020 38174
rect 47852 37938 47908 37950
rect 47852 37886 47854 37938
rect 47906 37886 47908 37938
rect 47852 37828 47908 37886
rect 47852 37762 47908 37772
rect 47964 37490 48020 38108
rect 48076 38052 48132 38062
rect 48076 37938 48132 37996
rect 48076 37886 48078 37938
rect 48130 37886 48132 37938
rect 48076 37874 48132 37886
rect 48188 37938 48244 38556
rect 48412 38500 48468 38510
rect 48412 38050 48468 38444
rect 48412 37998 48414 38050
rect 48466 37998 48468 38050
rect 48412 37986 48468 37998
rect 48748 38164 48804 38174
rect 48188 37886 48190 37938
rect 48242 37886 48244 37938
rect 48188 37874 48244 37886
rect 47964 37438 47966 37490
rect 48018 37438 48020 37490
rect 47964 37426 48020 37438
rect 48300 37826 48356 37838
rect 48300 37774 48302 37826
rect 48354 37774 48356 37826
rect 47740 37266 47796 37278
rect 47740 37214 47742 37266
rect 47794 37214 47796 37266
rect 47740 36708 47796 37214
rect 48188 37266 48244 37278
rect 48188 37214 48190 37266
rect 48242 37214 48244 37266
rect 48076 37154 48132 37166
rect 48076 37102 48078 37154
rect 48130 37102 48132 37154
rect 47852 36708 47908 36718
rect 47740 36652 47852 36708
rect 47852 36642 47908 36652
rect 47852 36484 47908 36494
rect 47628 36482 47908 36484
rect 47628 36430 47854 36482
rect 47906 36430 47908 36482
rect 47628 36428 47908 36430
rect 47852 36418 47908 36428
rect 48076 36370 48132 37102
rect 48188 36820 48244 37214
rect 48188 36754 48244 36764
rect 48188 36484 48244 36494
rect 48300 36484 48356 37774
rect 48412 37828 48468 37838
rect 48468 37772 48692 37828
rect 48412 37762 48468 37772
rect 48188 36482 48356 36484
rect 48188 36430 48190 36482
rect 48242 36430 48356 36482
rect 48188 36428 48356 36430
rect 48636 36484 48692 37772
rect 48748 37266 48804 38108
rect 48972 38050 49028 38062
rect 48972 37998 48974 38050
rect 49026 37998 49028 38050
rect 48972 37716 49028 37998
rect 49308 38052 49364 39790
rect 49420 39618 49476 39630
rect 49420 39566 49422 39618
rect 49474 39566 49476 39618
rect 49420 38724 49476 39566
rect 49420 38658 49476 38668
rect 49532 38836 49588 38846
rect 49532 38668 49588 38780
rect 49532 38612 49700 38668
rect 49308 37938 49364 37996
rect 49308 37886 49310 37938
rect 49362 37886 49364 37938
rect 49308 37874 49364 37886
rect 49532 37940 49588 37950
rect 48972 37650 49028 37660
rect 48860 37492 48916 37502
rect 48860 37398 48916 37436
rect 49420 37380 49476 37390
rect 49420 37286 49476 37324
rect 48748 37214 48750 37266
rect 48802 37214 48804 37266
rect 48748 37202 48804 37214
rect 49308 37266 49364 37278
rect 49308 37214 49310 37266
rect 49362 37214 49364 37266
rect 48748 37044 48804 37054
rect 48748 36706 48804 36988
rect 49308 37044 49364 37214
rect 49308 36978 49364 36988
rect 48748 36654 48750 36706
rect 48802 36654 48804 36706
rect 48748 36642 48804 36654
rect 49084 36708 49140 36718
rect 48748 36484 48804 36494
rect 48636 36482 48804 36484
rect 48636 36430 48750 36482
rect 48802 36430 48804 36482
rect 48636 36428 48804 36430
rect 48188 36418 48244 36428
rect 48076 36318 48078 36370
rect 48130 36318 48132 36370
rect 48076 36306 48132 36318
rect 48076 36148 48132 36158
rect 47628 35812 47684 35822
rect 47628 35718 47684 35756
rect 47852 35700 47908 35710
rect 47740 35588 47796 35598
rect 47740 35494 47796 35532
rect 47852 35364 47908 35644
rect 47740 35308 47908 35364
rect 48076 35308 48132 36092
rect 48748 35810 48804 36428
rect 49084 36370 49140 36652
rect 49084 36318 49086 36370
rect 49138 36318 49140 36370
rect 48748 35758 48750 35810
rect 48802 35758 48804 35810
rect 47740 34914 47796 35308
rect 47740 34862 47742 34914
rect 47794 34862 47796 34914
rect 47740 34354 47796 34862
rect 47740 34302 47742 34354
rect 47794 34302 47796 34354
rect 47740 34290 47796 34302
rect 47964 35252 48132 35308
rect 48188 35698 48244 35710
rect 48188 35646 48190 35698
rect 48242 35646 48244 35698
rect 47180 33404 47348 33460
rect 47404 33460 47460 33470
rect 47180 31948 47236 33404
rect 47404 33366 47460 33404
rect 47852 33124 47908 33134
rect 47852 33030 47908 33068
rect 47180 31892 47684 31948
rect 47180 31890 47236 31892
rect 47180 31838 47182 31890
rect 47234 31838 47236 31890
rect 47180 31826 47236 31838
rect 47068 31166 47070 31218
rect 47122 31166 47124 31218
rect 47068 31154 47124 31166
rect 47516 31778 47572 31790
rect 47516 31726 47518 31778
rect 47570 31726 47572 31778
rect 47404 30994 47460 31006
rect 47404 30942 47406 30994
rect 47458 30942 47460 30994
rect 46620 30370 46676 30380
rect 46732 30548 46788 30558
rect 46732 30212 46788 30492
rect 47404 30324 47460 30942
rect 47404 30258 47460 30268
rect 44716 29316 44772 29326
rect 44716 29222 44772 29260
rect 45052 29314 45108 29326
rect 45052 29262 45054 29314
rect 45106 29262 45108 29314
rect 45052 28868 45108 29262
rect 45836 29316 45892 29326
rect 45276 29204 45332 29214
rect 45276 29110 45332 29148
rect 45612 29202 45668 29214
rect 45612 29150 45614 29202
rect 45666 29150 45668 29202
rect 45052 28812 45332 28868
rect 45164 28642 45220 28654
rect 45164 28590 45166 28642
rect 45218 28590 45220 28642
rect 44828 28420 44884 28430
rect 44044 26002 44100 26012
rect 44156 26852 44436 26908
rect 44604 28418 44884 28420
rect 44604 28366 44830 28418
rect 44882 28366 44884 28418
rect 44604 28364 44884 28366
rect 43932 23314 43988 23324
rect 44156 22372 44212 26852
rect 44268 25508 44324 25518
rect 44268 25414 44324 25452
rect 44604 25172 44660 28364
rect 44828 28354 44884 28364
rect 45164 28308 45220 28590
rect 45164 28242 45220 28252
rect 45276 28644 45332 28812
rect 45388 28644 45444 28654
rect 45276 28642 45444 28644
rect 45276 28590 45390 28642
rect 45442 28590 45444 28642
rect 45276 28588 45444 28590
rect 44940 27300 44996 27310
rect 44716 27298 44996 27300
rect 44716 27246 44942 27298
rect 44994 27246 44996 27298
rect 44716 27244 44996 27246
rect 44716 26402 44772 27244
rect 44940 27234 44996 27244
rect 44828 26964 44884 27002
rect 44828 26898 44884 26908
rect 45052 26962 45108 26974
rect 45052 26910 45054 26962
rect 45106 26910 45108 26962
rect 44716 26350 44718 26402
rect 44770 26350 44772 26402
rect 44716 26338 44772 26350
rect 44828 26740 44884 26750
rect 44828 25730 44884 26684
rect 44828 25678 44830 25730
rect 44882 25678 44884 25730
rect 44828 25666 44884 25678
rect 45052 25732 45108 26910
rect 45276 26908 45332 28588
rect 45388 28578 45444 28588
rect 45612 27858 45668 29150
rect 45612 27806 45614 27858
rect 45666 27806 45668 27858
rect 45612 27794 45668 27806
rect 45724 28754 45780 28766
rect 45724 28702 45726 28754
rect 45778 28702 45780 28754
rect 45724 27636 45780 28702
rect 45836 28420 45892 29260
rect 45948 29202 46004 29214
rect 45948 29150 45950 29202
rect 46002 29150 46004 29202
rect 45948 28644 46004 29150
rect 45948 28578 46004 28588
rect 46060 28530 46116 28542
rect 46060 28478 46062 28530
rect 46114 28478 46116 28530
rect 45836 28418 46004 28420
rect 45836 28366 45838 28418
rect 45890 28366 46004 28418
rect 45836 28364 46004 28366
rect 45836 28354 45892 28364
rect 45948 28196 46004 28364
rect 45948 28130 46004 28140
rect 46060 27860 46116 28478
rect 46396 27860 46452 29932
rect 46620 30156 46788 30212
rect 46956 30212 47012 30222
rect 46508 29316 46564 29326
rect 46508 29222 46564 29260
rect 46060 27794 46116 27804
rect 46284 27804 46452 27860
rect 46508 28532 46564 28542
rect 46620 28532 46676 30156
rect 46956 29650 47012 30156
rect 46956 29598 46958 29650
rect 47010 29598 47012 29650
rect 46732 29204 46788 29214
rect 46732 28980 46788 29148
rect 46732 28642 46788 28924
rect 46956 28756 47012 29598
rect 47180 29988 47236 29998
rect 47516 29988 47572 31726
rect 47628 31220 47684 31892
rect 47628 31126 47684 31164
rect 47740 31108 47796 31118
rect 47964 31108 48020 35252
rect 48188 34914 48244 35646
rect 48188 34862 48190 34914
rect 48242 34862 48244 34914
rect 48188 34356 48244 34862
rect 48748 34916 48804 35758
rect 48860 35812 48916 35822
rect 48860 35810 49028 35812
rect 48860 35758 48862 35810
rect 48914 35758 49028 35810
rect 48860 35756 49028 35758
rect 48860 35746 48916 35756
rect 48860 35476 48916 35486
rect 48860 35382 48916 35420
rect 48748 34850 48804 34860
rect 48188 34290 48244 34300
rect 48748 34242 48804 34254
rect 48748 34190 48750 34242
rect 48802 34190 48804 34242
rect 48076 34018 48132 34030
rect 48076 33966 48078 34018
rect 48130 33966 48132 34018
rect 48076 33236 48132 33966
rect 48188 33908 48244 33918
rect 48188 33814 48244 33852
rect 48748 33460 48804 34190
rect 48972 33908 49028 35756
rect 49084 35138 49140 36318
rect 49420 36708 49476 36718
rect 49308 35698 49364 35710
rect 49308 35646 49310 35698
rect 49362 35646 49364 35698
rect 49308 35364 49364 35646
rect 49308 35298 49364 35308
rect 49420 35700 49476 36652
rect 49084 35086 49086 35138
rect 49138 35086 49140 35138
rect 49084 35074 49140 35086
rect 49196 35252 49252 35262
rect 49196 34914 49252 35196
rect 49196 34862 49198 34914
rect 49250 34862 49252 34914
rect 49196 34850 49252 34862
rect 49084 34244 49140 34254
rect 49084 34150 49140 34188
rect 48636 33404 48804 33460
rect 48860 33460 48916 33470
rect 48132 33180 48244 33236
rect 48076 33170 48132 33180
rect 48188 32450 48244 33180
rect 48636 33012 48692 33404
rect 48748 33236 48804 33246
rect 48748 33142 48804 33180
rect 48636 32956 48804 33012
rect 48188 32398 48190 32450
rect 48242 32398 48244 32450
rect 48188 32386 48244 32398
rect 48300 32340 48356 32350
rect 48188 31556 48244 31566
rect 47740 31106 48020 31108
rect 47740 31054 47742 31106
rect 47794 31054 48020 31106
rect 47740 31052 48020 31054
rect 48076 31500 48188 31556
rect 47740 31042 47796 31052
rect 47740 30884 47796 30894
rect 47740 30882 48020 30884
rect 47740 30830 47742 30882
rect 47794 30830 48020 30882
rect 47740 30828 48020 30830
rect 47740 30818 47796 30828
rect 47628 30212 47684 30222
rect 47628 30098 47684 30156
rect 47628 30046 47630 30098
rect 47682 30046 47684 30098
rect 47628 30034 47684 30046
rect 47180 29986 47572 29988
rect 47180 29934 47182 29986
rect 47234 29934 47572 29986
rect 47180 29932 47572 29934
rect 47180 29204 47236 29932
rect 47292 29428 47348 29438
rect 47292 29334 47348 29372
rect 47852 29428 47908 29438
rect 47852 29334 47908 29372
rect 47180 29138 47236 29148
rect 47068 28868 47124 28878
rect 47068 28866 47236 28868
rect 47068 28814 47070 28866
rect 47122 28814 47236 28866
rect 47068 28812 47236 28814
rect 47068 28802 47124 28812
rect 46956 28690 47012 28700
rect 46732 28590 46734 28642
rect 46786 28590 46788 28642
rect 46732 28578 46788 28590
rect 47068 28642 47124 28654
rect 47068 28590 47070 28642
rect 47122 28590 47124 28642
rect 46508 28530 46676 28532
rect 46508 28478 46510 28530
rect 46562 28478 46676 28530
rect 46508 28476 46676 28478
rect 46508 27860 46564 28476
rect 46732 27860 46788 27870
rect 46508 27804 46732 27860
rect 45388 27580 45780 27636
rect 45388 27298 45444 27580
rect 45388 27246 45390 27298
rect 45442 27246 45444 27298
rect 45388 27234 45444 27246
rect 45612 27300 45668 27310
rect 45612 27206 45668 27244
rect 46172 27076 46228 27114
rect 46172 27010 46228 27020
rect 46284 26908 46340 27804
rect 46732 27766 46788 27804
rect 46396 27636 46452 27646
rect 46396 27542 46452 27580
rect 45164 26852 45332 26908
rect 45948 26852 46340 26908
rect 46508 27524 46564 27534
rect 45164 26628 45220 26852
rect 45164 26562 45220 26572
rect 45052 25506 45108 25676
rect 45276 26292 45332 26302
rect 45164 25620 45220 25630
rect 45164 25526 45220 25564
rect 45052 25454 45054 25506
rect 45106 25454 45108 25506
rect 45052 25442 45108 25454
rect 44604 25106 44660 25116
rect 44940 25284 44996 25294
rect 44268 24724 44324 24734
rect 44268 23154 44324 24668
rect 44492 24722 44548 24734
rect 44492 24670 44494 24722
rect 44546 24670 44548 24722
rect 44380 24164 44436 24174
rect 44380 24070 44436 24108
rect 44268 23102 44270 23154
rect 44322 23102 44324 23154
rect 44268 23090 44324 23102
rect 43820 21606 43876 21644
rect 43932 22316 44212 22372
rect 43596 21588 43652 21598
rect 43596 21494 43652 21532
rect 43148 20290 43204 20300
rect 43260 20748 43428 20804
rect 43484 20804 43540 20814
rect 43036 20244 43092 20254
rect 42924 20242 43092 20244
rect 42924 20190 43038 20242
rect 43090 20190 43092 20242
rect 42924 20188 43092 20190
rect 43036 20178 43092 20188
rect 43036 19572 43092 19582
rect 43036 19234 43092 19516
rect 43036 19182 43038 19234
rect 43090 19182 43092 19234
rect 43036 19170 43092 19182
rect 42700 19122 42756 19134
rect 42700 19070 42702 19122
rect 42754 19070 42756 19122
rect 42700 18676 42756 19070
rect 42812 19012 42868 19022
rect 42812 19010 42980 19012
rect 42812 18958 42814 19010
rect 42866 18958 42980 19010
rect 42812 18956 42980 18958
rect 42812 18946 42868 18956
rect 42700 18610 42756 18620
rect 42812 18564 42868 18574
rect 42700 18452 42756 18462
rect 42700 18358 42756 18396
rect 42812 18450 42868 18508
rect 42812 18398 42814 18450
rect 42866 18398 42868 18450
rect 42812 18386 42868 18398
rect 42812 18116 42868 18126
rect 42924 18116 42980 18956
rect 43148 18450 43204 18462
rect 43148 18398 43150 18450
rect 43202 18398 43204 18450
rect 43036 18340 43092 18350
rect 43036 18246 43092 18284
rect 43148 18228 43204 18398
rect 43148 18162 43204 18172
rect 42868 18060 42980 18116
rect 42812 18050 42868 18060
rect 42812 17668 42868 17678
rect 42700 17666 42868 17668
rect 42700 17614 42814 17666
rect 42866 17614 42868 17666
rect 42700 17612 42868 17614
rect 42476 16706 42532 16716
rect 42588 17554 42644 17566
rect 42588 17502 42590 17554
rect 42642 17502 42644 17554
rect 42588 16882 42644 17502
rect 42588 16830 42590 16882
rect 42642 16830 42644 16882
rect 42364 16100 42420 16110
rect 42252 16098 42420 16100
rect 42252 16046 42366 16098
rect 42418 16046 42420 16098
rect 42252 16044 42420 16046
rect 42028 16034 42084 16044
rect 42364 16034 42420 16044
rect 42476 16100 42532 16110
rect 42140 15986 42196 15998
rect 42140 15934 42142 15986
rect 42194 15934 42196 15986
rect 41804 15708 41972 15764
rect 41804 15540 41860 15550
rect 41692 15428 41748 15466
rect 41804 15446 41860 15484
rect 41692 15362 41748 15372
rect 41692 15204 41748 15214
rect 41580 15202 41748 15204
rect 41580 15150 41694 15202
rect 41746 15150 41748 15202
rect 41580 15148 41748 15150
rect 41468 15138 41524 15148
rect 41692 15138 41748 15148
rect 41916 14980 41972 15708
rect 42028 15316 42084 15326
rect 42028 15222 42084 15260
rect 41916 14914 41972 14924
rect 42140 14756 42196 15934
rect 42140 14690 42196 14700
rect 42252 15204 42308 15214
rect 42476 15148 42532 16044
rect 42588 15540 42644 16830
rect 42588 15474 42644 15484
rect 42700 15316 42756 17612
rect 42812 17602 42868 17612
rect 43148 17442 43204 17454
rect 43148 17390 43150 17442
rect 43202 17390 43204 17442
rect 42924 16658 42980 16670
rect 42924 16606 42926 16658
rect 42978 16606 42980 16658
rect 42812 15988 42868 15998
rect 42812 15894 42868 15932
rect 42924 15428 42980 16606
rect 42924 15334 42980 15372
rect 43036 16098 43092 16110
rect 43036 16046 43038 16098
rect 43090 16046 43092 16098
rect 42812 15316 42868 15326
rect 42700 15260 42812 15316
rect 42812 15250 42868 15260
rect 42252 15092 42532 15148
rect 41244 14642 41412 14644
rect 41244 14590 41246 14642
rect 41298 14590 41412 14642
rect 41244 14588 41412 14590
rect 41244 14578 41300 14588
rect 41916 14532 41972 14542
rect 40908 14478 40910 14530
rect 40962 14478 40964 14530
rect 40908 14466 40964 14478
rect 41468 14530 41972 14532
rect 41468 14478 41918 14530
rect 41970 14478 41972 14530
rect 41468 14476 41972 14478
rect 41020 14420 41076 14430
rect 40796 14252 40964 14308
rect 40908 13748 40964 14252
rect 41020 13972 41076 14364
rect 41244 14418 41300 14430
rect 41244 14366 41246 14418
rect 41298 14366 41300 14418
rect 41132 14308 41188 14318
rect 41132 14214 41188 14252
rect 41132 13972 41188 13982
rect 41020 13970 41188 13972
rect 41020 13918 41134 13970
rect 41186 13918 41188 13970
rect 41020 13916 41188 13918
rect 41132 13906 41188 13916
rect 41020 13748 41076 13758
rect 40908 13746 41076 13748
rect 40908 13694 41022 13746
rect 41074 13694 41076 13746
rect 40908 13692 41076 13694
rect 41020 13682 41076 13692
rect 41132 13748 41188 13758
rect 40796 13636 40852 13646
rect 40796 13524 40852 13580
rect 40796 13468 41076 13524
rect 40684 13244 40964 13300
rect 40684 13076 40740 13086
rect 40684 12982 40740 13020
rect 40348 11342 40350 11394
rect 40402 11342 40404 11394
rect 40348 11330 40404 11342
rect 40460 11340 40628 11396
rect 40684 12852 40740 12862
rect 40348 10498 40404 10510
rect 40348 10446 40350 10498
rect 40402 10446 40404 10498
rect 40236 10388 40292 10398
rect 39900 9874 39956 9884
rect 40012 10386 40292 10388
rect 40012 10334 40238 10386
rect 40290 10334 40292 10386
rect 40012 10332 40292 10334
rect 39676 9604 39732 9614
rect 39676 9510 39732 9548
rect 39788 9602 39844 9614
rect 39788 9550 39790 9602
rect 39842 9550 39844 9602
rect 39564 9090 39620 9100
rect 39788 9044 39844 9550
rect 39340 8978 39396 8988
rect 39676 8988 39844 9044
rect 39900 9602 39956 9614
rect 39900 9550 39902 9602
rect 39954 9550 39956 9602
rect 39900 9044 39956 9550
rect 40012 9044 40068 10332
rect 40236 10322 40292 10332
rect 40348 10052 40404 10446
rect 40348 9986 40404 9996
rect 40124 9826 40180 9838
rect 40348 9828 40404 9838
rect 40124 9774 40126 9826
rect 40178 9774 40180 9826
rect 40124 9268 40180 9774
rect 40124 9202 40180 9212
rect 40236 9826 40404 9828
rect 40236 9774 40350 9826
rect 40402 9774 40404 9826
rect 40236 9772 40404 9774
rect 40124 9044 40180 9054
rect 40012 8988 40124 9044
rect 39564 8932 39620 8942
rect 39564 8838 39620 8876
rect 39228 8204 39508 8260
rect 39004 8082 39060 8092
rect 39116 8146 39172 8158
rect 39116 8094 39118 8146
rect 39170 8094 39172 8146
rect 39116 7924 39172 8094
rect 38892 7868 39172 7924
rect 39228 8036 39284 8046
rect 38780 7756 38948 7812
rect 38780 7474 38836 7486
rect 38780 7422 38782 7474
rect 38834 7422 38836 7474
rect 38780 5906 38836 7422
rect 38780 5854 38782 5906
rect 38834 5854 38836 5906
rect 38780 5348 38836 5854
rect 38780 5282 38836 5292
rect 38500 4844 38612 4900
rect 38668 4900 38724 4910
rect 38444 4834 38500 4844
rect 38332 3726 38334 3778
rect 38386 3726 38388 3778
rect 38332 3714 38388 3726
rect 38332 3556 38388 3566
rect 38332 3442 38388 3500
rect 38444 3556 38500 3566
rect 38668 3556 38724 4844
rect 38892 3668 38948 7756
rect 39228 7586 39284 7980
rect 39228 7534 39230 7586
rect 39282 7534 39284 7586
rect 39228 7522 39284 7534
rect 39340 7588 39396 7598
rect 39340 7494 39396 7532
rect 39340 7028 39396 7038
rect 39340 6804 39396 6972
rect 39340 6738 39396 6748
rect 39228 6580 39284 6590
rect 39452 6580 39508 8204
rect 39284 6524 39508 6580
rect 39564 7474 39620 7486
rect 39564 7422 39566 7474
rect 39618 7422 39620 7474
rect 39228 6486 39284 6524
rect 39564 6130 39620 7422
rect 39676 6804 39732 8988
rect 39900 8978 39956 8988
rect 40124 8950 40180 8988
rect 39788 8818 39844 8830
rect 39788 8766 39790 8818
rect 39842 8766 39844 8818
rect 39788 8146 39844 8766
rect 39900 8820 39956 8830
rect 39900 8370 39956 8764
rect 40236 8818 40292 9772
rect 40348 9762 40404 9772
rect 40348 9156 40404 9166
rect 40460 9156 40516 11340
rect 40684 11282 40740 12796
rect 40684 11230 40686 11282
rect 40738 11230 40740 11282
rect 40572 11170 40628 11182
rect 40572 11118 40574 11170
rect 40626 11118 40628 11170
rect 40572 10836 40628 11118
rect 40572 10770 40628 10780
rect 40684 9940 40740 11230
rect 40908 11060 40964 13244
rect 41020 12962 41076 13468
rect 41020 12910 41022 12962
rect 41074 12910 41076 12962
rect 41020 12898 41076 12910
rect 41132 11620 41188 13692
rect 41244 13636 41300 14366
rect 41356 14420 41412 14430
rect 41356 14326 41412 14364
rect 41356 13972 41412 13982
rect 41468 13972 41524 14476
rect 41916 14466 41972 14476
rect 41356 13970 41524 13972
rect 41356 13918 41358 13970
rect 41410 13918 41524 13970
rect 41356 13916 41524 13918
rect 41356 13906 41412 13916
rect 42140 13858 42196 13870
rect 42140 13806 42142 13858
rect 42194 13806 42196 13858
rect 41356 13636 41412 13646
rect 41244 13580 41356 13636
rect 41356 13570 41412 13580
rect 41916 13636 41972 13646
rect 42140 13636 42196 13806
rect 42252 13746 42308 15092
rect 42588 14532 42644 14542
rect 42364 14420 42420 14430
rect 42364 14418 42532 14420
rect 42364 14366 42366 14418
rect 42418 14366 42532 14418
rect 42364 14364 42532 14366
rect 42364 14354 42420 14364
rect 42252 13694 42254 13746
rect 42306 13694 42308 13746
rect 42252 13682 42308 13694
rect 41972 13580 42196 13636
rect 41916 13186 41972 13580
rect 41916 13134 41918 13186
rect 41970 13134 41972 13186
rect 41916 13122 41972 13134
rect 41468 12964 41524 12974
rect 41468 12870 41524 12908
rect 41468 12404 41524 12414
rect 41468 12310 41524 12348
rect 41244 12292 41300 12302
rect 41244 12198 41300 12236
rect 41692 12290 41748 12302
rect 41692 12238 41694 12290
rect 41746 12238 41748 12290
rect 41692 12180 41748 12238
rect 41916 12180 41972 12190
rect 41132 11554 41188 11564
rect 41580 12124 41692 12180
rect 41244 11396 41300 11406
rect 41244 11302 41300 11340
rect 41468 11284 41524 11294
rect 41580 11284 41636 12124
rect 41692 12114 41748 12124
rect 41804 12178 41972 12180
rect 41804 12126 41918 12178
rect 41970 12126 41972 12178
rect 41804 12124 41972 12126
rect 41804 12066 41860 12124
rect 41916 12114 41972 12124
rect 42028 12180 42084 12190
rect 41804 12014 41806 12066
rect 41858 12014 41860 12066
rect 41804 12002 41860 12014
rect 41468 11282 41636 11284
rect 41468 11230 41470 11282
rect 41522 11230 41636 11282
rect 41468 11228 41636 11230
rect 41804 11844 41860 11854
rect 41804 11394 41860 11788
rect 41804 11342 41806 11394
rect 41858 11342 41860 11394
rect 41468 11218 41524 11228
rect 40908 10994 40964 11004
rect 40684 9874 40740 9884
rect 41020 10780 41524 10836
rect 41020 10722 41076 10780
rect 41020 10670 41022 10722
rect 41074 10670 41076 10722
rect 41020 9714 41076 10670
rect 41356 10612 41412 10650
rect 41356 10546 41412 10556
rect 41468 10500 41524 10780
rect 41692 10724 41748 10734
rect 41804 10724 41860 11342
rect 42028 11394 42084 12124
rect 42476 12068 42532 14364
rect 42588 13524 42644 14476
rect 43036 14532 43092 16046
rect 43148 16098 43204 17390
rect 43260 17444 43316 20748
rect 43372 20580 43428 20590
rect 43484 20580 43540 20748
rect 43372 20578 43540 20580
rect 43372 20526 43374 20578
rect 43426 20526 43540 20578
rect 43372 20524 43540 20526
rect 43820 20580 43876 20590
rect 43372 20514 43428 20524
rect 43820 20486 43876 20524
rect 43932 19236 43988 22316
rect 44156 22148 44212 22158
rect 44156 22146 44324 22148
rect 44156 22094 44158 22146
rect 44210 22094 44324 22146
rect 44156 22092 44324 22094
rect 44156 22082 44212 22092
rect 44156 21698 44212 21710
rect 44156 21646 44158 21698
rect 44210 21646 44212 21698
rect 44156 21364 44212 21646
rect 44268 21588 44324 22092
rect 44492 21812 44548 24670
rect 44716 24610 44772 24622
rect 44716 24558 44718 24610
rect 44770 24558 44772 24610
rect 44604 23268 44660 23278
rect 44604 23174 44660 23212
rect 44716 22820 44772 24558
rect 44940 24050 44996 25228
rect 45052 24724 45108 24734
rect 45052 24630 45108 24668
rect 44940 23998 44942 24050
rect 44994 23998 44996 24050
rect 44940 23986 44996 23998
rect 45276 23828 45332 26236
rect 45612 26180 45668 26190
rect 45500 26068 45556 26078
rect 45388 25844 45444 25854
rect 45388 25730 45444 25788
rect 45388 25678 45390 25730
rect 45442 25678 45444 25730
rect 45388 25666 45444 25678
rect 45500 25284 45556 26012
rect 45612 25730 45668 26124
rect 45612 25678 45614 25730
rect 45666 25678 45668 25730
rect 45612 25666 45668 25678
rect 45836 26066 45892 26078
rect 45836 26014 45838 26066
rect 45890 26014 45892 26066
rect 45500 25218 45556 25228
rect 45164 23826 45332 23828
rect 45164 23774 45278 23826
rect 45330 23774 45332 23826
rect 45164 23772 45332 23774
rect 44716 22754 44772 22764
rect 44828 23714 44884 23726
rect 44828 23662 44830 23714
rect 44882 23662 44884 23714
rect 44828 22596 44884 23662
rect 45052 23714 45108 23726
rect 45052 23662 45054 23714
rect 45106 23662 45108 23714
rect 45052 23604 45108 23662
rect 45052 23538 45108 23548
rect 44940 23156 44996 23166
rect 44940 23062 44996 23100
rect 44828 22530 44884 22540
rect 44828 22372 44884 22382
rect 45164 22372 45220 23772
rect 45276 23762 45332 23772
rect 45388 24724 45444 24734
rect 45276 22484 45332 22494
rect 45276 22390 45332 22428
rect 44828 22278 44884 22316
rect 44940 22370 45220 22372
rect 44940 22318 45166 22370
rect 45218 22318 45220 22370
rect 44940 22316 45220 22318
rect 44940 22036 44996 22316
rect 45164 22306 45220 22316
rect 45388 22370 45444 24668
rect 45388 22318 45390 22370
rect 45442 22318 45444 22370
rect 45388 22306 45444 22318
rect 45500 24722 45556 24734
rect 45500 24670 45502 24722
rect 45554 24670 45556 24722
rect 44492 21718 44548 21756
rect 44604 21980 44996 22036
rect 44380 21588 44436 21598
rect 44268 21532 44380 21588
rect 44380 21522 44436 21532
rect 44604 21364 44660 21980
rect 45388 21812 45444 21822
rect 45500 21812 45556 24670
rect 45836 23716 45892 26014
rect 45948 24164 46004 26852
rect 46508 26516 46564 27468
rect 47068 27074 47124 28590
rect 47180 28084 47236 28812
rect 47964 28530 48020 30828
rect 48076 30660 48132 31500
rect 48188 31462 48244 31500
rect 48188 30996 48244 31006
rect 48188 30902 48244 30940
rect 48076 30594 48132 30604
rect 48076 29540 48132 29550
rect 48076 29446 48132 29484
rect 47964 28478 47966 28530
rect 48018 28478 48020 28530
rect 47964 28466 48020 28478
rect 47292 28420 47348 28430
rect 47292 28418 47460 28420
rect 47292 28366 47294 28418
rect 47346 28366 47460 28418
rect 47292 28364 47460 28366
rect 47292 28354 47348 28364
rect 47180 28018 47236 28028
rect 47292 28196 47348 28206
rect 47292 27860 47348 28140
rect 47068 27022 47070 27074
rect 47122 27022 47124 27074
rect 47068 26908 47124 27022
rect 46508 26450 46564 26460
rect 46956 26852 47124 26908
rect 47180 27858 47348 27860
rect 47180 27806 47294 27858
rect 47346 27806 47348 27858
rect 47180 27804 47348 27806
rect 46060 26404 46116 26414
rect 46060 25732 46116 26348
rect 46060 25638 46116 25676
rect 46172 26402 46228 26414
rect 46172 26350 46174 26402
rect 46226 26350 46228 26402
rect 46172 25396 46228 26350
rect 46620 26404 46676 26414
rect 46620 26402 46788 26404
rect 46620 26350 46622 26402
rect 46674 26350 46788 26402
rect 46620 26348 46788 26350
rect 46620 26338 46676 26348
rect 46620 26068 46676 26078
rect 46396 25844 46452 25854
rect 46172 25302 46228 25340
rect 46284 25788 46396 25844
rect 45948 24108 46228 24164
rect 45948 23940 46004 23950
rect 45948 23938 46116 23940
rect 45948 23886 45950 23938
rect 46002 23886 46116 23938
rect 45948 23884 46116 23886
rect 45948 23874 46004 23884
rect 45612 23660 45892 23716
rect 45948 23714 46004 23726
rect 45948 23662 45950 23714
rect 46002 23662 46004 23714
rect 45612 23268 45668 23660
rect 45612 23202 45668 23212
rect 45948 23268 46004 23662
rect 45388 21810 45556 21812
rect 45388 21758 45390 21810
rect 45442 21758 45556 21810
rect 45388 21756 45556 21758
rect 45724 23154 45780 23166
rect 45724 23102 45726 23154
rect 45778 23102 45780 23154
rect 45388 21746 45444 21756
rect 44716 21700 44772 21710
rect 44772 21644 44884 21700
rect 44716 21634 44772 21644
rect 44828 21586 44884 21644
rect 44828 21534 44830 21586
rect 44882 21534 44884 21586
rect 44828 21522 44884 21534
rect 45052 21588 45108 21598
rect 45052 21494 45108 21532
rect 45724 21588 45780 23102
rect 45948 23042 46004 23212
rect 45948 22990 45950 23042
rect 46002 22990 46004 23042
rect 45948 22978 46004 22990
rect 45836 22484 45892 22494
rect 45836 22390 45892 22428
rect 45836 21812 45892 21822
rect 45836 21718 45892 21756
rect 45724 21494 45780 21532
rect 46060 21476 46116 23884
rect 44156 21308 44660 21364
rect 45948 21420 46116 21476
rect 44156 21140 44212 21150
rect 44044 21084 44156 21140
rect 44044 19348 44100 21084
rect 44156 21074 44212 21084
rect 45948 20916 46004 21420
rect 45164 20804 45220 20814
rect 45164 20710 45220 20748
rect 45612 20804 45668 20814
rect 44156 20578 44212 20590
rect 44156 20526 44158 20578
rect 44210 20526 44212 20578
rect 44156 20468 44212 20526
rect 44156 20412 44660 20468
rect 44156 20244 44212 20254
rect 44156 20150 44212 20188
rect 44044 19292 44212 19348
rect 43820 19180 43988 19236
rect 43708 19122 43764 19134
rect 43708 19070 43710 19122
rect 43762 19070 43764 19122
rect 43596 18340 43652 18350
rect 43596 18246 43652 18284
rect 43708 18228 43764 19070
rect 43708 18162 43764 18172
rect 43820 17668 43876 19180
rect 44044 19122 44100 19134
rect 44044 19070 44046 19122
rect 44098 19070 44100 19122
rect 43932 19012 43988 19022
rect 43932 18918 43988 18956
rect 44044 18900 44100 19070
rect 44156 19012 44212 19292
rect 44268 19236 44324 19246
rect 44604 19236 44660 20412
rect 45500 20020 45556 20030
rect 45500 19926 45556 19964
rect 45612 19908 45668 20748
rect 45948 20130 46004 20860
rect 45948 20078 45950 20130
rect 46002 20078 46004 20130
rect 45948 20066 46004 20078
rect 45052 19458 45108 19470
rect 45052 19406 45054 19458
rect 45106 19406 45108 19458
rect 44828 19236 44884 19246
rect 44268 19234 44436 19236
rect 44268 19182 44270 19234
rect 44322 19182 44436 19234
rect 44268 19180 44436 19182
rect 44604 19234 44884 19236
rect 44604 19182 44830 19234
rect 44882 19182 44884 19234
rect 44604 19180 44884 19182
rect 44268 19170 44324 19180
rect 44156 18956 44324 19012
rect 44044 18844 44212 18900
rect 44044 18676 44100 18686
rect 44044 18450 44100 18620
rect 44156 18564 44212 18844
rect 44156 18498 44212 18508
rect 44044 18398 44046 18450
rect 44098 18398 44100 18450
rect 44044 18386 44100 18398
rect 44268 18004 44324 18956
rect 44380 18452 44436 19180
rect 44828 18452 44884 19180
rect 44940 18900 44996 18910
rect 44940 18562 44996 18844
rect 44940 18510 44942 18562
rect 44994 18510 44996 18562
rect 44940 18498 44996 18510
rect 44380 18396 44772 18452
rect 44380 18228 44436 18238
rect 44380 18226 44660 18228
rect 44380 18174 44382 18226
rect 44434 18174 44660 18226
rect 44380 18172 44660 18174
rect 44380 18162 44436 18172
rect 44268 17948 44436 18004
rect 43820 17666 44324 17668
rect 43820 17614 43822 17666
rect 43874 17614 44324 17666
rect 43820 17612 44324 17614
rect 43820 17602 43876 17612
rect 43708 17556 43764 17566
rect 43708 17462 43764 17500
rect 43260 16994 43316 17388
rect 43596 17442 43652 17454
rect 43596 17390 43598 17442
rect 43650 17390 43652 17442
rect 43596 17332 43652 17390
rect 43596 17266 43652 17276
rect 43260 16942 43262 16994
rect 43314 16942 43316 16994
rect 43260 16930 43316 16942
rect 43148 16046 43150 16098
rect 43202 16046 43204 16098
rect 43148 15876 43204 16046
rect 43596 16660 43652 16670
rect 43596 15876 43652 16604
rect 43148 15820 43428 15876
rect 43036 14466 43092 14476
rect 43148 15316 43204 15326
rect 42588 13458 42644 13468
rect 42700 14308 42756 14318
rect 42700 13748 42756 14252
rect 42700 12962 42756 13692
rect 43036 13636 43092 13646
rect 42700 12910 42702 12962
rect 42754 12910 42756 12962
rect 42700 12898 42756 12910
rect 42812 13524 42868 13534
rect 42812 12292 42868 13468
rect 42700 12180 42756 12190
rect 42700 12086 42756 12124
rect 42588 12068 42644 12078
rect 42476 12066 42644 12068
rect 42476 12014 42590 12066
rect 42642 12014 42644 12066
rect 42476 12012 42644 12014
rect 42476 11844 42532 12012
rect 42588 12002 42644 12012
rect 42476 11778 42532 11788
rect 42812 11732 42868 12236
rect 43036 12404 43092 13580
rect 42812 11676 42980 11732
rect 42812 11508 42868 11518
rect 42028 11342 42030 11394
rect 42082 11342 42084 11394
rect 41692 10722 41860 10724
rect 41692 10670 41694 10722
rect 41746 10670 41860 10722
rect 41692 10668 41860 10670
rect 41916 11170 41972 11182
rect 41916 11118 41918 11170
rect 41970 11118 41972 11170
rect 41692 10658 41748 10668
rect 41916 10612 41972 11118
rect 41804 10556 41972 10612
rect 42028 10610 42084 11342
rect 42364 11506 42868 11508
rect 42364 11454 42814 11506
rect 42866 11454 42868 11506
rect 42364 11452 42868 11454
rect 42364 11394 42420 11452
rect 42812 11442 42868 11452
rect 42364 11342 42366 11394
rect 42418 11342 42420 11394
rect 42028 10558 42030 10610
rect 42082 10558 42084 10610
rect 41804 10500 41860 10556
rect 42028 10546 42084 10558
rect 42140 10612 42196 10622
rect 42252 10612 42308 10622
rect 42196 10610 42308 10612
rect 42196 10558 42254 10610
rect 42306 10558 42308 10610
rect 42196 10556 42308 10558
rect 41468 10444 41860 10500
rect 41356 10388 41412 10398
rect 41356 10386 41748 10388
rect 41356 10334 41358 10386
rect 41410 10334 41748 10386
rect 41356 10332 41748 10334
rect 41356 10322 41412 10332
rect 41580 9828 41636 9838
rect 41580 9734 41636 9772
rect 41020 9662 41022 9714
rect 41074 9662 41076 9714
rect 41020 9650 41076 9662
rect 41356 9716 41412 9726
rect 41356 9622 41412 9660
rect 40348 9154 40516 9156
rect 40348 9102 40350 9154
rect 40402 9102 40516 9154
rect 40348 9100 40516 9102
rect 41468 9604 41524 9614
rect 40348 9090 40404 9100
rect 41020 9044 41076 9054
rect 40236 8766 40238 8818
rect 40290 8766 40292 8818
rect 40236 8754 40292 8766
rect 40796 8988 41020 9044
rect 39900 8318 39902 8370
rect 39954 8318 39956 8370
rect 39900 8306 39956 8318
rect 40012 8596 40068 8606
rect 39788 8094 39790 8146
rect 39842 8094 39844 8146
rect 39788 7476 39844 8094
rect 39788 7410 39844 7420
rect 39788 7252 39844 7262
rect 39788 7158 39844 7196
rect 40012 6916 40068 8540
rect 40236 8258 40292 8270
rect 40236 8206 40238 8258
rect 40290 8206 40292 8258
rect 40124 7252 40180 7262
rect 40124 7158 40180 7196
rect 39676 6738 39732 6748
rect 39788 6860 40068 6916
rect 39564 6078 39566 6130
rect 39618 6078 39620 6130
rect 39564 6066 39620 6078
rect 39788 6132 39844 6860
rect 40236 6692 40292 8206
rect 40796 7474 40852 8988
rect 41020 8950 41076 8988
rect 41468 9042 41524 9548
rect 41468 8990 41470 9042
rect 41522 8990 41524 9042
rect 41468 8978 41524 8990
rect 41692 9042 41748 10332
rect 41916 9602 41972 9614
rect 41916 9550 41918 9602
rect 41970 9550 41972 9602
rect 41692 8990 41694 9042
rect 41746 8990 41748 9042
rect 41692 8978 41748 8990
rect 41804 9266 41860 9278
rect 41804 9214 41806 9266
rect 41858 9214 41860 9266
rect 41580 8932 41636 8942
rect 40908 8820 40964 8830
rect 40908 8818 41300 8820
rect 40908 8766 40910 8818
rect 40962 8766 41300 8818
rect 40908 8764 41300 8766
rect 40908 8754 40964 8764
rect 40796 7422 40798 7474
rect 40850 7422 40852 7474
rect 40796 7410 40852 7422
rect 41020 8146 41076 8158
rect 41020 8094 41022 8146
rect 41074 8094 41076 8146
rect 40236 6626 40292 6636
rect 40348 7362 40404 7374
rect 40348 7310 40350 7362
rect 40402 7310 40404 7362
rect 39788 6038 39844 6076
rect 40012 6468 40068 6478
rect 40348 6468 40404 7310
rect 41020 7252 41076 8094
rect 41244 7700 41300 8764
rect 41356 8036 41412 8046
rect 41356 7942 41412 7980
rect 41356 7700 41412 7710
rect 41244 7698 41412 7700
rect 41244 7646 41358 7698
rect 41410 7646 41412 7698
rect 41244 7644 41412 7646
rect 41356 7634 41412 7644
rect 41468 7700 41524 7710
rect 41580 7700 41636 8876
rect 41468 7698 41636 7700
rect 41468 7646 41470 7698
rect 41522 7646 41636 7698
rect 41468 7644 41636 7646
rect 41468 7634 41524 7644
rect 41804 7588 41860 9214
rect 41692 7532 41860 7588
rect 41916 7588 41972 9550
rect 41244 7476 41300 7486
rect 41244 7382 41300 7420
rect 40012 6466 40404 6468
rect 40012 6414 40014 6466
rect 40066 6414 40404 6466
rect 40012 6412 40404 6414
rect 40460 6804 40516 6814
rect 40012 5908 40068 6412
rect 40012 5842 40068 5852
rect 40124 5906 40180 5918
rect 40124 5854 40126 5906
rect 40178 5854 40180 5906
rect 39676 5796 39732 5806
rect 39116 5794 39732 5796
rect 39116 5742 39678 5794
rect 39730 5742 39732 5794
rect 39116 5740 39732 5742
rect 39116 5234 39172 5740
rect 39676 5730 39732 5740
rect 39116 5182 39118 5234
rect 39170 5182 39172 5234
rect 39116 5170 39172 5182
rect 39900 5122 39956 5134
rect 39900 5070 39902 5122
rect 39954 5070 39956 5122
rect 39900 3780 39956 5070
rect 40124 5124 40180 5854
rect 40124 5058 40180 5068
rect 40236 5572 40292 5582
rect 40236 4452 40292 5516
rect 40236 4338 40292 4396
rect 40236 4286 40238 4338
rect 40290 4286 40292 4338
rect 40236 4274 40292 4286
rect 39004 3668 39060 3678
rect 38892 3666 39060 3668
rect 38892 3614 39006 3666
rect 39058 3614 39060 3666
rect 38892 3612 39060 3614
rect 39004 3602 39060 3612
rect 38444 3554 38668 3556
rect 38444 3502 38446 3554
rect 38498 3502 38668 3554
rect 38444 3500 38668 3502
rect 38444 3490 38500 3500
rect 38668 3462 38724 3500
rect 39900 3554 39956 3724
rect 40460 3668 40516 6748
rect 40572 6692 40628 6702
rect 40572 6356 40628 6636
rect 40572 5346 40628 6300
rect 40572 5294 40574 5346
rect 40626 5294 40628 5346
rect 40572 5282 40628 5294
rect 41020 6580 41076 7196
rect 41692 6580 41748 7532
rect 41916 7522 41972 7532
rect 42028 8146 42084 8158
rect 42028 8094 42030 8146
rect 42082 8094 42084 8146
rect 41916 7364 41972 7374
rect 41916 7270 41972 7308
rect 41804 6580 41860 6590
rect 41692 6578 41860 6580
rect 41692 6526 41806 6578
rect 41858 6526 41860 6578
rect 41692 6524 41860 6526
rect 41020 4562 41076 6524
rect 41804 6514 41860 6524
rect 41580 6018 41636 6030
rect 41580 5966 41582 6018
rect 41634 5966 41636 6018
rect 41020 4510 41022 4562
rect 41074 4510 41076 4562
rect 41020 4498 41076 4510
rect 41356 5906 41412 5918
rect 41356 5854 41358 5906
rect 41410 5854 41412 5906
rect 41356 4340 41412 5854
rect 41580 5124 41636 5966
rect 41916 5908 41972 5918
rect 41916 5814 41972 5852
rect 42028 5236 42084 8094
rect 42140 8036 42196 10556
rect 42252 10546 42308 10556
rect 42252 10388 42308 10398
rect 42364 10388 42420 11342
rect 42700 11284 42756 11294
rect 42924 11284 42980 11676
rect 43036 11394 43092 12348
rect 43036 11342 43038 11394
rect 43090 11342 43092 11394
rect 43036 11330 43092 11342
rect 42700 11282 42980 11284
rect 42700 11230 42702 11282
rect 42754 11230 42980 11282
rect 42700 11228 42980 11230
rect 42700 11218 42756 11228
rect 43148 11060 43204 15260
rect 43372 14642 43428 15820
rect 43372 14590 43374 14642
rect 43426 14590 43428 14642
rect 43372 14578 43428 14590
rect 43484 15820 43652 15876
rect 43260 14532 43316 14542
rect 43260 13746 43316 14476
rect 43260 13694 43262 13746
rect 43314 13694 43316 13746
rect 43260 13682 43316 13694
rect 43484 13524 43540 15820
rect 43260 13468 43540 13524
rect 43596 15314 43652 15326
rect 43596 15262 43598 15314
rect 43650 15262 43652 15314
rect 43596 14420 43652 15262
rect 43708 14756 43764 14766
rect 43764 14700 43876 14756
rect 43708 14690 43764 14700
rect 43708 14420 43764 14430
rect 43652 14418 43764 14420
rect 43652 14366 43710 14418
rect 43762 14366 43764 14418
rect 43652 14364 43764 14366
rect 43260 12964 43316 13468
rect 43372 13076 43428 13086
rect 43596 13076 43652 14364
rect 43708 14354 43764 14364
rect 43708 13748 43764 13758
rect 43708 13654 43764 13692
rect 43372 13074 43652 13076
rect 43372 13022 43374 13074
rect 43426 13022 43652 13074
rect 43372 13020 43652 13022
rect 43372 13010 43428 13020
rect 43260 12898 43316 12908
rect 43820 12962 43876 14700
rect 43820 12910 43822 12962
rect 43874 12910 43876 12962
rect 43820 12898 43876 12910
rect 43372 12292 43428 12302
rect 43372 12198 43428 12236
rect 43260 12180 43316 12190
rect 43260 11396 43316 12124
rect 43260 11302 43316 11340
rect 43036 11004 43204 11060
rect 42476 10836 42532 10846
rect 42476 10834 42868 10836
rect 42476 10782 42478 10834
rect 42530 10782 42868 10834
rect 42476 10780 42868 10782
rect 42476 10770 42532 10780
rect 42252 10386 42420 10388
rect 42252 10334 42254 10386
rect 42306 10334 42420 10386
rect 42252 10332 42420 10334
rect 42252 10322 42308 10332
rect 42252 10052 42308 10062
rect 42252 9044 42308 9996
rect 42700 9828 42756 9838
rect 42700 9734 42756 9772
rect 42476 9716 42532 9726
rect 42476 9602 42532 9660
rect 42476 9550 42478 9602
rect 42530 9550 42532 9602
rect 42364 9268 42420 9306
rect 42364 9202 42420 9212
rect 42364 9044 42420 9054
rect 42252 8988 42364 9044
rect 42364 8950 42420 8988
rect 42476 8484 42532 9550
rect 42588 9604 42644 9614
rect 42588 9510 42644 9548
rect 42700 9044 42756 9054
rect 42812 9044 42868 10780
rect 42700 9042 42868 9044
rect 42700 8990 42702 9042
rect 42754 8990 42868 9042
rect 42700 8988 42868 8990
rect 42924 9042 42980 9054
rect 42924 8990 42926 9042
rect 42978 8990 42980 9042
rect 42700 8978 42756 8988
rect 42476 8428 42756 8484
rect 42140 5906 42196 7980
rect 42364 8258 42420 8270
rect 42364 8206 42366 8258
rect 42418 8206 42420 8258
rect 42364 7700 42420 8206
rect 42364 7698 42644 7700
rect 42364 7646 42366 7698
rect 42418 7646 42644 7698
rect 42364 7644 42644 7646
rect 42364 7634 42420 7644
rect 42476 6916 42532 6926
rect 42476 6130 42532 6860
rect 42588 6914 42644 7644
rect 42700 7364 42756 8428
rect 42812 8036 42868 8046
rect 42924 8036 42980 8990
rect 43036 8372 43092 11004
rect 43484 10948 43540 10958
rect 43260 9940 43316 9950
rect 43148 9828 43204 9838
rect 43148 9154 43204 9772
rect 43148 9102 43150 9154
rect 43202 9102 43204 9154
rect 43148 8596 43204 9102
rect 43148 8530 43204 8540
rect 43148 8372 43204 8382
rect 43036 8370 43204 8372
rect 43036 8318 43150 8370
rect 43202 8318 43204 8370
rect 43036 8316 43204 8318
rect 43148 8306 43204 8316
rect 43260 8148 43316 9884
rect 43484 9714 43540 10892
rect 43596 10836 43652 10846
rect 43596 10722 43652 10780
rect 43596 10670 43598 10722
rect 43650 10670 43652 10722
rect 43596 10658 43652 10670
rect 43596 10052 43652 10062
rect 43596 9826 43652 9996
rect 43596 9774 43598 9826
rect 43650 9774 43652 9826
rect 43596 9762 43652 9774
rect 43484 9662 43486 9714
rect 43538 9662 43540 9714
rect 43484 9650 43540 9662
rect 43596 9268 43652 9278
rect 43596 9174 43652 9212
rect 43820 9044 43876 9054
rect 43708 8708 43764 8718
rect 42868 7980 42980 8036
rect 43148 8092 43316 8148
rect 43596 8258 43652 8270
rect 43596 8206 43598 8258
rect 43650 8206 43652 8258
rect 42812 7970 42868 7980
rect 42924 7588 42980 7598
rect 42924 7474 42980 7532
rect 42924 7422 42926 7474
rect 42978 7422 42980 7474
rect 42924 7410 42980 7422
rect 42700 7298 42756 7308
rect 42588 6862 42590 6914
rect 42642 6862 42644 6914
rect 42588 6850 42644 6862
rect 42700 6580 42756 6590
rect 42700 6486 42756 6524
rect 42476 6078 42478 6130
rect 42530 6078 42532 6130
rect 42476 6066 42532 6078
rect 42140 5854 42142 5906
rect 42194 5854 42196 5906
rect 42140 5842 42196 5854
rect 42252 5236 42308 5246
rect 42028 5180 42252 5236
rect 42252 5170 42308 5180
rect 43036 5236 43092 5246
rect 43036 5142 43092 5180
rect 41580 5068 42084 5124
rect 42028 5012 42084 5068
rect 42084 4956 42196 5012
rect 42028 4918 42084 4956
rect 42140 4562 42196 4956
rect 42140 4510 42142 4562
rect 42194 4510 42196 4562
rect 42140 4498 42196 4510
rect 41356 4274 41412 4284
rect 42700 4340 42756 4350
rect 40572 3668 40628 3678
rect 40460 3666 40628 3668
rect 40460 3614 40574 3666
rect 40626 3614 40628 3666
rect 40460 3612 40628 3614
rect 40572 3602 40628 3612
rect 42700 3668 42756 4284
rect 43148 4340 43204 8092
rect 43372 7588 43428 7598
rect 43372 7494 43428 7532
rect 43484 7586 43540 7598
rect 43484 7534 43486 7586
rect 43538 7534 43540 7586
rect 43484 7476 43540 7534
rect 43484 7410 43540 7420
rect 43372 7362 43428 7374
rect 43372 7310 43374 7362
rect 43426 7310 43428 7362
rect 43260 6692 43316 6702
rect 43260 6598 43316 6636
rect 43260 6468 43316 6478
rect 43260 6374 43316 6412
rect 43260 6020 43316 6030
rect 43372 6020 43428 7310
rect 43596 6916 43652 8206
rect 43708 7698 43764 8652
rect 43708 7646 43710 7698
rect 43762 7646 43764 7698
rect 43708 7634 43764 7646
rect 43596 6850 43652 6860
rect 43260 6018 43428 6020
rect 43260 5966 43262 6018
rect 43314 5966 43428 6018
rect 43260 5964 43428 5966
rect 43708 6132 43764 6142
rect 43260 5954 43316 5964
rect 43372 5122 43428 5134
rect 43372 5070 43374 5122
rect 43426 5070 43428 5122
rect 43372 5012 43428 5070
rect 43372 4946 43428 4956
rect 43148 4274 43204 4284
rect 43708 3668 43764 6076
rect 43820 5122 43876 8988
rect 43932 8708 43988 17612
rect 44044 17444 44100 17454
rect 44044 17350 44100 17388
rect 44268 16882 44324 17612
rect 44268 16830 44270 16882
rect 44322 16830 44324 16882
rect 44268 16818 44324 16830
rect 44268 16100 44324 16110
rect 44268 16006 44324 16044
rect 44268 15540 44324 15550
rect 44044 15316 44100 15326
rect 44044 15222 44100 15260
rect 44268 15314 44324 15484
rect 44268 15262 44270 15314
rect 44322 15262 44324 15314
rect 44268 15148 44324 15262
rect 44156 15092 44324 15148
rect 44156 12402 44212 15092
rect 44268 14644 44324 14654
rect 44380 14644 44436 17948
rect 44604 15148 44660 18172
rect 44716 17892 44772 18396
rect 44828 18340 44884 18396
rect 44828 18284 44996 18340
rect 44828 17892 44884 17902
rect 44716 17890 44884 17892
rect 44716 17838 44830 17890
rect 44882 17838 44884 17890
rect 44716 17836 44884 17838
rect 44828 16098 44884 17836
rect 44940 17778 44996 18284
rect 44940 17726 44942 17778
rect 44994 17726 44996 17778
rect 44940 17714 44996 17726
rect 44828 16046 44830 16098
rect 44882 16046 44884 16098
rect 44828 16034 44884 16046
rect 45052 16322 45108 19406
rect 45612 19348 45668 19852
rect 46172 19684 46228 24108
rect 46284 23378 46340 25788
rect 46396 25778 46452 25788
rect 46620 25620 46676 26012
rect 46508 25618 46676 25620
rect 46508 25566 46622 25618
rect 46674 25566 46676 25618
rect 46508 25564 46676 25566
rect 46396 24724 46452 24734
rect 46396 24630 46452 24668
rect 46508 23380 46564 25564
rect 46620 25554 46676 25564
rect 46620 25284 46676 25294
rect 46620 23716 46676 25228
rect 46732 24498 46788 26348
rect 46956 25396 47012 26852
rect 47180 26740 47236 27804
rect 47292 27794 47348 27804
rect 47068 26684 47236 26740
rect 47292 27076 47348 27086
rect 47068 26516 47124 26684
rect 47292 26628 47348 27020
rect 47068 26450 47124 26460
rect 47180 26572 47348 26628
rect 47068 26066 47124 26078
rect 47068 26014 47070 26066
rect 47122 26014 47124 26066
rect 47068 25620 47124 26014
rect 47068 25554 47124 25564
rect 47068 25396 47124 25406
rect 46956 25340 47068 25396
rect 47068 24834 47124 25340
rect 47068 24782 47070 24834
rect 47122 24782 47124 24834
rect 47068 24770 47124 24782
rect 47180 24836 47236 26572
rect 47404 26516 47460 28364
rect 48300 28196 48356 32284
rect 48748 31892 48804 32956
rect 48860 32674 48916 33404
rect 48972 32786 49028 33852
rect 49308 33236 49364 33246
rect 48972 32734 48974 32786
rect 49026 32734 49028 32786
rect 48972 32722 49028 32734
rect 49196 32788 49252 32798
rect 49196 32694 49252 32732
rect 48860 32622 48862 32674
rect 48914 32622 48916 32674
rect 48860 32610 48916 32622
rect 48748 31826 48804 31836
rect 49308 31666 49364 33180
rect 49308 31614 49310 31666
rect 49362 31614 49364 31666
rect 49308 31106 49364 31614
rect 49308 31054 49310 31106
rect 49362 31054 49364 31106
rect 49308 31042 49364 31054
rect 49420 30884 49476 35644
rect 49532 32676 49588 37884
rect 49532 32610 49588 32620
rect 49532 32450 49588 32462
rect 49532 32398 49534 32450
rect 49586 32398 49588 32450
rect 49532 32338 49588 32398
rect 49532 32286 49534 32338
rect 49586 32286 49588 32338
rect 49532 32274 49588 32286
rect 49196 30828 49476 30884
rect 48300 28130 48356 28140
rect 48636 30210 48692 30222
rect 48636 30158 48638 30210
rect 48690 30158 48692 30210
rect 48636 29092 48692 30158
rect 48860 29428 48916 29438
rect 48748 29316 48804 29326
rect 48748 29222 48804 29260
rect 47516 27972 47572 27982
rect 47516 27878 47572 27916
rect 48076 27746 48132 27758
rect 48076 27694 48078 27746
rect 48130 27694 48132 27746
rect 48076 26908 48132 27694
rect 47292 26460 47460 26516
rect 47964 26852 48132 26908
rect 47292 26290 47348 26460
rect 47292 26238 47294 26290
rect 47346 26238 47348 26290
rect 47292 26226 47348 26238
rect 47516 26290 47572 26302
rect 47516 26238 47518 26290
rect 47570 26238 47572 26290
rect 47516 25060 47572 26238
rect 47740 26290 47796 26302
rect 47740 26238 47742 26290
rect 47794 26238 47796 26290
rect 47628 26180 47684 26190
rect 47628 26086 47684 26124
rect 47740 25956 47796 26238
rect 47740 25890 47796 25900
rect 47964 25508 48020 26852
rect 47516 25004 47908 25060
rect 47292 24836 47348 24846
rect 47628 24836 47684 24846
rect 47180 24834 47348 24836
rect 47180 24782 47294 24834
rect 47346 24782 47348 24834
rect 47180 24780 47348 24782
rect 47292 24770 47348 24780
rect 47516 24780 47628 24836
rect 46732 24446 46734 24498
rect 46786 24446 46788 24498
rect 46732 24164 46788 24446
rect 46732 24098 46788 24108
rect 46732 23940 46788 23950
rect 47516 23940 47572 24780
rect 47628 24770 47684 24780
rect 46732 23846 46788 23884
rect 47404 23938 47572 23940
rect 47404 23886 47518 23938
rect 47570 23886 47572 23938
rect 47404 23884 47572 23886
rect 46844 23826 46900 23838
rect 46844 23774 46846 23826
rect 46898 23774 46900 23826
rect 46844 23716 46900 23774
rect 46620 23660 46788 23716
rect 46284 23326 46286 23378
rect 46338 23326 46340 23378
rect 46284 23314 46340 23326
rect 46396 23324 46564 23380
rect 46620 23492 46676 23502
rect 46396 23156 46452 23324
rect 46620 23268 46676 23436
rect 46396 23090 46452 23100
rect 46508 23266 46676 23268
rect 46508 23214 46622 23266
rect 46674 23214 46676 23266
rect 46508 23212 46676 23214
rect 46508 22932 46564 23212
rect 46620 23202 46676 23212
rect 46396 22876 46564 22932
rect 45612 19282 45668 19292
rect 45724 19628 46228 19684
rect 46284 20802 46340 20814
rect 46284 20750 46286 20802
rect 46338 20750 46340 20802
rect 45388 19122 45444 19134
rect 45388 19070 45390 19122
rect 45442 19070 45444 19122
rect 45164 18452 45220 18462
rect 45388 18452 45444 19070
rect 45500 19124 45556 19134
rect 45500 19030 45556 19068
rect 45612 19122 45668 19134
rect 45612 19070 45614 19122
rect 45666 19070 45668 19122
rect 45164 18450 45388 18452
rect 45164 18398 45166 18450
rect 45218 18398 45388 18450
rect 45164 18396 45388 18398
rect 45164 17556 45220 18396
rect 45388 18358 45444 18396
rect 45612 18900 45668 19070
rect 45500 18340 45556 18350
rect 45276 17892 45332 17902
rect 45276 17798 45332 17836
rect 45164 17500 45444 17556
rect 45052 16270 45054 16322
rect 45106 16270 45108 16322
rect 44828 15876 44884 15886
rect 44828 15782 44884 15820
rect 44604 15092 44884 15148
rect 44268 14642 44436 14644
rect 44268 14590 44270 14642
rect 44322 14590 44436 14642
rect 44268 14588 44436 14590
rect 44268 14578 44324 14588
rect 44492 13524 44548 13534
rect 44492 13430 44548 13468
rect 44268 12852 44324 12862
rect 44268 12758 44324 12796
rect 44156 12350 44158 12402
rect 44210 12350 44212 12402
rect 44156 12338 44212 12350
rect 44716 12290 44772 12302
rect 44716 12238 44718 12290
rect 44770 12238 44772 12290
rect 44268 12180 44324 12190
rect 44268 12086 44324 12124
rect 44156 11394 44212 11406
rect 44156 11342 44158 11394
rect 44210 11342 44212 11394
rect 44156 11284 44212 11342
rect 44156 11218 44212 11228
rect 44716 11284 44772 12238
rect 44828 11508 44884 15092
rect 44940 14756 44996 14766
rect 44940 14662 44996 14700
rect 44940 12852 44996 12862
rect 44940 12758 44996 12796
rect 45052 12402 45108 16270
rect 45388 15986 45444 17500
rect 45388 15934 45390 15986
rect 45442 15934 45444 15986
rect 45388 15148 45444 15934
rect 45500 15540 45556 18284
rect 45612 16098 45668 18844
rect 45724 17780 45780 19628
rect 46060 19348 46116 19358
rect 45948 19234 46004 19246
rect 45948 19182 45950 19234
rect 46002 19182 46004 19234
rect 45948 18452 46004 19182
rect 46060 18562 46116 19292
rect 46060 18510 46062 18562
rect 46114 18510 46116 18562
rect 46060 18498 46116 18510
rect 46172 19236 46228 19246
rect 45948 18386 46004 18396
rect 45724 17332 45780 17724
rect 45724 16882 45780 17276
rect 45724 16830 45726 16882
rect 45778 16830 45780 16882
rect 45724 16818 45780 16830
rect 45836 18116 45892 18126
rect 45836 16996 45892 18060
rect 46172 17106 46228 19180
rect 46284 18452 46340 20750
rect 46396 19906 46452 22876
rect 46620 22372 46676 22382
rect 46620 21810 46676 22316
rect 46620 21758 46622 21810
rect 46674 21758 46676 21810
rect 46620 21746 46676 21758
rect 46732 20020 46788 23660
rect 46844 23650 46900 23660
rect 47404 23492 47460 23884
rect 47516 23874 47572 23884
rect 47180 23268 47236 23278
rect 47180 23174 47236 23212
rect 47404 23266 47460 23436
rect 47628 23826 47684 23838
rect 47628 23774 47630 23826
rect 47682 23774 47684 23826
rect 47516 23380 47572 23390
rect 47516 23286 47572 23324
rect 47404 23214 47406 23266
rect 47458 23214 47460 23266
rect 47404 23202 47460 23214
rect 46844 23156 46900 23166
rect 46844 23062 46900 23100
rect 47068 22820 47124 22830
rect 47068 22260 47124 22764
rect 47628 22596 47684 23774
rect 46956 21588 47012 21598
rect 47068 21588 47124 22204
rect 46956 21586 47124 21588
rect 46956 21534 46958 21586
rect 47010 21534 47124 21586
rect 46956 21532 47124 21534
rect 47404 22540 47684 22596
rect 46956 21522 47012 21532
rect 47404 20804 47460 22540
rect 47180 20748 47460 20804
rect 47628 22370 47684 22382
rect 47628 22318 47630 22370
rect 47682 22318 47684 22370
rect 47628 21588 47684 22318
rect 47740 21924 47796 25004
rect 47852 24724 47908 25004
rect 47964 24948 48020 25452
rect 47964 24882 48020 24892
rect 48188 26516 48244 26526
rect 48636 26516 48692 29036
rect 48860 28868 48916 29372
rect 48748 28532 48804 28542
rect 48748 27076 48804 28476
rect 48860 28082 48916 28812
rect 48860 28030 48862 28082
rect 48914 28030 48916 28082
rect 48860 28018 48916 28030
rect 48972 29204 49028 29214
rect 48748 26962 48804 27020
rect 48748 26910 48750 26962
rect 48802 26910 48804 26962
rect 48748 26898 48804 26910
rect 48748 26516 48804 26526
rect 48636 26514 48804 26516
rect 48636 26462 48750 26514
rect 48802 26462 48804 26514
rect 48636 26460 48804 26462
rect 48076 24834 48132 24846
rect 48076 24782 48078 24834
rect 48130 24782 48132 24834
rect 47964 24724 48020 24734
rect 47852 24722 48020 24724
rect 47852 24670 47966 24722
rect 48018 24670 48020 24722
rect 47852 24668 48020 24670
rect 47964 24658 48020 24668
rect 47852 24050 47908 24062
rect 47852 23998 47854 24050
rect 47906 23998 47908 24050
rect 47852 23156 47908 23998
rect 47852 22596 47908 23100
rect 47852 22530 47908 22540
rect 47964 23940 48020 23950
rect 47964 22482 48020 23884
rect 47964 22430 47966 22482
rect 48018 22430 48020 22482
rect 47964 22418 48020 22430
rect 47852 22370 47908 22382
rect 47852 22318 47854 22370
rect 47906 22318 47908 22370
rect 47852 22260 47908 22318
rect 47852 22194 47908 22204
rect 48076 22148 48132 24782
rect 48188 23044 48244 26460
rect 48748 26450 48804 26460
rect 48972 26290 49028 29148
rect 48972 26238 48974 26290
rect 49026 26238 49028 26290
rect 48972 26226 49028 26238
rect 48748 26180 48804 26190
rect 48748 25618 48804 26124
rect 48748 25566 48750 25618
rect 48802 25566 48804 25618
rect 48748 25554 48804 25566
rect 48972 25508 49028 25518
rect 48636 25284 48692 25294
rect 48300 24722 48356 24734
rect 48300 24670 48302 24722
rect 48354 24670 48356 24722
rect 48300 23156 48356 24670
rect 48636 23938 48692 25228
rect 48636 23886 48638 23938
rect 48690 23886 48692 23938
rect 48636 23874 48692 23886
rect 48860 24612 48916 24622
rect 48860 23828 48916 24556
rect 48860 23762 48916 23772
rect 48972 23548 49028 25452
rect 48972 23492 49140 23548
rect 48748 23156 48804 23166
rect 48300 23154 48804 23156
rect 48300 23102 48750 23154
rect 48802 23102 48804 23154
rect 48300 23100 48804 23102
rect 48748 23090 48804 23100
rect 48188 22950 48244 22988
rect 48524 22260 48580 22270
rect 48076 22092 48468 22148
rect 47740 21858 47796 21868
rect 47964 21812 48020 21822
rect 47628 20802 47684 21532
rect 47628 20750 47630 20802
rect 47682 20750 47684 20802
rect 46396 19854 46398 19906
rect 46450 19854 46452 19906
rect 46396 19842 46452 19854
rect 46508 19964 46788 20020
rect 47068 20020 47124 20030
rect 46396 19348 46452 19358
rect 46396 19234 46452 19292
rect 46396 19182 46398 19234
rect 46450 19182 46452 19234
rect 46396 19170 46452 19182
rect 46284 18358 46340 18396
rect 46172 17054 46174 17106
rect 46226 17054 46228 17106
rect 46172 17042 46228 17054
rect 46396 18338 46452 18350
rect 46396 18286 46398 18338
rect 46450 18286 46452 18338
rect 45612 16046 45614 16098
rect 45666 16046 45668 16098
rect 45612 16034 45668 16046
rect 45500 15474 45556 15484
rect 45276 15092 45332 15102
rect 45388 15092 45668 15148
rect 45276 13636 45332 15036
rect 45276 13570 45332 13580
rect 45388 13522 45444 13534
rect 45388 13470 45390 13522
rect 45442 13470 45444 13522
rect 45388 13412 45444 13470
rect 45052 12350 45054 12402
rect 45106 12350 45108 12402
rect 45052 12338 45108 12350
rect 45276 13356 45444 13412
rect 45052 12178 45108 12190
rect 45052 12126 45054 12178
rect 45106 12126 45108 12178
rect 44940 11508 44996 11518
rect 44828 11506 44996 11508
rect 44828 11454 44942 11506
rect 44994 11454 44996 11506
rect 44828 11452 44996 11454
rect 44940 11442 44996 11452
rect 44716 11218 44772 11228
rect 44828 11284 44884 11294
rect 45052 11284 45108 12126
rect 45276 12180 45332 13356
rect 45388 13186 45444 13198
rect 45388 13134 45390 13186
rect 45442 13134 45444 13186
rect 45388 13074 45444 13134
rect 45388 13022 45390 13074
rect 45442 13022 45444 13074
rect 45388 13010 45444 13022
rect 45276 12114 45332 12124
rect 45612 12178 45668 15092
rect 45836 13186 45892 16940
rect 46060 15874 46116 15886
rect 46060 15822 46062 15874
rect 46114 15822 46116 15874
rect 46060 13748 46116 15822
rect 46172 14420 46228 14430
rect 46172 14326 46228 14364
rect 46060 13682 46116 13692
rect 45836 13134 45838 13186
rect 45890 13134 45892 13186
rect 45836 13122 45892 13134
rect 46060 13412 46116 13422
rect 46396 13412 46452 18286
rect 46508 18340 46564 19964
rect 46844 19908 46900 19918
rect 46508 18274 46564 18284
rect 46620 19906 46900 19908
rect 46620 19854 46846 19906
rect 46898 19854 46900 19906
rect 46620 19852 46900 19854
rect 46508 17892 46564 17902
rect 46620 17892 46676 19852
rect 46844 19842 46900 19852
rect 47068 19684 47124 19964
rect 46844 19628 47124 19684
rect 46844 19348 46900 19628
rect 47180 19572 47236 20748
rect 47628 20738 47684 20750
rect 47740 21698 47796 21710
rect 47740 21646 47742 21698
rect 47794 21646 47796 21698
rect 47516 20692 47572 20702
rect 46564 17836 46676 17892
rect 46732 19292 46844 19348
rect 46732 18564 46788 19292
rect 46844 19282 46900 19292
rect 46956 19516 47236 19572
rect 47292 20690 47572 20692
rect 47292 20638 47518 20690
rect 47570 20638 47572 20690
rect 47292 20636 47572 20638
rect 47292 20020 47348 20636
rect 47516 20626 47572 20636
rect 46844 19124 46900 19134
rect 46844 19030 46900 19068
rect 46956 18900 47012 19516
rect 47180 19346 47236 19358
rect 47180 19294 47182 19346
rect 47234 19294 47236 19346
rect 47068 19012 47124 19022
rect 47068 18918 47124 18956
rect 46956 18834 47012 18844
rect 46508 16994 46564 17836
rect 46508 16942 46510 16994
rect 46562 16942 46564 16994
rect 46508 16930 46564 16942
rect 46732 16770 46788 18508
rect 47180 17554 47236 19294
rect 47180 17502 47182 17554
rect 47234 17502 47236 17554
rect 47180 17490 47236 17502
rect 47068 17108 47124 17118
rect 47292 17108 47348 19964
rect 47628 20356 47684 20366
rect 47404 19796 47460 19806
rect 47404 19794 47572 19796
rect 47404 19742 47406 19794
rect 47458 19742 47572 19794
rect 47404 19740 47572 19742
rect 47404 19730 47460 19740
rect 47516 18452 47572 19740
rect 47628 19572 47684 20300
rect 47740 20132 47796 21646
rect 47740 20066 47796 20076
rect 47852 21476 47908 21486
rect 47852 20130 47908 21420
rect 47852 20078 47854 20130
rect 47906 20078 47908 20130
rect 47852 20066 47908 20078
rect 47964 20130 48020 21756
rect 48300 21700 48356 21710
rect 48300 21026 48356 21644
rect 48412 21364 48468 22092
rect 48524 21812 48580 22204
rect 48860 22258 48916 22270
rect 48860 22206 48862 22258
rect 48914 22206 48916 22258
rect 48860 21924 48916 22206
rect 49084 22260 49140 23492
rect 49084 22194 49140 22204
rect 48860 21868 49140 21924
rect 48524 21756 48804 21812
rect 48748 21698 48804 21756
rect 48748 21646 48750 21698
rect 48802 21646 48804 21698
rect 48748 21634 48804 21646
rect 48860 21700 48916 21868
rect 48860 21634 48916 21644
rect 48972 21698 49028 21710
rect 48972 21646 48974 21698
rect 49026 21646 49028 21698
rect 48972 21588 49028 21646
rect 49084 21698 49140 21868
rect 49084 21646 49086 21698
rect 49138 21646 49140 21698
rect 49084 21634 49140 21646
rect 48860 21476 48916 21486
rect 48972 21476 49028 21532
rect 49084 21476 49140 21486
rect 48972 21420 49084 21476
rect 48860 21382 48916 21420
rect 49084 21410 49140 21420
rect 48412 21298 48468 21308
rect 48300 20974 48302 21026
rect 48354 20974 48356 21026
rect 48300 20962 48356 20974
rect 48748 20692 48804 20702
rect 48748 20580 48804 20636
rect 47964 20078 47966 20130
rect 48018 20078 48020 20130
rect 47964 20066 48020 20078
rect 48636 20578 48804 20580
rect 48636 20526 48750 20578
rect 48802 20526 48804 20578
rect 48636 20524 48804 20526
rect 47852 19796 47908 19806
rect 47852 19794 48580 19796
rect 47852 19742 47854 19794
rect 47906 19742 48580 19794
rect 47852 19740 48580 19742
rect 47852 19730 47908 19740
rect 47628 19516 48020 19572
rect 47740 19236 47796 19246
rect 47628 18452 47684 18462
rect 47516 18450 47684 18452
rect 47516 18398 47630 18450
rect 47682 18398 47684 18450
rect 47516 18396 47684 18398
rect 47628 18386 47684 18396
rect 47068 17106 47348 17108
rect 47068 17054 47070 17106
rect 47122 17054 47348 17106
rect 47068 17052 47348 17054
rect 47068 17042 47124 17052
rect 46732 16718 46734 16770
rect 46786 16718 46788 16770
rect 46732 16706 46788 16718
rect 47404 16994 47460 17006
rect 47404 16942 47406 16994
rect 47458 16942 47460 16994
rect 47292 16658 47348 16670
rect 47292 16606 47294 16658
rect 47346 16606 47348 16658
rect 46508 16212 46564 16222
rect 46508 15428 46564 16156
rect 46620 16100 46676 16110
rect 47068 16100 47124 16110
rect 46620 16098 47124 16100
rect 46620 16046 46622 16098
rect 46674 16046 47070 16098
rect 47122 16046 47124 16098
rect 46620 16044 47124 16046
rect 46620 16034 46676 16044
rect 46620 15428 46676 15438
rect 46508 15426 46676 15428
rect 46508 15374 46622 15426
rect 46674 15374 46676 15426
rect 46508 15372 46676 15374
rect 46508 14420 46564 15372
rect 46620 15362 46676 15372
rect 47068 15428 47124 16044
rect 47068 15362 47124 15372
rect 47180 14980 47236 14990
rect 47180 14754 47236 14924
rect 47180 14702 47182 14754
rect 47234 14702 47236 14754
rect 47180 14690 47236 14702
rect 47068 14420 47124 14430
rect 46564 14364 46788 14420
rect 46508 14354 46564 14364
rect 46732 13970 46788 14364
rect 47068 14326 47124 14364
rect 46732 13918 46734 13970
rect 46786 13918 46788 13970
rect 46732 13906 46788 13918
rect 46844 14308 46900 14318
rect 46732 13748 46788 13758
rect 46396 13356 46564 13412
rect 46060 12850 46116 13356
rect 46060 12798 46062 12850
rect 46114 12798 46116 12850
rect 46060 12786 46116 12798
rect 45612 12126 45614 12178
rect 45666 12126 45668 12178
rect 45612 12114 45668 12126
rect 46172 12178 46228 12190
rect 46172 12126 46174 12178
rect 46226 12126 46228 12178
rect 46172 11508 46228 12126
rect 45388 11506 46228 11508
rect 45388 11454 46174 11506
rect 46226 11454 46228 11506
rect 45388 11452 46228 11454
rect 45388 11394 45444 11452
rect 46172 11442 46228 11452
rect 45388 11342 45390 11394
rect 45442 11342 45444 11394
rect 45388 11330 45444 11342
rect 46396 11394 46452 11406
rect 46396 11342 46398 11394
rect 46450 11342 46452 11394
rect 44828 11282 45108 11284
rect 44828 11230 44830 11282
rect 44882 11230 45108 11282
rect 44828 11228 45108 11230
rect 45164 11284 45220 11294
rect 44044 11170 44100 11182
rect 44044 11118 44046 11170
rect 44098 11118 44100 11170
rect 44044 8820 44100 11118
rect 44604 10164 44660 10174
rect 44268 9828 44324 9838
rect 44268 9734 44324 9772
rect 44156 9602 44212 9614
rect 44156 9550 44158 9602
rect 44210 9550 44212 9602
rect 44156 9044 44212 9550
rect 44604 9268 44660 10108
rect 44828 9828 44884 11228
rect 45164 11172 45220 11228
rect 45724 11282 45780 11294
rect 45724 11230 45726 11282
rect 45778 11230 45780 11282
rect 45724 11172 45780 11230
rect 45164 11116 45780 11172
rect 45948 11282 46004 11294
rect 45948 11230 45950 11282
rect 46002 11230 46004 11282
rect 45164 10834 45220 11116
rect 45948 10948 46004 11230
rect 45948 10882 46004 10892
rect 45164 10782 45166 10834
rect 45218 10782 45220 10834
rect 45164 10770 45220 10782
rect 46396 10836 46452 11342
rect 46396 10770 46452 10780
rect 46508 10834 46564 13356
rect 46732 12962 46788 13692
rect 46844 13074 46900 14252
rect 46844 13022 46846 13074
rect 46898 13022 46900 13074
rect 46844 13010 46900 13022
rect 47068 13076 47124 13086
rect 46732 12910 46734 12962
rect 46786 12910 46788 12962
rect 46732 12898 46788 12910
rect 46956 12178 47012 12190
rect 46956 12126 46958 12178
rect 47010 12126 47012 12178
rect 46844 11508 46900 11518
rect 46844 11414 46900 11452
rect 46956 10836 47012 12126
rect 47068 12066 47124 13020
rect 47292 12962 47348 16606
rect 47404 16210 47460 16942
rect 47628 16884 47684 16894
rect 47404 16158 47406 16210
rect 47458 16158 47460 16210
rect 47404 16100 47460 16158
rect 47404 16034 47460 16044
rect 47516 16882 47684 16884
rect 47516 16830 47630 16882
rect 47682 16830 47684 16882
rect 47516 16828 47684 16830
rect 47516 15148 47572 16828
rect 47628 16818 47684 16828
rect 47740 16772 47796 19180
rect 47852 17668 47908 17678
rect 47964 17668 48020 19516
rect 48412 19122 48468 19134
rect 48412 19070 48414 19122
rect 48466 19070 48468 19122
rect 48300 17780 48356 17790
rect 48412 17780 48468 19070
rect 48300 17778 48468 17780
rect 48300 17726 48302 17778
rect 48354 17726 48468 17778
rect 48300 17724 48468 17726
rect 48300 17714 48356 17724
rect 48188 17668 48244 17678
rect 47964 17666 48244 17668
rect 47964 17614 48190 17666
rect 48242 17614 48244 17666
rect 47964 17612 48244 17614
rect 47852 17574 47908 17612
rect 48188 17602 48244 17612
rect 48412 17556 48468 17566
rect 48524 17556 48580 19740
rect 48636 17892 48692 20524
rect 48748 20514 48804 20524
rect 49084 20580 49140 20590
rect 48860 20132 48916 20142
rect 48860 20038 48916 20076
rect 48748 20018 48804 20030
rect 48748 19966 48750 20018
rect 48802 19966 48804 20018
rect 48748 19908 48804 19966
rect 48748 19842 48804 19852
rect 48972 20018 49028 20030
rect 48972 19966 48974 20018
rect 49026 19966 49028 20018
rect 48748 18564 48804 18574
rect 48748 18450 48804 18508
rect 48748 18398 48750 18450
rect 48802 18398 48804 18450
rect 48748 18386 48804 18398
rect 48860 18452 48916 18462
rect 48972 18452 49028 19966
rect 49084 19236 49140 20524
rect 49196 19460 49252 30828
rect 49420 30212 49476 30222
rect 49308 30210 49476 30212
rect 49308 30158 49422 30210
rect 49474 30158 49476 30210
rect 49308 30156 49476 30158
rect 49308 29650 49364 30156
rect 49420 30146 49476 30156
rect 49308 29598 49310 29650
rect 49362 29598 49364 29650
rect 49308 29586 49364 29598
rect 49644 26908 49700 38612
rect 49756 30098 49812 40348
rect 49980 39618 50036 39630
rect 49980 39566 49982 39618
rect 50034 39566 50036 39618
rect 49980 39508 50036 39566
rect 49980 39442 50036 39452
rect 50092 39284 50148 40460
rect 49980 39228 50148 39284
rect 49868 38836 49924 38846
rect 49868 38742 49924 38780
rect 49980 38668 50036 39228
rect 50204 38668 50260 40908
rect 50316 40290 50372 42028
rect 50428 40404 50484 44044
rect 50652 44034 50708 44044
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50764 43540 50820 43550
rect 50764 42980 50820 43484
rect 50876 43540 50932 43550
rect 50988 43540 51044 44270
rect 50876 43538 51044 43540
rect 50876 43486 50878 43538
rect 50930 43486 51044 43538
rect 50876 43484 51044 43486
rect 50876 43474 50932 43484
rect 51324 43428 51380 45838
rect 51436 44994 51492 46060
rect 51548 46004 51604 46014
rect 51548 45910 51604 45948
rect 51660 45668 51716 46284
rect 51436 44942 51438 44994
rect 51490 44942 51492 44994
rect 51436 44930 51492 44942
rect 51548 45612 51716 45668
rect 51772 46284 51884 46340
rect 51548 45444 51604 45612
rect 51324 43362 51380 43372
rect 50876 42980 50932 42990
rect 50764 42978 50932 42980
rect 50764 42926 50878 42978
rect 50930 42926 50932 42978
rect 50764 42924 50932 42926
rect 50876 42914 50932 42924
rect 51212 42980 51268 42990
rect 51212 42886 51268 42924
rect 51548 42756 51604 45388
rect 51772 44772 51828 46284
rect 51884 46274 51940 46284
rect 51996 45780 52052 45790
rect 51884 45668 51940 45678
rect 51884 45574 51940 45612
rect 51548 42690 51604 42700
rect 51660 44716 51828 44772
rect 51884 45444 51940 45454
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 51548 42196 51604 42206
rect 50540 41860 50596 41870
rect 50540 41766 50596 41804
rect 51100 41858 51156 41870
rect 51100 41806 51102 41858
rect 51154 41806 51156 41858
rect 50764 40964 50820 41002
rect 50764 40898 50820 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50428 40338 50484 40348
rect 50316 40238 50318 40290
rect 50370 40238 50372 40290
rect 50316 39732 50372 40238
rect 50316 39666 50372 39676
rect 50428 39620 50484 39630
rect 49868 38612 50036 38668
rect 50092 38612 50260 38668
rect 50316 39508 50372 39518
rect 50316 38948 50372 39452
rect 50428 39060 50484 39564
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50428 38994 50484 39004
rect 50316 38724 50372 38892
rect 50764 38724 50820 38734
rect 50316 38722 50484 38724
rect 50316 38670 50318 38722
rect 50370 38670 50484 38722
rect 50316 38668 50484 38670
rect 50316 38658 50372 38668
rect 49868 37940 49924 38612
rect 49868 37874 49924 37884
rect 49868 37716 49924 37726
rect 49868 35812 49924 37660
rect 50092 36148 50148 38612
rect 50316 37938 50372 37950
rect 50316 37886 50318 37938
rect 50370 37886 50372 37938
rect 50316 37380 50372 37886
rect 50428 37380 50484 38668
rect 50764 38052 50820 38668
rect 50764 37958 50820 37996
rect 50876 38722 50932 38734
rect 50876 38670 50878 38722
rect 50930 38670 50932 38722
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50428 37324 50596 37380
rect 50316 37286 50372 37324
rect 50204 37266 50260 37278
rect 50204 37214 50206 37266
rect 50258 37214 50260 37266
rect 50204 37044 50260 37214
rect 50204 36978 50260 36988
rect 50204 36820 50260 36830
rect 50204 36482 50260 36764
rect 50540 36708 50596 37324
rect 50540 36642 50596 36652
rect 50204 36430 50206 36482
rect 50258 36430 50260 36482
rect 50204 36418 50260 36430
rect 50428 36482 50484 36494
rect 50428 36430 50430 36482
rect 50482 36430 50484 36482
rect 50092 36092 50372 36148
rect 49868 35756 50148 35812
rect 50092 35700 50148 35756
rect 50092 35698 50260 35700
rect 50092 35646 50094 35698
rect 50146 35646 50260 35698
rect 50092 35644 50260 35646
rect 50092 35634 50148 35644
rect 49868 35364 49924 35374
rect 49924 35308 50148 35364
rect 49868 34130 49924 35308
rect 50092 35138 50148 35308
rect 50092 35086 50094 35138
rect 50146 35086 50148 35138
rect 50092 35074 50148 35086
rect 49868 34078 49870 34130
rect 49922 34078 49924 34130
rect 49868 34066 49924 34078
rect 49980 34916 50036 34926
rect 49980 34130 50036 34860
rect 50204 34356 50260 35644
rect 49980 34078 49982 34130
rect 50034 34078 50036 34130
rect 49980 34066 50036 34078
rect 50092 34300 50260 34356
rect 50092 33460 50148 34300
rect 50092 33394 50148 33404
rect 50204 34132 50260 34142
rect 50204 32900 50260 34076
rect 50316 33572 50372 36092
rect 50428 35252 50484 36430
rect 50876 36372 50932 38670
rect 51100 37828 51156 41806
rect 51324 41188 51380 41198
rect 51324 41186 51492 41188
rect 51324 41134 51326 41186
rect 51378 41134 51492 41186
rect 51324 41132 51492 41134
rect 51324 41122 51380 41132
rect 51436 39620 51492 41132
rect 51436 39554 51492 39564
rect 51548 38836 51604 42140
rect 51660 41860 51716 44716
rect 51772 44546 51828 44558
rect 51772 44494 51774 44546
rect 51826 44494 51828 44546
rect 51772 43540 51828 44494
rect 51884 44212 51940 45388
rect 51996 44436 52052 45724
rect 51996 44380 52164 44436
rect 51996 44212 52052 44222
rect 51884 44210 52052 44212
rect 51884 44158 51998 44210
rect 52050 44158 52052 44210
rect 51884 44156 52052 44158
rect 51996 44146 52052 44156
rect 51996 43764 52052 43774
rect 51772 43474 51828 43484
rect 51884 43708 51996 43764
rect 51772 42868 51828 42878
rect 51772 42754 51828 42812
rect 51772 42702 51774 42754
rect 51826 42702 51828 42754
rect 51772 42690 51828 42702
rect 51660 41794 51716 41804
rect 51884 41412 51940 43708
rect 51996 43698 52052 43708
rect 52108 43540 52164 44380
rect 51996 43484 52164 43540
rect 51996 42642 52052 43484
rect 51996 42590 51998 42642
rect 52050 42590 52052 42642
rect 51996 42578 52052 42590
rect 52108 42756 52164 42766
rect 51996 42084 52052 42094
rect 51996 41990 52052 42028
rect 51772 41356 51940 41412
rect 51996 41860 52052 41870
rect 51772 40740 51828 41356
rect 51996 41298 52052 41804
rect 51996 41246 51998 41298
rect 52050 41246 52052 41298
rect 51996 41234 52052 41246
rect 52108 41076 52164 42700
rect 52444 42532 52500 47180
rect 52668 46340 52724 47182
rect 52892 46900 52948 48974
rect 53116 48020 53172 49644
rect 53116 47964 53396 48020
rect 53228 47796 53284 47806
rect 53116 47572 53172 47582
rect 52892 46834 52948 46844
rect 53004 47570 53172 47572
rect 53004 47518 53118 47570
rect 53170 47518 53172 47570
rect 53004 47516 53172 47518
rect 52668 46274 52724 46284
rect 53004 46004 53060 47516
rect 53116 47506 53172 47516
rect 52668 45948 53060 46004
rect 52668 44996 52724 45948
rect 53116 45892 53172 45902
rect 52892 45890 53172 45892
rect 52892 45838 53118 45890
rect 53170 45838 53172 45890
rect 52892 45836 53172 45838
rect 53228 45892 53284 47740
rect 53340 46898 53396 47964
rect 53340 46846 53342 46898
rect 53394 46846 53396 46898
rect 53340 46834 53396 46846
rect 53340 45892 53396 45902
rect 53228 45836 53340 45892
rect 52668 44322 52724 44940
rect 52668 44270 52670 44322
rect 52722 44270 52724 44322
rect 52668 43538 52724 44270
rect 52780 45666 52836 45678
rect 52780 45614 52782 45666
rect 52834 45614 52836 45666
rect 52780 43764 52836 45614
rect 52892 43988 52948 45836
rect 53116 45826 53172 45836
rect 53340 45778 53396 45836
rect 53340 45726 53342 45778
rect 53394 45726 53396 45778
rect 53340 45714 53396 45726
rect 53340 45556 53396 45566
rect 53228 45108 53284 45118
rect 53228 44994 53284 45052
rect 53340 45106 53396 45500
rect 53340 45054 53342 45106
rect 53394 45054 53396 45106
rect 53340 45042 53396 45054
rect 53228 44942 53230 44994
rect 53282 44942 53284 44994
rect 53228 44930 53284 44942
rect 53340 44660 53396 44670
rect 52892 43922 52948 43932
rect 53116 44548 53172 44558
rect 53116 44210 53172 44492
rect 53228 44436 53284 44446
rect 53340 44436 53396 44604
rect 53228 44434 53396 44436
rect 53228 44382 53230 44434
rect 53282 44382 53396 44434
rect 53228 44380 53396 44382
rect 53228 44370 53284 44380
rect 53452 44324 53508 50372
rect 53564 47682 53620 50540
rect 53676 50148 53732 50158
rect 53676 49588 53732 50092
rect 53788 49812 53844 52556
rect 53788 49746 53844 49756
rect 53900 52388 53956 52398
rect 53900 52162 53956 52332
rect 54124 52276 54180 55134
rect 54236 54068 54292 55916
rect 54460 54514 54516 57374
rect 54796 57426 54852 57438
rect 54796 57374 54798 57426
rect 54850 57374 54852 57426
rect 54796 56868 54852 57374
rect 55020 57092 55076 57102
rect 55020 56998 55076 57036
rect 54796 56308 54852 56812
rect 54796 56242 54852 56252
rect 54908 56644 54964 56654
rect 54908 56082 54964 56588
rect 55356 56306 55412 57820
rect 56700 57876 56756 57886
rect 56756 57820 56868 57876
rect 56700 57810 56756 57820
rect 55916 57764 55972 57774
rect 55804 57650 55860 57662
rect 55804 57598 55806 57650
rect 55858 57598 55860 57650
rect 55468 57540 55524 57550
rect 55524 57484 55636 57540
rect 55468 57446 55524 57484
rect 55468 56754 55524 56766
rect 55468 56702 55470 56754
rect 55522 56702 55524 56754
rect 55468 56644 55524 56702
rect 55580 56644 55636 57484
rect 55804 57092 55860 57598
rect 55804 57026 55860 57036
rect 55692 56868 55748 56878
rect 55692 56774 55748 56812
rect 55580 56588 55748 56644
rect 55468 56578 55524 56588
rect 55356 56254 55358 56306
rect 55410 56254 55412 56306
rect 55356 56242 55412 56254
rect 55580 56196 55636 56206
rect 55580 56102 55636 56140
rect 54908 56030 54910 56082
rect 54962 56030 54964 56082
rect 54908 56018 54964 56030
rect 55132 56082 55188 56094
rect 55132 56030 55134 56082
rect 55186 56030 55188 56082
rect 55132 55524 55188 56030
rect 55356 55970 55412 55982
rect 55356 55918 55358 55970
rect 55410 55918 55412 55970
rect 55356 55636 55412 55918
rect 55356 55580 55524 55636
rect 55188 55468 55412 55524
rect 55132 55458 55188 55468
rect 55356 55188 55412 55468
rect 55468 55412 55524 55580
rect 55468 55346 55524 55356
rect 55580 55300 55636 55310
rect 55692 55300 55748 56588
rect 55804 55524 55860 55534
rect 55916 55524 55972 57708
rect 56812 57762 56868 57820
rect 56812 57710 56814 57762
rect 56866 57710 56868 57762
rect 56364 57092 56420 57102
rect 56364 56978 56420 57036
rect 56364 56926 56366 56978
rect 56418 56926 56420 56978
rect 56364 56914 56420 56926
rect 55804 55522 55972 55524
rect 55804 55470 55806 55522
rect 55858 55470 55972 55522
rect 55804 55468 55972 55470
rect 55804 55458 55860 55468
rect 55580 55298 55748 55300
rect 55580 55246 55582 55298
rect 55634 55246 55748 55298
rect 55580 55244 55748 55246
rect 55468 55188 55524 55198
rect 55356 55186 55524 55188
rect 55356 55134 55470 55186
rect 55522 55134 55524 55186
rect 55356 55132 55524 55134
rect 55468 55122 55524 55132
rect 55580 54964 55636 55244
rect 55916 55188 55972 55468
rect 55916 55122 55972 55132
rect 56028 56642 56084 56654
rect 56028 56590 56030 56642
rect 56082 56590 56084 56642
rect 55468 54908 55636 54964
rect 54460 54462 54462 54514
rect 54514 54462 54516 54514
rect 54460 54450 54516 54462
rect 54684 54516 54740 54526
rect 54348 54292 54404 54302
rect 54348 54198 54404 54236
rect 54236 54012 54516 54068
rect 54236 52946 54292 52958
rect 54236 52894 54238 52946
rect 54290 52894 54292 52946
rect 54236 52612 54292 52894
rect 54348 52836 54404 52846
rect 54348 52742 54404 52780
rect 54348 52612 54404 52622
rect 54236 52556 54348 52612
rect 54348 52546 54404 52556
rect 54460 52500 54516 54012
rect 54460 52434 54516 52444
rect 54124 52220 54628 52276
rect 53900 52110 53902 52162
rect 53954 52110 53956 52162
rect 53788 49588 53844 49598
rect 53676 49532 53788 49588
rect 53788 49028 53844 49532
rect 53564 47630 53566 47682
rect 53618 47630 53620 47682
rect 53564 47618 53620 47630
rect 53676 49026 53844 49028
rect 53676 48974 53790 49026
rect 53842 48974 53844 49026
rect 53676 48972 53844 48974
rect 53676 47570 53732 48972
rect 53788 48962 53844 48972
rect 53900 48468 53956 52110
rect 54124 52050 54180 52062
rect 54124 51998 54126 52050
rect 54178 51998 54180 52050
rect 54124 51044 54180 51998
rect 54124 50978 54180 50988
rect 54236 52052 54292 52062
rect 54236 51380 54292 51996
rect 54572 51940 54628 52220
rect 54684 52164 54740 54460
rect 55132 53732 55188 53742
rect 55132 53638 55188 53676
rect 55132 53172 55188 53182
rect 55020 53060 55076 53070
rect 55020 52966 55076 53004
rect 54796 52946 54852 52958
rect 54796 52894 54798 52946
rect 54850 52894 54852 52946
rect 54796 52500 54852 52894
rect 54796 52434 54852 52444
rect 54796 52164 54852 52174
rect 54684 52162 54852 52164
rect 54684 52110 54798 52162
rect 54850 52110 54852 52162
rect 54684 52108 54852 52110
rect 54796 52098 54852 52108
rect 54572 51884 54964 51940
rect 54348 51380 54404 51390
rect 54236 51378 54404 51380
rect 54236 51326 54350 51378
rect 54402 51326 54404 51378
rect 54236 51324 54404 51326
rect 54236 50594 54292 51324
rect 54348 51314 54404 51324
rect 54572 51380 54628 51390
rect 54572 51286 54628 51324
rect 54236 50542 54238 50594
rect 54290 50542 54292 50594
rect 54236 50428 54292 50542
rect 54236 50372 54852 50428
rect 54796 50034 54852 50372
rect 54796 49982 54798 50034
rect 54850 49982 54852 50034
rect 54796 49970 54852 49982
rect 54908 50036 54964 51884
rect 55020 51156 55076 51166
rect 55132 51156 55188 53116
rect 55020 51154 55188 51156
rect 55020 51102 55022 51154
rect 55074 51102 55188 51154
rect 55020 51100 55188 51102
rect 55356 53060 55412 53070
rect 55020 51090 55076 51100
rect 54908 49970 54964 49980
rect 55244 50594 55300 50606
rect 55244 50542 55246 50594
rect 55298 50542 55300 50594
rect 55244 50036 55300 50542
rect 55356 50428 55412 53004
rect 55468 52612 55524 54908
rect 56028 54852 56084 56590
rect 56476 56644 56532 56654
rect 56140 55972 56196 55982
rect 56140 55970 56308 55972
rect 56140 55918 56142 55970
rect 56194 55918 56308 55970
rect 56140 55916 56308 55918
rect 56140 55906 56196 55916
rect 56028 54786 56084 54796
rect 56140 55524 56196 55534
rect 55692 54740 55748 54750
rect 55692 54402 55748 54684
rect 55692 54350 55694 54402
rect 55746 54350 55748 54402
rect 55580 53730 55636 53742
rect 55580 53678 55582 53730
rect 55634 53678 55636 53730
rect 55580 53172 55636 53678
rect 55580 53106 55636 53116
rect 55580 52724 55636 52734
rect 55580 52630 55636 52668
rect 55468 52162 55524 52556
rect 55692 52274 55748 54350
rect 55916 54628 55972 54638
rect 56140 54628 56196 55468
rect 55916 54626 56196 54628
rect 55916 54574 55918 54626
rect 55970 54574 56196 54626
rect 55916 54572 56196 54574
rect 55916 53730 55972 54572
rect 55916 53678 55918 53730
rect 55970 53678 55972 53730
rect 55916 53666 55972 53678
rect 56252 53172 56308 55916
rect 56476 55524 56532 56588
rect 56812 56308 56868 57710
rect 56700 55860 56756 55870
rect 56476 55458 56532 55468
rect 56588 55858 56756 55860
rect 56588 55806 56702 55858
rect 56754 55806 56756 55858
rect 56588 55804 56756 55806
rect 56588 54740 56644 55804
rect 56700 55794 56756 55804
rect 56812 55636 56868 56252
rect 56924 56980 56980 56990
rect 56924 56084 56980 56924
rect 57820 56980 57876 56990
rect 57820 56886 57876 56924
rect 57036 56868 57092 56878
rect 57036 56754 57092 56812
rect 57036 56702 57038 56754
rect 57090 56702 57092 56754
rect 57036 56690 57092 56702
rect 57260 56866 57316 56878
rect 57260 56814 57262 56866
rect 57314 56814 57316 56866
rect 57260 56756 57316 56814
rect 57260 56690 57316 56700
rect 58268 56756 58324 56766
rect 58268 56662 58324 56700
rect 59052 56756 59108 56766
rect 59108 56700 59220 56756
rect 59052 56690 59108 56700
rect 57708 56364 58324 56420
rect 57036 56084 57092 56094
rect 56924 56082 57092 56084
rect 56924 56030 57038 56082
rect 57090 56030 57092 56082
rect 56924 56028 57092 56030
rect 57036 56018 57092 56028
rect 57708 56082 57764 56364
rect 57820 56196 57876 56206
rect 57876 56140 58212 56196
rect 57820 56102 57876 56140
rect 57708 56030 57710 56082
rect 57762 56030 57764 56082
rect 57708 56018 57764 56030
rect 56700 55580 56868 55636
rect 57260 55636 57316 55646
rect 56700 55298 56756 55580
rect 56700 55246 56702 55298
rect 56754 55246 56756 55298
rect 56700 55234 56756 55246
rect 56812 55412 56868 55422
rect 56588 54674 56644 54684
rect 56588 54514 56644 54526
rect 56588 54462 56590 54514
rect 56642 54462 56644 54514
rect 56588 54404 56644 54462
rect 56588 54338 56644 54348
rect 56700 54290 56756 54302
rect 56700 54238 56702 54290
rect 56754 54238 56756 54290
rect 56700 53732 56756 54238
rect 56700 53666 56756 53676
rect 55692 52222 55694 52274
rect 55746 52222 55748 52274
rect 55692 52210 55748 52222
rect 55916 52722 55972 52734
rect 55916 52670 55918 52722
rect 55970 52670 55972 52722
rect 55468 52110 55470 52162
rect 55522 52110 55524 52162
rect 55468 52098 55524 52110
rect 55916 51604 55972 52670
rect 55916 51538 55972 51548
rect 55692 50596 55748 50634
rect 55748 50540 55860 50596
rect 55692 50530 55748 50540
rect 55356 50372 55748 50428
rect 55244 49970 55300 49980
rect 55692 49922 55748 50372
rect 55692 49870 55694 49922
rect 55746 49870 55748 49922
rect 54236 49812 54292 49822
rect 54236 49718 54292 49756
rect 55356 49700 55412 49710
rect 55244 49644 55356 49700
rect 55132 49588 55188 49598
rect 54348 49586 55188 49588
rect 54348 49534 55134 49586
rect 55186 49534 55188 49586
rect 54348 49532 55188 49534
rect 54348 49140 54404 49532
rect 55132 49522 55188 49532
rect 54572 49252 54628 49262
rect 54572 49158 54628 49196
rect 54012 49084 54404 49140
rect 54012 48914 54068 49084
rect 54012 48862 54014 48914
rect 54066 48862 54068 48914
rect 54012 48850 54068 48862
rect 53900 48412 54292 48468
rect 53676 47518 53678 47570
rect 53730 47518 53732 47570
rect 53676 47506 53732 47518
rect 53900 47236 53956 47246
rect 53676 46900 53732 46910
rect 53676 46806 53732 46844
rect 53900 46786 53956 47180
rect 53900 46734 53902 46786
rect 53954 46734 53956 46786
rect 53900 46722 53956 46734
rect 54236 46788 54292 48412
rect 54348 48466 54404 49084
rect 54348 48414 54350 48466
rect 54402 48414 54404 48466
rect 54348 48402 54404 48414
rect 54908 48802 54964 48814
rect 54908 48750 54910 48802
rect 54962 48750 54964 48802
rect 54572 48242 54628 48254
rect 54572 48190 54574 48242
rect 54626 48190 54628 48242
rect 54460 46788 54516 46798
rect 54236 46786 54516 46788
rect 54236 46734 54462 46786
rect 54514 46734 54516 46786
rect 54236 46732 54516 46734
rect 54460 46722 54516 46732
rect 53788 46564 53844 46574
rect 53564 46450 53620 46462
rect 53564 46398 53566 46450
rect 53618 46398 53620 46450
rect 53564 45556 53620 46398
rect 53564 45490 53620 45500
rect 53788 45330 53844 46508
rect 54348 46562 54404 46574
rect 54348 46510 54350 46562
rect 54402 46510 54404 46562
rect 54348 46452 54404 46510
rect 53788 45278 53790 45330
rect 53842 45278 53844 45330
rect 53676 45218 53732 45230
rect 53676 45166 53678 45218
rect 53730 45166 53732 45218
rect 53676 45108 53732 45166
rect 53676 45042 53732 45052
rect 53452 44268 53732 44324
rect 53116 44158 53118 44210
rect 53170 44158 53172 44210
rect 52780 43698 52836 43708
rect 52668 43486 52670 43538
rect 52722 43486 52724 43538
rect 52668 43474 52724 43486
rect 52892 43540 52948 43550
rect 52892 43446 52948 43484
rect 52780 43092 52836 43102
rect 52780 42978 52836 43036
rect 52780 42926 52782 42978
rect 52834 42926 52836 42978
rect 52780 42914 52836 42926
rect 52892 42756 52948 42766
rect 52892 42662 52948 42700
rect 53116 42644 53172 44158
rect 53228 44098 53284 44110
rect 53228 44046 53230 44098
rect 53282 44046 53284 44098
rect 53228 43876 53284 44046
rect 53228 43810 53284 43820
rect 53452 44098 53508 44110
rect 53452 44046 53454 44098
rect 53506 44046 53508 44098
rect 53452 42980 53508 44046
rect 53564 43988 53620 43998
rect 53564 43316 53620 43932
rect 53564 43250 53620 43260
rect 53452 42756 53508 42924
rect 53452 42690 53508 42700
rect 53228 42644 53284 42654
rect 53116 42642 53284 42644
rect 53116 42590 53230 42642
rect 53282 42590 53284 42642
rect 53116 42588 53284 42590
rect 53228 42578 53284 42588
rect 52444 42476 53060 42532
rect 52332 42084 52388 42094
rect 51884 41020 52164 41076
rect 52220 42028 52332 42084
rect 51884 40962 51940 41020
rect 51884 40910 51886 40962
rect 51938 40910 51940 40962
rect 51884 40898 51940 40910
rect 51772 40684 52052 40740
rect 51996 39618 52052 40684
rect 52108 39844 52164 39854
rect 52220 39844 52276 42028
rect 52332 42018 52388 42028
rect 52668 41972 52724 41982
rect 52108 39842 52276 39844
rect 52108 39790 52110 39842
rect 52162 39790 52276 39842
rect 52108 39788 52276 39790
rect 52332 41188 52388 41198
rect 52108 39778 52164 39788
rect 51996 39566 51998 39618
rect 52050 39566 52052 39618
rect 51996 39554 52052 39566
rect 51772 39396 51828 39406
rect 51772 38946 51828 39340
rect 51772 38894 51774 38946
rect 51826 38894 51828 38946
rect 51772 38882 51828 38894
rect 52108 39284 52164 39294
rect 51548 38770 51604 38780
rect 51996 38834 52052 38846
rect 51996 38782 51998 38834
rect 52050 38782 52052 38834
rect 51212 38612 51268 38622
rect 51212 38518 51268 38556
rect 51548 38612 51604 38622
rect 51604 38556 51716 38612
rect 51548 38546 51604 38556
rect 51100 37762 51156 37772
rect 51212 37492 51268 37502
rect 51212 37490 51492 37492
rect 51212 37438 51214 37490
rect 51266 37438 51492 37490
rect 51212 37436 51492 37438
rect 51212 37426 51268 37436
rect 51100 37268 51156 37278
rect 50876 36306 50932 36316
rect 50988 36820 51044 36830
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50988 35924 51044 36764
rect 50428 35186 50484 35196
rect 50652 35868 51044 35924
rect 50428 34916 50484 34926
rect 50652 34916 50708 35868
rect 50428 34914 50708 34916
rect 50428 34862 50430 34914
rect 50482 34862 50708 34914
rect 50428 34860 50708 34862
rect 50988 35588 51044 35598
rect 50428 34356 50484 34860
rect 50988 34802 51044 35532
rect 50988 34750 50990 34802
rect 51042 34750 51044 34802
rect 50988 34738 51044 34750
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50428 34290 50484 34300
rect 51100 34244 51156 37212
rect 50876 34188 51156 34244
rect 51212 35252 51268 35262
rect 51212 34914 51268 35196
rect 51212 34862 51214 34914
rect 51266 34862 51268 34914
rect 50764 33572 50820 33582
rect 50876 33572 50932 34188
rect 50316 33516 50484 33572
rect 49980 32844 50260 32900
rect 49980 32338 50036 32844
rect 50428 32788 50484 33516
rect 50764 33570 50932 33572
rect 50764 33518 50766 33570
rect 50818 33518 50932 33570
rect 50764 33516 50932 33518
rect 50988 34020 51044 34030
rect 51212 34020 51268 34862
rect 51212 33964 51380 34020
rect 50764 33506 50820 33516
rect 50988 33124 51044 33964
rect 51324 33570 51380 33964
rect 51324 33518 51326 33570
rect 51378 33518 51380 33570
rect 51324 33506 51380 33518
rect 50876 33068 50988 33124
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50428 32732 50596 32788
rect 50540 32562 50596 32732
rect 50540 32510 50542 32562
rect 50594 32510 50596 32562
rect 50428 32450 50484 32462
rect 50428 32398 50430 32450
rect 50482 32398 50484 32450
rect 49980 32286 49982 32338
rect 50034 32286 50036 32338
rect 49980 32116 50036 32286
rect 49980 32050 50036 32060
rect 50204 32338 50260 32350
rect 50204 32286 50206 32338
rect 50258 32286 50260 32338
rect 50204 30324 50260 32286
rect 49756 30046 49758 30098
rect 49810 30046 49812 30098
rect 49756 30034 49812 30046
rect 49980 30268 50260 30324
rect 49756 29540 49812 29550
rect 49812 29484 49924 29540
rect 49756 29474 49812 29484
rect 49756 28980 49812 28990
rect 49756 28420 49812 28924
rect 49868 28866 49924 29484
rect 49868 28814 49870 28866
rect 49922 28814 49924 28866
rect 49868 28644 49924 28814
rect 49868 28578 49924 28588
rect 49756 28364 49924 28420
rect 49756 27300 49812 27310
rect 49756 27206 49812 27244
rect 49532 26852 49700 26908
rect 49756 26964 49812 26974
rect 49420 25508 49476 25518
rect 49420 25414 49476 25452
rect 49308 25396 49364 25406
rect 49308 24946 49364 25340
rect 49532 24948 49588 26852
rect 49756 26514 49812 26908
rect 49868 26962 49924 28364
rect 49980 27748 50036 30268
rect 50204 30100 50260 30110
rect 50092 30044 50204 30100
rect 50092 28532 50148 30044
rect 50204 30034 50260 30044
rect 50204 29540 50260 29550
rect 50204 29538 50372 29540
rect 50204 29486 50206 29538
rect 50258 29486 50372 29538
rect 50204 29484 50372 29486
rect 50204 29474 50260 29484
rect 50204 28532 50260 28542
rect 50092 28530 50260 28532
rect 50092 28478 50206 28530
rect 50258 28478 50260 28530
rect 50092 28476 50260 28478
rect 50204 28466 50260 28476
rect 49980 27682 50036 27692
rect 50092 27972 50148 27982
rect 49868 26910 49870 26962
rect 49922 26910 49924 26962
rect 49868 26898 49924 26910
rect 50092 27298 50148 27916
rect 50204 27970 50260 27982
rect 50204 27918 50206 27970
rect 50258 27918 50260 27970
rect 50204 27860 50260 27918
rect 50204 27524 50260 27804
rect 50204 27458 50260 27468
rect 50092 27246 50094 27298
rect 50146 27246 50148 27298
rect 50092 26964 50148 27246
rect 50316 27188 50372 29484
rect 50316 27122 50372 27132
rect 50428 27074 50484 32398
rect 50540 32004 50596 32510
rect 50540 31938 50596 31948
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50540 31220 50596 31230
rect 50876 31220 50932 33068
rect 50988 33058 51044 33068
rect 51324 33348 51380 33358
rect 51212 32564 51268 32574
rect 51212 32470 51268 32508
rect 50540 31218 50932 31220
rect 50540 31166 50542 31218
rect 50594 31166 50932 31218
rect 50540 31164 50932 31166
rect 51100 32116 51156 32126
rect 51100 31218 51156 32060
rect 51324 32002 51380 33292
rect 51324 31950 51326 32002
rect 51378 31950 51380 32002
rect 51324 31938 51380 31950
rect 51100 31166 51102 31218
rect 51154 31166 51156 31218
rect 50540 31154 50596 31164
rect 51100 31154 51156 31166
rect 51436 31220 51492 37436
rect 51548 37266 51604 37278
rect 51548 37214 51550 37266
rect 51602 37214 51604 37266
rect 51548 37044 51604 37214
rect 51548 36978 51604 36988
rect 51660 36820 51716 38556
rect 51996 38052 52052 38782
rect 51996 37492 52052 37996
rect 52108 38612 52164 39228
rect 52108 38050 52164 38556
rect 52108 37998 52110 38050
rect 52162 37998 52164 38050
rect 52108 37986 52164 37998
rect 52332 39060 52388 41132
rect 52668 41186 52724 41916
rect 52668 41134 52670 41186
rect 52722 41134 52724 41186
rect 52668 41122 52724 41134
rect 52892 41188 52948 41198
rect 52892 41094 52948 41132
rect 52780 40962 52836 40974
rect 52780 40910 52782 40962
rect 52834 40910 52836 40962
rect 52780 40628 52836 40910
rect 52444 40572 52836 40628
rect 52444 40514 52500 40572
rect 52444 40462 52446 40514
rect 52498 40462 52500 40514
rect 52444 40450 52500 40462
rect 52668 39396 52724 39406
rect 52668 39394 52836 39396
rect 52668 39342 52670 39394
rect 52722 39342 52836 39394
rect 52668 39340 52836 39342
rect 52668 39330 52724 39340
rect 52332 39004 52724 39060
rect 52332 37940 52388 39004
rect 52668 38946 52724 39004
rect 52668 38894 52670 38946
rect 52722 38894 52724 38946
rect 52668 38882 52724 38894
rect 52444 38836 52500 38846
rect 52444 38052 52500 38780
rect 52780 38724 52836 39340
rect 53004 38946 53060 42476
rect 53452 42196 53508 42206
rect 53452 42102 53508 42140
rect 53228 41748 53284 41758
rect 53116 40964 53172 40974
rect 53116 40870 53172 40908
rect 53228 40516 53284 41692
rect 53228 40402 53284 40460
rect 53228 40350 53230 40402
rect 53282 40350 53284 40402
rect 53228 40338 53284 40350
rect 53676 41410 53732 44268
rect 53788 43988 53844 45278
rect 53900 45778 53956 45790
rect 53900 45726 53902 45778
rect 53954 45726 53956 45778
rect 53900 44100 53956 45726
rect 54012 45108 54068 45118
rect 54348 45108 54404 46396
rect 54012 45106 54404 45108
rect 54012 45054 54014 45106
rect 54066 45054 54404 45106
rect 54012 45052 54404 45054
rect 54012 44436 54068 45052
rect 54572 44772 54628 48190
rect 54796 48242 54852 48254
rect 54796 48190 54798 48242
rect 54850 48190 54852 48242
rect 54684 48130 54740 48142
rect 54684 48078 54686 48130
rect 54738 48078 54740 48130
rect 54684 45780 54740 48078
rect 54796 47684 54852 48190
rect 54796 47618 54852 47628
rect 54908 47460 54964 48750
rect 55244 48468 55300 49644
rect 55356 49634 55412 49644
rect 55692 49252 55748 49870
rect 55804 49810 55860 50540
rect 55804 49758 55806 49810
rect 55858 49758 55860 49810
rect 55804 49746 55860 49758
rect 55692 49186 55748 49196
rect 55804 49476 55860 49486
rect 55132 48412 55300 48468
rect 55468 49028 55524 49038
rect 55468 48802 55524 48972
rect 55468 48750 55470 48802
rect 55522 48750 55524 48802
rect 55468 48468 55524 48750
rect 55468 48412 55748 48468
rect 54908 47394 54964 47404
rect 55020 48132 55076 48142
rect 55020 47458 55076 48076
rect 55020 47406 55022 47458
rect 55074 47406 55076 47458
rect 55020 47394 55076 47406
rect 55132 47068 55188 48412
rect 55020 47012 55188 47068
rect 55244 48242 55300 48254
rect 55244 48190 55246 48242
rect 55298 48190 55300 48242
rect 55244 47124 55300 48190
rect 55468 48242 55524 48254
rect 55468 48190 55470 48242
rect 55522 48190 55524 48242
rect 55468 47796 55524 48190
rect 55468 47730 55524 47740
rect 55244 47058 55300 47068
rect 55356 47684 55412 47694
rect 54796 46674 54852 46686
rect 54796 46622 54798 46674
rect 54850 46622 54852 46674
rect 54796 46564 54852 46622
rect 54796 46498 54852 46508
rect 55020 46452 55076 47012
rect 55244 46676 55300 46686
rect 55020 46386 55076 46396
rect 55132 46674 55300 46676
rect 55132 46622 55246 46674
rect 55298 46622 55300 46674
rect 55132 46620 55300 46622
rect 54684 45714 54740 45724
rect 54012 44370 54068 44380
rect 54124 44716 54572 44772
rect 54124 44322 54180 44716
rect 54572 44678 54628 44716
rect 54684 45108 54740 45118
rect 54460 44548 54516 44558
rect 54460 44454 54516 44492
rect 54124 44270 54126 44322
rect 54178 44270 54180 44322
rect 54124 44258 54180 44270
rect 53900 44034 53956 44044
rect 54012 44212 54068 44222
rect 53788 43922 53844 43932
rect 54012 43652 54068 44156
rect 53900 43538 53956 43550
rect 53900 43486 53902 43538
rect 53954 43486 53956 43538
rect 53900 43316 53956 43486
rect 53900 43250 53956 43260
rect 53900 43092 53956 43102
rect 53676 41358 53678 41410
rect 53730 41358 53732 41410
rect 53228 40068 53284 40078
rect 53228 39732 53284 40012
rect 53116 39730 53284 39732
rect 53116 39678 53230 39730
rect 53282 39678 53284 39730
rect 53116 39676 53284 39678
rect 53116 39060 53172 39676
rect 53228 39666 53284 39676
rect 53564 39732 53620 39742
rect 53564 39638 53620 39676
rect 53116 38994 53172 39004
rect 53228 39004 53508 39060
rect 53004 38894 53006 38946
rect 53058 38894 53060 38946
rect 53004 38836 53060 38894
rect 53004 38770 53060 38780
rect 52556 38612 52836 38724
rect 52668 38052 52724 38062
rect 52444 38050 52724 38052
rect 52444 37998 52670 38050
rect 52722 37998 52724 38050
rect 52444 37996 52724 37998
rect 52668 37986 52724 37996
rect 52332 37874 52388 37884
rect 52668 37492 52724 37502
rect 51996 37490 52724 37492
rect 51996 37438 52670 37490
rect 52722 37438 52724 37490
rect 51996 37436 52724 37438
rect 52668 37426 52724 37436
rect 51884 37380 51940 37390
rect 51884 37266 51940 37324
rect 51884 37214 51886 37266
rect 51938 37214 51940 37266
rect 51884 37202 51940 37214
rect 52220 37266 52276 37278
rect 52220 37214 52222 37266
rect 52274 37214 52276 37266
rect 51548 36764 51716 36820
rect 51772 37154 51828 37166
rect 51772 37102 51774 37154
rect 51826 37102 51828 37154
rect 51548 33572 51604 36764
rect 51772 36708 51828 37102
rect 51772 36652 51940 36708
rect 51884 36484 51940 36652
rect 52220 36596 52276 37214
rect 52556 37268 52612 37278
rect 52780 37268 52836 38612
rect 52612 37212 52836 37268
rect 52892 38722 52948 38734
rect 52892 38670 52894 38722
rect 52946 38670 52948 38722
rect 52556 37174 52612 37212
rect 52892 37044 52948 38670
rect 53228 38668 53284 39004
rect 53452 38946 53508 39004
rect 53452 38894 53454 38946
rect 53506 38894 53508 38946
rect 53452 38882 53508 38894
rect 52892 36978 52948 36988
rect 53004 38612 53284 38668
rect 53340 38834 53396 38846
rect 53340 38782 53342 38834
rect 53394 38782 53396 38834
rect 53340 38724 53396 38782
rect 52220 36530 52276 36540
rect 52892 36596 52948 36606
rect 51884 36418 51940 36428
rect 52780 36484 52836 36494
rect 51772 36372 51828 36382
rect 51772 35700 51828 36316
rect 52220 36260 52276 36270
rect 52108 36204 52220 36260
rect 51884 35700 51940 35710
rect 51772 35698 51940 35700
rect 51772 35646 51886 35698
rect 51938 35646 51940 35698
rect 51772 35644 51940 35646
rect 51772 35028 51828 35038
rect 51772 34934 51828 34972
rect 51660 34914 51716 34926
rect 51660 34862 51662 34914
rect 51714 34862 51716 34914
rect 51660 34020 51716 34862
rect 51884 34130 51940 35644
rect 51996 35700 52052 35710
rect 51996 35606 52052 35644
rect 52108 35364 52164 36204
rect 52220 36194 52276 36204
rect 52668 35924 52724 35934
rect 51996 35308 52164 35364
rect 52220 35698 52276 35710
rect 52220 35646 52222 35698
rect 52274 35646 52276 35698
rect 51996 34244 52052 35308
rect 52108 34244 52164 34254
rect 51996 34242 52164 34244
rect 51996 34190 52110 34242
rect 52162 34190 52164 34242
rect 51996 34188 52164 34190
rect 52108 34178 52164 34188
rect 51884 34078 51886 34130
rect 51938 34078 51940 34130
rect 51884 34066 51940 34078
rect 51660 33954 51716 33964
rect 51996 34020 52052 34030
rect 51548 33516 51716 33572
rect 51548 33348 51604 33358
rect 51548 33254 51604 33292
rect 51660 32228 51716 33516
rect 51996 32674 52052 33964
rect 51996 32622 51998 32674
rect 52050 32622 52052 32674
rect 51996 32610 52052 32622
rect 52108 33684 52164 33694
rect 51436 31154 51492 31164
rect 51548 32172 51716 32228
rect 51996 32452 52052 32462
rect 51436 30996 51492 31006
rect 51212 30994 51492 30996
rect 51212 30942 51438 30994
rect 51490 30942 51492 30994
rect 51212 30940 51492 30942
rect 51212 30548 51268 30940
rect 51436 30930 51492 30940
rect 50876 30492 51268 30548
rect 50876 30434 50932 30492
rect 50876 30382 50878 30434
rect 50930 30382 50932 30434
rect 50876 30370 50932 30382
rect 51212 30210 51268 30222
rect 51212 30158 51214 30210
rect 51266 30158 51268 30210
rect 50540 29988 50596 29998
rect 50540 29986 50932 29988
rect 50540 29934 50542 29986
rect 50594 29934 50932 29986
rect 50540 29932 50932 29934
rect 50540 29922 50596 29932
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50540 29428 50596 29438
rect 50540 28868 50596 29372
rect 50540 28642 50596 28812
rect 50540 28590 50542 28642
rect 50594 28590 50596 28642
rect 50540 28578 50596 28590
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50764 27860 50820 27870
rect 50540 27188 50596 27198
rect 50540 27094 50596 27132
rect 50428 27022 50430 27074
rect 50482 27022 50484 27074
rect 50428 27010 50484 27022
rect 50764 27074 50820 27804
rect 50876 27412 50932 29932
rect 51212 29540 51268 30158
rect 51212 28868 51268 29484
rect 51324 28868 51380 28878
rect 51212 28866 51380 28868
rect 51212 28814 51326 28866
rect 51378 28814 51380 28866
rect 51212 28812 51380 28814
rect 51324 28802 51380 28812
rect 50988 28644 51044 28654
rect 51548 28644 51604 32172
rect 50988 28550 51044 28588
rect 51212 28588 51604 28644
rect 51660 32004 51716 32014
rect 50876 27346 50932 27356
rect 50764 27022 50766 27074
rect 50818 27022 50820 27074
rect 50764 27010 50820 27022
rect 50988 27076 51044 27086
rect 50988 26982 51044 27020
rect 50092 26898 50148 26908
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 49756 26462 49758 26514
rect 49810 26462 49812 26514
rect 49756 26450 49812 26462
rect 50092 26404 50148 26414
rect 50092 26310 50148 26348
rect 49644 26292 49700 26302
rect 49644 26198 49700 26236
rect 49868 26290 49924 26302
rect 49868 26238 49870 26290
rect 49922 26238 49924 26290
rect 49868 25844 49924 26238
rect 50988 26290 51044 26302
rect 50988 26238 50990 26290
rect 51042 26238 51044 26290
rect 49868 25778 49924 25788
rect 50540 25844 50596 25854
rect 50540 25620 50596 25788
rect 50988 25732 51044 26238
rect 50988 25666 51044 25676
rect 50540 25564 50708 25620
rect 50092 25508 50148 25518
rect 49756 25284 49812 25294
rect 49756 25190 49812 25228
rect 49868 25282 49924 25294
rect 49868 25230 49870 25282
rect 49922 25230 49924 25282
rect 49308 24894 49310 24946
rect 49362 24894 49364 24946
rect 49308 23826 49364 24894
rect 49420 24892 49588 24948
rect 49420 24164 49476 24892
rect 49868 24836 49924 25230
rect 49868 24770 49924 24780
rect 50092 25282 50148 25452
rect 50316 25396 50372 25406
rect 50092 25230 50094 25282
rect 50146 25230 50148 25282
rect 50092 24836 50148 25230
rect 50204 25394 50372 25396
rect 50204 25342 50318 25394
rect 50370 25342 50372 25394
rect 50204 25340 50372 25342
rect 50204 25060 50260 25340
rect 50316 25330 50372 25340
rect 50540 25396 50596 25406
rect 50540 25302 50596 25340
rect 50652 25394 50708 25564
rect 50876 25508 50932 25518
rect 50876 25414 50932 25452
rect 50652 25342 50654 25394
rect 50706 25342 50708 25394
rect 50652 25330 50708 25342
rect 51100 25394 51156 25406
rect 51100 25342 51102 25394
rect 51154 25342 51156 25394
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50204 24994 50260 25004
rect 50540 24948 50596 24958
rect 50092 24770 50148 24780
rect 50316 24892 50540 24948
rect 49532 24724 49588 24734
rect 49532 24630 49588 24668
rect 49756 24724 49812 24734
rect 49756 24630 49812 24668
rect 49644 24610 49700 24622
rect 49644 24558 49646 24610
rect 49698 24558 49700 24610
rect 49420 24108 49588 24164
rect 49308 23774 49310 23826
rect 49362 23774 49364 23826
rect 49308 23762 49364 23774
rect 49420 23938 49476 23950
rect 49420 23886 49422 23938
rect 49474 23886 49476 23938
rect 49420 23828 49476 23886
rect 49308 22370 49364 22382
rect 49308 22318 49310 22370
rect 49362 22318 49364 22370
rect 49308 22260 49364 22318
rect 49308 22194 49364 22204
rect 49308 21698 49364 21710
rect 49308 21646 49310 21698
rect 49362 21646 49364 21698
rect 49308 21364 49364 21646
rect 49420 21700 49476 23772
rect 49420 21634 49476 21644
rect 49532 21588 49588 24108
rect 49644 24052 49700 24558
rect 50204 24500 50260 24510
rect 49644 23986 49700 23996
rect 49868 24498 50260 24500
rect 49868 24446 50206 24498
rect 50258 24446 50260 24498
rect 49868 24444 50260 24446
rect 49644 23828 49700 23838
rect 49644 23266 49700 23772
rect 49644 23214 49646 23266
rect 49698 23214 49700 23266
rect 49644 23202 49700 23214
rect 49868 23156 49924 24444
rect 50204 24434 50260 24444
rect 49980 23828 50036 23838
rect 49980 23826 50148 23828
rect 49980 23774 49982 23826
rect 50034 23774 50148 23826
rect 49980 23772 50148 23774
rect 49980 23762 50036 23772
rect 49868 23062 49924 23100
rect 49980 22596 50036 22606
rect 49980 22502 50036 22540
rect 49756 22370 49812 22382
rect 49756 22318 49758 22370
rect 49810 22318 49812 22370
rect 49532 21522 49588 21532
rect 49644 21700 49700 21710
rect 49308 21298 49364 21308
rect 49644 21252 49700 21644
rect 49644 21186 49700 21196
rect 49532 20916 49588 20926
rect 49532 20822 49588 20860
rect 49308 20020 49364 20030
rect 49308 19926 49364 19964
rect 49196 19404 49364 19460
rect 49084 19170 49140 19180
rect 48916 18396 49028 18452
rect 48860 18338 48916 18396
rect 48860 18286 48862 18338
rect 48914 18286 48916 18338
rect 48860 18274 48916 18286
rect 48636 17826 48692 17836
rect 49084 17668 49140 17678
rect 49084 17574 49140 17612
rect 49308 17668 49364 19404
rect 49420 18900 49476 18910
rect 49420 18562 49476 18844
rect 49644 18676 49700 18686
rect 49420 18510 49422 18562
rect 49474 18510 49476 18562
rect 49420 18498 49476 18510
rect 49532 18564 49588 18574
rect 49644 18564 49700 18620
rect 49532 18562 49700 18564
rect 49532 18510 49534 18562
rect 49586 18510 49700 18562
rect 49532 18508 49700 18510
rect 49532 18498 49588 18508
rect 49756 18450 49812 22318
rect 49868 21586 49924 21598
rect 49868 21534 49870 21586
rect 49922 21534 49924 21586
rect 49868 20916 49924 21534
rect 49980 21476 50036 21486
rect 49980 21382 50036 21420
rect 50092 21140 50148 23772
rect 50316 23548 50372 24892
rect 50540 24882 50596 24892
rect 50988 24722 51044 24734
rect 50988 24670 50990 24722
rect 51042 24670 51044 24722
rect 50540 24500 50596 24510
rect 50540 24164 50596 24444
rect 50988 24500 51044 24670
rect 50988 24434 51044 24444
rect 50540 24098 50596 24108
rect 50652 24276 50708 24286
rect 50652 23938 50708 24220
rect 50652 23886 50654 23938
rect 50706 23886 50708 23938
rect 50652 23874 50708 23886
rect 51100 23940 51156 25342
rect 51100 23846 51156 23884
rect 50876 23828 50932 23838
rect 50876 23734 50932 23772
rect 50092 21074 50148 21084
rect 50204 23492 50372 23548
rect 50428 23716 50484 23726
rect 49868 20850 49924 20860
rect 50204 20692 50260 23492
rect 50204 20626 50260 20636
rect 50204 18676 50260 18686
rect 50428 18676 50484 23660
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50540 23156 50596 23166
rect 50540 22370 50596 23100
rect 50540 22318 50542 22370
rect 50594 22318 50596 22370
rect 50540 22306 50596 22318
rect 51100 22594 51156 22606
rect 51100 22542 51102 22594
rect 51154 22542 51156 22594
rect 51100 22372 51156 22542
rect 51100 22306 51156 22316
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 51212 20916 51268 28588
rect 51548 27860 51604 27870
rect 51660 27860 51716 31948
rect 51996 31890 52052 32396
rect 52108 32002 52164 33628
rect 52220 32788 52276 35646
rect 52332 35476 52388 35486
rect 52332 34130 52388 35420
rect 52332 34078 52334 34130
rect 52386 34078 52388 34130
rect 52332 34066 52388 34078
rect 52220 32722 52276 32732
rect 52108 31950 52110 32002
rect 52162 31950 52164 32002
rect 52108 31938 52164 31950
rect 52220 32004 52276 32014
rect 51996 31838 51998 31890
rect 52050 31838 52052 31890
rect 51996 31826 52052 31838
rect 51772 31106 51828 31118
rect 51772 31054 51774 31106
rect 51826 31054 51828 31106
rect 51772 30996 51828 31054
rect 51772 30930 51828 30940
rect 52108 30994 52164 31006
rect 52108 30942 52110 30994
rect 52162 30942 52164 30994
rect 51884 30212 51940 30222
rect 51884 30118 51940 30156
rect 51996 30098 52052 30110
rect 51996 30046 51998 30098
rect 52050 30046 52052 30098
rect 51996 29316 52052 30046
rect 52108 29428 52164 30942
rect 52108 29362 52164 29372
rect 52220 29316 52276 31948
rect 52668 31892 52724 35868
rect 52780 35588 52836 36428
rect 52780 35522 52836 35532
rect 52892 36482 52948 36540
rect 52892 36430 52894 36482
rect 52946 36430 52948 36482
rect 52892 35700 52948 36430
rect 53004 35924 53060 38612
rect 53228 38050 53284 38062
rect 53228 37998 53230 38050
rect 53282 37998 53284 38050
rect 53228 36820 53284 37998
rect 53340 36932 53396 38668
rect 53452 38612 53508 38622
rect 53452 38610 53620 38612
rect 53452 38558 53454 38610
rect 53506 38558 53620 38610
rect 53452 38556 53620 38558
rect 53452 38546 53508 38556
rect 53340 36866 53396 36876
rect 53452 37938 53508 37950
rect 53452 37886 53454 37938
rect 53506 37886 53508 37938
rect 53228 36754 53284 36764
rect 53116 36484 53172 36494
rect 53116 36390 53172 36428
rect 53228 36370 53284 36382
rect 53228 36318 53230 36370
rect 53282 36318 53284 36370
rect 53228 36260 53284 36318
rect 53004 35858 53060 35868
rect 53116 36148 53172 36158
rect 52780 33346 52836 33358
rect 52780 33294 52782 33346
rect 52834 33294 52836 33346
rect 52780 33236 52836 33294
rect 52892 33348 52948 35644
rect 53004 35140 53060 35150
rect 53116 35140 53172 36092
rect 53228 35698 53284 36204
rect 53228 35646 53230 35698
rect 53282 35646 53284 35698
rect 53228 35634 53284 35646
rect 53340 35810 53396 35822
rect 53340 35758 53342 35810
rect 53394 35758 53396 35810
rect 53340 35700 53396 35758
rect 53340 35634 53396 35644
rect 53060 35084 53172 35140
rect 53004 35046 53060 35084
rect 53452 35028 53508 37886
rect 53564 37266 53620 38556
rect 53564 37214 53566 37266
rect 53618 37214 53620 37266
rect 53564 37202 53620 37214
rect 53676 36484 53732 41358
rect 53788 42980 53844 42990
rect 53788 41186 53844 42924
rect 53900 41970 53956 43036
rect 54012 42082 54068 43596
rect 54236 43876 54292 43886
rect 54236 43650 54292 43820
rect 54236 43598 54238 43650
rect 54290 43598 54292 43650
rect 54236 43586 54292 43598
rect 54348 43764 54404 43774
rect 54012 42030 54014 42082
rect 54066 42030 54068 42082
rect 54012 42018 54068 42030
rect 54236 42196 54292 42206
rect 53900 41918 53902 41970
rect 53954 41918 53956 41970
rect 53900 41906 53956 41918
rect 54236 41410 54292 42140
rect 54236 41358 54238 41410
rect 54290 41358 54292 41410
rect 54236 41346 54292 41358
rect 54348 41412 54404 43708
rect 54572 42868 54628 42878
rect 54572 42754 54628 42812
rect 54572 42702 54574 42754
rect 54626 42702 54628 42754
rect 54572 42690 54628 42702
rect 54460 41412 54516 41422
rect 54348 41410 54516 41412
rect 54348 41358 54462 41410
rect 54514 41358 54516 41410
rect 54348 41356 54516 41358
rect 54460 41346 54516 41356
rect 54684 41300 54740 45052
rect 54796 45106 54852 45118
rect 54796 45054 54798 45106
rect 54850 45054 54852 45106
rect 54796 44324 54852 45054
rect 55132 45108 55188 46620
rect 55244 46610 55300 46620
rect 55132 45042 55188 45052
rect 55244 46452 55300 46462
rect 55244 44994 55300 46396
rect 55244 44942 55246 44994
rect 55298 44942 55300 44994
rect 55244 44930 55300 44942
rect 54908 44324 54964 44334
rect 55356 44324 55412 47628
rect 55468 47460 55524 47470
rect 55468 46002 55524 47404
rect 55468 45950 55470 46002
rect 55522 45950 55524 46002
rect 55468 45938 55524 45950
rect 55580 46788 55636 46798
rect 55580 46228 55636 46732
rect 55692 46674 55748 48412
rect 55804 47346 55860 49420
rect 55804 47294 55806 47346
rect 55858 47294 55860 47346
rect 55804 47282 55860 47294
rect 56028 48018 56084 48030
rect 56028 47966 56030 48018
rect 56082 47966 56084 48018
rect 56028 47796 56084 47966
rect 56028 47068 56084 47740
rect 56252 47124 56308 53116
rect 56812 52946 56868 55356
rect 56924 55076 56980 55086
rect 56924 53954 56980 55020
rect 56924 53902 56926 53954
rect 56978 53902 56980 53954
rect 56924 53844 56980 53902
rect 56924 53778 56980 53788
rect 56812 52894 56814 52946
rect 56866 52894 56868 52946
rect 56812 52882 56868 52894
rect 56588 52836 56644 52846
rect 56588 52742 56644 52780
rect 57148 52724 57204 52734
rect 57148 52630 57204 52668
rect 57036 51492 57092 51502
rect 57036 51378 57092 51436
rect 57036 51326 57038 51378
rect 57090 51326 57092 51378
rect 56700 51266 56756 51278
rect 56700 51214 56702 51266
rect 56754 51214 56756 51266
rect 56700 50260 56756 51214
rect 57036 50932 57092 51326
rect 57036 50866 57092 50876
rect 57260 50820 57316 55580
rect 58156 55300 58212 56140
rect 58156 55206 58212 55244
rect 58268 56082 58324 56364
rect 58380 56308 58436 56318
rect 58380 56214 58436 56252
rect 58268 56030 58270 56082
rect 58322 56030 58324 56082
rect 57596 54852 57652 54862
rect 57484 53060 57540 53070
rect 57484 52966 57540 53004
rect 57596 52164 57652 54796
rect 57932 54292 57988 54302
rect 58268 54292 58324 56030
rect 58716 55188 58772 55198
rect 58772 55132 58884 55188
rect 58716 55094 58772 55132
rect 57932 54290 58324 54292
rect 57932 54238 57934 54290
rect 57986 54238 58324 54290
rect 57932 54236 58324 54238
rect 58380 55074 58436 55086
rect 58380 55022 58382 55074
rect 58434 55022 58436 55074
rect 57708 53956 57764 53994
rect 57708 53890 57764 53900
rect 57932 53508 57988 54236
rect 58156 53842 58212 53854
rect 58156 53790 58158 53842
rect 58210 53790 58212 53842
rect 57932 53442 57988 53452
rect 58044 53732 58100 53742
rect 57820 52946 57876 52958
rect 57820 52894 57822 52946
rect 57874 52894 57876 52946
rect 57708 52164 57764 52174
rect 57596 52162 57764 52164
rect 57596 52110 57710 52162
rect 57762 52110 57764 52162
rect 57596 52108 57764 52110
rect 57708 52098 57764 52108
rect 57820 51604 57876 52894
rect 58044 52164 58100 53676
rect 58156 52276 58212 53790
rect 58380 53730 58436 55022
rect 58380 53678 58382 53730
rect 58434 53678 58436 53730
rect 58380 53666 58436 53678
rect 58492 55074 58548 55086
rect 58492 55022 58494 55074
rect 58546 55022 58548 55074
rect 58492 53732 58548 55022
rect 58492 53666 58548 53676
rect 58828 53058 58884 55132
rect 58940 55186 58996 55198
rect 58940 55134 58942 55186
rect 58994 55134 58996 55186
rect 58940 53844 58996 55134
rect 59164 55188 59220 56700
rect 59276 56308 59332 56318
rect 59276 56214 59332 56252
rect 62748 55300 62804 55310
rect 59276 55188 59332 55198
rect 59388 55188 59444 55198
rect 59164 55186 59388 55188
rect 59164 55134 59278 55186
rect 59330 55134 59388 55186
rect 59164 55132 59388 55134
rect 59276 55122 59332 55132
rect 59388 54738 59444 55132
rect 59612 55188 59668 55198
rect 61068 55188 61124 55198
rect 59612 55186 60004 55188
rect 59612 55134 59614 55186
rect 59666 55134 60004 55186
rect 59612 55132 60004 55134
rect 59612 55122 59668 55132
rect 59388 54686 59390 54738
rect 59442 54686 59444 54738
rect 59388 54674 59444 54686
rect 58940 53508 58996 53788
rect 59052 53732 59108 53742
rect 59052 53638 59108 53676
rect 59612 53508 59668 53518
rect 58940 53452 59108 53508
rect 58828 53006 58830 53058
rect 58882 53006 58884 53058
rect 58828 52994 58884 53006
rect 59052 52946 59108 53452
rect 59052 52894 59054 52946
rect 59106 52894 59108 52946
rect 59052 52882 59108 52894
rect 59612 52946 59668 53452
rect 59612 52894 59614 52946
rect 59666 52894 59668 52946
rect 59612 52882 59668 52894
rect 58380 52834 58436 52846
rect 58380 52782 58382 52834
rect 58434 52782 58436 52834
rect 58268 52276 58324 52286
rect 58156 52274 58324 52276
rect 58156 52222 58270 52274
rect 58322 52222 58324 52274
rect 58156 52220 58324 52222
rect 58044 52108 58212 52164
rect 57708 51548 57876 51604
rect 57260 50754 57316 50764
rect 57484 51492 57540 51502
rect 57036 50708 57092 50718
rect 56924 50484 56980 50522
rect 56588 50036 56644 50046
rect 56588 49942 56644 49980
rect 56700 48916 56756 50204
rect 56700 48850 56756 48860
rect 56812 50428 56924 50484
rect 56812 48914 56868 50428
rect 56924 50418 56980 50428
rect 56924 49812 56980 49822
rect 56924 49718 56980 49756
rect 56812 48862 56814 48914
rect 56866 48862 56868 48914
rect 56812 48850 56868 48862
rect 56364 48804 56420 48814
rect 56364 47458 56420 48748
rect 57036 48692 57092 50652
rect 57484 50148 57540 51436
rect 57708 51156 57764 51548
rect 57820 51268 57876 51278
rect 57820 51174 57876 51212
rect 57708 51090 57764 51100
rect 57932 51156 57988 51166
rect 57484 50082 57540 50092
rect 57820 50370 57876 50382
rect 57820 50318 57822 50370
rect 57874 50318 57876 50370
rect 57148 49924 57204 49934
rect 57148 49810 57204 49868
rect 57148 49758 57150 49810
rect 57202 49758 57204 49810
rect 57148 49140 57204 49758
rect 57484 49700 57540 49710
rect 57148 49074 57204 49084
rect 57260 49698 57540 49700
rect 57260 49646 57486 49698
rect 57538 49646 57540 49698
rect 57260 49644 57540 49646
rect 57036 48626 57092 48636
rect 56700 48468 56756 48478
rect 56700 48374 56756 48412
rect 57036 48356 57092 48366
rect 56924 47908 56980 47918
rect 56364 47406 56366 47458
rect 56418 47406 56420 47458
rect 56364 47394 56420 47406
rect 56812 47852 56924 47908
rect 56812 47458 56868 47852
rect 56924 47842 56980 47852
rect 56812 47406 56814 47458
rect 56866 47406 56868 47458
rect 56812 47394 56868 47406
rect 56028 47012 56196 47068
rect 55692 46622 55694 46674
rect 55746 46622 55748 46674
rect 55692 46610 55748 46622
rect 55580 45890 55636 46172
rect 55580 45838 55582 45890
rect 55634 45838 55636 45890
rect 55580 45826 55636 45838
rect 55692 46114 55748 46126
rect 55692 46062 55694 46114
rect 55746 46062 55748 46114
rect 55692 45444 55748 46062
rect 54796 44268 54908 44324
rect 54908 44258 54964 44268
rect 55020 44322 55412 44324
rect 55020 44270 55358 44322
rect 55410 44270 55412 44322
rect 55020 44268 55412 44270
rect 54796 43876 54852 43886
rect 54796 41970 54852 43820
rect 55020 43540 55076 44268
rect 55356 44258 55412 44268
rect 55468 45388 55748 45444
rect 55356 43988 55412 43998
rect 55020 43446 55076 43484
rect 55244 43538 55300 43550
rect 55244 43486 55246 43538
rect 55298 43486 55300 43538
rect 54796 41918 54798 41970
rect 54850 41918 54852 41970
rect 54796 41524 54852 41918
rect 54908 42194 54964 42206
rect 54908 42142 54910 42194
rect 54962 42142 54964 42194
rect 54908 41636 54964 42142
rect 55244 41636 55300 43486
rect 55356 41970 55412 43932
rect 55356 41918 55358 41970
rect 55410 41918 55412 41970
rect 55356 41860 55412 41918
rect 55356 41794 55412 41804
rect 54908 41580 55300 41636
rect 54796 41468 55188 41524
rect 54796 41300 54852 41310
rect 54684 41298 54852 41300
rect 54684 41246 54798 41298
rect 54850 41246 54852 41298
rect 54684 41244 54852 41246
rect 54796 41234 54852 41244
rect 53788 41134 53790 41186
rect 53842 41134 53844 41186
rect 53788 41122 53844 41134
rect 54572 41188 54628 41198
rect 54572 40962 54628 41132
rect 54572 40910 54574 40962
rect 54626 40910 54628 40962
rect 54572 40898 54628 40910
rect 55132 40852 55188 41468
rect 55132 40786 55188 40796
rect 54572 40740 54628 40750
rect 54236 40516 54292 40526
rect 54236 40422 54292 40460
rect 54572 40514 54628 40684
rect 54572 40462 54574 40514
rect 54626 40462 54628 40514
rect 53788 40292 53844 40302
rect 53788 39730 53844 40236
rect 53788 39678 53790 39730
rect 53842 39678 53844 39730
rect 53788 39666 53844 39678
rect 54348 40180 54404 40190
rect 53788 38836 53844 38846
rect 53788 38050 53844 38780
rect 53788 37998 53790 38050
rect 53842 37998 53844 38050
rect 53788 37986 53844 37998
rect 53900 37940 53956 37950
rect 53900 37846 53956 37884
rect 54012 37492 54068 37502
rect 54012 37398 54068 37436
rect 54236 37268 54292 37278
rect 54236 37174 54292 37212
rect 54124 37156 54180 37166
rect 54124 37062 54180 37100
rect 54012 37044 54068 37054
rect 53788 36820 53844 36830
rect 53844 36764 53956 36820
rect 53788 36754 53844 36764
rect 53564 36428 53732 36484
rect 53564 36148 53620 36428
rect 53564 36082 53620 36092
rect 53676 36258 53732 36270
rect 53676 36206 53678 36258
rect 53730 36206 53732 36258
rect 53564 35586 53620 35598
rect 53564 35534 53566 35586
rect 53618 35534 53620 35586
rect 53564 35140 53620 35534
rect 53564 35046 53620 35084
rect 53116 34972 53452 35028
rect 53116 33570 53172 34972
rect 53452 34962 53508 34972
rect 53676 34916 53732 36206
rect 53788 35252 53844 35262
rect 53788 35138 53844 35196
rect 53788 35086 53790 35138
rect 53842 35086 53844 35138
rect 53788 35074 53844 35086
rect 53676 34850 53732 34860
rect 53228 34802 53284 34814
rect 53228 34750 53230 34802
rect 53282 34750 53284 34802
rect 53228 33684 53284 34750
rect 53340 34802 53396 34814
rect 53340 34750 53342 34802
rect 53394 34750 53396 34802
rect 53340 34130 53396 34750
rect 53900 34356 53956 36764
rect 54012 36708 54068 36988
rect 54012 36652 54180 36708
rect 54012 36484 54068 36494
rect 54012 36390 54068 36428
rect 54012 35588 54068 35598
rect 54012 35494 54068 35532
rect 54124 34916 54180 36652
rect 54348 35700 54404 40124
rect 54572 39284 54628 40462
rect 54684 40404 54740 40414
rect 54684 39506 54740 40348
rect 55132 40402 55188 40414
rect 55132 40350 55134 40402
rect 55186 40350 55188 40402
rect 54796 40180 54852 40190
rect 55132 40180 55188 40350
rect 54796 40178 54964 40180
rect 54796 40126 54798 40178
rect 54850 40126 54964 40178
rect 54796 40124 54964 40126
rect 54796 40114 54852 40124
rect 54684 39454 54686 39506
rect 54738 39454 54740 39506
rect 54684 39442 54740 39454
rect 54796 39956 54852 39966
rect 54908 39956 54964 40124
rect 55132 40114 55188 40124
rect 54908 39900 55188 39956
rect 54796 39506 54852 39900
rect 54796 39454 54798 39506
rect 54850 39454 54852 39506
rect 54796 39442 54852 39454
rect 54908 39394 54964 39406
rect 54908 39342 54910 39394
rect 54962 39342 54964 39394
rect 54908 39284 54964 39342
rect 54572 39228 54964 39284
rect 54796 38946 54852 38958
rect 54796 38894 54798 38946
rect 54850 38894 54852 38946
rect 54796 38612 54852 38894
rect 54796 38546 54852 38556
rect 54796 38050 54852 38062
rect 54796 37998 54798 38050
rect 54850 37998 54852 38050
rect 54796 37716 54852 37998
rect 54908 38052 54964 39228
rect 54908 37986 54964 37996
rect 55020 39394 55076 39406
rect 55020 39342 55022 39394
rect 55074 39342 55076 39394
rect 55020 37940 55076 39342
rect 55020 37874 55076 37884
rect 55132 39394 55188 39900
rect 55244 39620 55300 41580
rect 55356 41300 55412 41310
rect 55468 41300 55524 45388
rect 55916 45220 55972 45230
rect 55916 45126 55972 45164
rect 55580 45106 55636 45118
rect 55580 45054 55582 45106
rect 55634 45054 55636 45106
rect 55580 44996 55636 45054
rect 55580 44930 55636 44940
rect 55916 44996 55972 45006
rect 55916 44902 55972 44940
rect 55916 44436 55972 44446
rect 55692 44380 55916 44436
rect 55580 44100 55636 44110
rect 55580 43650 55636 44044
rect 55580 43598 55582 43650
rect 55634 43598 55636 43650
rect 55580 43586 55636 43598
rect 55468 41244 55636 41300
rect 55356 41074 55412 41244
rect 55356 41022 55358 41074
rect 55410 41022 55412 41074
rect 55356 39844 55412 41022
rect 55468 40964 55524 40974
rect 55468 40626 55524 40908
rect 55468 40574 55470 40626
rect 55522 40574 55524 40626
rect 55468 40562 55524 40574
rect 55580 39956 55636 41244
rect 55692 40740 55748 44380
rect 55916 44370 55972 44380
rect 56140 44324 56196 47012
rect 56028 44322 56196 44324
rect 56028 44270 56142 44322
rect 56194 44270 56196 44322
rect 56028 44268 56196 44270
rect 55804 43652 55860 43662
rect 55804 43558 55860 43596
rect 55916 43538 55972 43550
rect 55916 43486 55918 43538
rect 55970 43486 55972 43538
rect 55916 43092 55972 43486
rect 55916 43026 55972 43036
rect 56028 42868 56084 44268
rect 56140 44258 56196 44268
rect 56252 44212 56308 47068
rect 56700 47348 56756 47358
rect 56700 47012 56756 47292
rect 56924 47346 56980 47358
rect 56924 47294 56926 47346
rect 56978 47294 56980 47346
rect 56700 46956 56868 47012
rect 56700 46788 56756 46798
rect 56588 46786 56756 46788
rect 56588 46734 56702 46786
rect 56754 46734 56756 46786
rect 56588 46732 56756 46734
rect 56476 45890 56532 45902
rect 56476 45838 56478 45890
rect 56530 45838 56532 45890
rect 56476 44436 56532 45838
rect 56588 44660 56644 46732
rect 56700 46722 56756 46732
rect 56812 46786 56868 46956
rect 56812 46734 56814 46786
rect 56866 46734 56868 46786
rect 56812 46722 56868 46734
rect 56588 44594 56644 44604
rect 56700 46450 56756 46462
rect 56700 46398 56702 46450
rect 56754 46398 56756 46450
rect 56476 44370 56532 44380
rect 56252 44146 56308 44156
rect 56700 43876 56756 46398
rect 56924 45556 56980 47294
rect 57036 45778 57092 48300
rect 57036 45726 57038 45778
rect 57090 45726 57092 45778
rect 57036 45714 57092 45726
rect 57148 48242 57204 48254
rect 57148 48190 57150 48242
rect 57202 48190 57204 48242
rect 57148 45556 57204 48190
rect 57260 46788 57316 49644
rect 57484 49634 57540 49644
rect 57820 49588 57876 50318
rect 57932 49700 57988 51100
rect 58044 50596 58100 50606
rect 58044 50502 58100 50540
rect 57932 49634 57988 49644
rect 58044 49810 58100 49822
rect 58044 49758 58046 49810
rect 58098 49758 58100 49810
rect 57820 49522 57876 49532
rect 58044 49364 58100 49758
rect 57484 49252 57540 49262
rect 57260 46722 57316 46732
rect 57372 48018 57428 48030
rect 57372 47966 57374 48018
rect 57426 47966 57428 48018
rect 57260 46564 57316 46574
rect 57372 46564 57428 47966
rect 57484 46786 57540 49196
rect 57820 48802 57876 48814
rect 57820 48750 57822 48802
rect 57874 48750 57876 48802
rect 57820 48356 57876 48750
rect 57820 48290 57876 48300
rect 57708 48242 57764 48254
rect 57708 48190 57710 48242
rect 57762 48190 57764 48242
rect 57484 46734 57486 46786
rect 57538 46734 57540 46786
rect 57484 46722 57540 46734
rect 57596 47458 57652 47470
rect 57596 47406 57598 47458
rect 57650 47406 57652 47458
rect 57596 46788 57652 47406
rect 57596 46722 57652 46732
rect 57708 47124 57764 48190
rect 57932 48244 57988 48254
rect 57932 48150 57988 48188
rect 57260 46562 57428 46564
rect 57260 46510 57262 46562
rect 57314 46510 57428 46562
rect 57260 46508 57428 46510
rect 57260 46452 57316 46508
rect 57260 46386 57316 46396
rect 56924 45500 57092 45556
rect 57148 45500 57428 45556
rect 57036 45444 57092 45500
rect 57036 45388 57204 45444
rect 56924 45332 56980 45342
rect 56924 45218 56980 45276
rect 56924 45166 56926 45218
rect 56978 45166 56980 45218
rect 56924 45154 56980 45166
rect 57036 44324 57092 44334
rect 56812 44212 56868 44222
rect 56812 44118 56868 44156
rect 56700 43810 56756 43820
rect 56700 43652 56756 43662
rect 56588 43650 56756 43652
rect 56588 43598 56702 43650
rect 56754 43598 56756 43650
rect 56588 43596 56756 43598
rect 56476 43538 56532 43550
rect 56476 43486 56478 43538
rect 56530 43486 56532 43538
rect 56476 43428 56532 43486
rect 56028 42802 56084 42812
rect 56140 43372 56532 43428
rect 55916 42756 55972 42766
rect 55916 42662 55972 42700
rect 55916 41970 55972 41982
rect 55916 41918 55918 41970
rect 55970 41918 55972 41970
rect 55692 40674 55748 40684
rect 55804 41412 55860 41422
rect 55692 40514 55748 40526
rect 55692 40462 55694 40514
rect 55746 40462 55748 40514
rect 55692 39956 55748 40462
rect 55804 40516 55860 41356
rect 55916 41300 55972 41918
rect 55916 41234 55972 41244
rect 56028 41186 56084 41198
rect 56028 41134 56030 41186
rect 56082 41134 56084 41186
rect 55916 41076 55972 41086
rect 55916 40982 55972 41020
rect 55804 40422 55860 40460
rect 56028 40292 56084 41134
rect 55916 39956 55972 39966
rect 55692 39900 55916 39956
rect 55356 39788 55524 39844
rect 55356 39620 55412 39630
rect 55244 39564 55356 39620
rect 55356 39554 55412 39564
rect 55468 39396 55524 39788
rect 55580 39508 55636 39900
rect 55916 39890 55972 39900
rect 55580 39442 55636 39452
rect 55132 39342 55134 39394
rect 55186 39342 55188 39394
rect 55132 37716 55188 39342
rect 54796 37660 55188 37716
rect 55244 39340 55524 39396
rect 54908 37266 54964 37278
rect 54908 37214 54910 37266
rect 54962 37214 54964 37266
rect 54908 36708 54964 37214
rect 54908 36642 54964 36652
rect 54348 35634 54404 35644
rect 54460 36482 54516 36494
rect 54460 36430 54462 36482
rect 54514 36430 54516 36482
rect 54460 35698 54516 36430
rect 54796 36372 54852 36382
rect 54796 36278 54852 36316
rect 54460 35646 54462 35698
rect 54514 35646 54516 35698
rect 54460 35476 54516 35646
rect 54460 35410 54516 35420
rect 54796 35364 54852 35374
rect 55020 35308 55076 37660
rect 55244 37268 55300 39340
rect 55916 38836 55972 38846
rect 55916 38742 55972 38780
rect 55804 38276 55860 38286
rect 55804 37378 55860 38220
rect 55916 38052 55972 38062
rect 55916 37958 55972 37996
rect 55804 37326 55806 37378
rect 55858 37326 55860 37378
rect 55804 37314 55860 37326
rect 55132 37212 55300 37268
rect 56028 37266 56084 40236
rect 56140 39618 56196 43372
rect 56364 42980 56420 42990
rect 56364 42886 56420 42924
rect 56476 42868 56532 42878
rect 56476 42774 56532 42812
rect 56140 39566 56142 39618
rect 56194 39566 56196 39618
rect 56140 39554 56196 39566
rect 56252 41860 56308 41870
rect 56252 38668 56308 41804
rect 56476 41412 56532 41422
rect 56476 41318 56532 41356
rect 56364 41074 56420 41086
rect 56364 41022 56366 41074
rect 56418 41022 56420 41074
rect 56364 40404 56420 41022
rect 56476 41076 56532 41086
rect 56588 41076 56644 43596
rect 56700 43586 56756 43596
rect 56812 43540 56868 43550
rect 56812 43538 56980 43540
rect 56812 43486 56814 43538
rect 56866 43486 56980 43538
rect 56812 43484 56980 43486
rect 56812 43474 56868 43484
rect 56476 41074 56644 41076
rect 56476 41022 56478 41074
rect 56530 41022 56644 41074
rect 56476 41020 56644 41022
rect 56476 41010 56532 41020
rect 56588 40964 56644 41020
rect 56588 40898 56644 40908
rect 56812 41412 56868 41422
rect 56364 40338 56420 40348
rect 56700 40516 56756 40526
rect 56028 37214 56030 37266
rect 56082 37214 56084 37266
rect 55132 36708 55188 37212
rect 56028 37202 56084 37214
rect 56140 38612 56308 38668
rect 56364 39844 56420 39854
rect 56364 39506 56420 39788
rect 56364 39454 56366 39506
rect 56418 39454 56420 39506
rect 55356 37156 55412 37166
rect 55132 36642 55188 36652
rect 55244 37154 55412 37156
rect 55244 37102 55358 37154
rect 55410 37102 55412 37154
rect 55244 37100 55412 37102
rect 54236 34916 54292 34926
rect 54124 34914 54292 34916
rect 54124 34862 54238 34914
rect 54290 34862 54292 34914
rect 54124 34860 54292 34862
rect 54236 34850 54292 34860
rect 54572 34916 54628 34926
rect 54572 34802 54628 34860
rect 54572 34750 54574 34802
rect 54626 34750 54628 34802
rect 54572 34738 54628 34750
rect 54684 34802 54740 34814
rect 54684 34750 54686 34802
rect 54738 34750 54740 34802
rect 54348 34690 54404 34702
rect 54348 34638 54350 34690
rect 54402 34638 54404 34690
rect 54348 34580 54404 34638
rect 54348 34514 54404 34524
rect 54460 34690 54516 34702
rect 54460 34638 54462 34690
rect 54514 34638 54516 34690
rect 54460 34356 54516 34638
rect 54684 34356 54740 34750
rect 53900 34300 54180 34356
rect 53340 34078 53342 34130
rect 53394 34078 53396 34130
rect 53340 34066 53396 34078
rect 53788 34132 53844 34142
rect 53788 34038 53844 34076
rect 54012 34132 54068 34142
rect 54012 34038 54068 34076
rect 53228 33618 53284 33628
rect 53564 34018 53620 34030
rect 53564 33966 53566 34018
rect 53618 33966 53620 34018
rect 53116 33518 53118 33570
rect 53170 33518 53172 33570
rect 53116 33506 53172 33518
rect 53452 33460 53508 33470
rect 53564 33460 53620 33966
rect 53900 34020 53956 34030
rect 53900 33926 53956 33964
rect 54124 33572 54180 34300
rect 54348 34300 54516 34356
rect 54572 34300 54740 34356
rect 54348 34244 54404 34300
rect 53452 33458 53620 33460
rect 53452 33406 53454 33458
rect 53506 33406 53620 33458
rect 53452 33404 53620 33406
rect 53900 33516 54180 33572
rect 54236 34188 54404 34244
rect 54236 33572 54292 34188
rect 54460 34132 54516 34142
rect 53452 33394 53508 33404
rect 52892 33282 52948 33292
rect 53340 33348 53396 33358
rect 53340 33254 53396 33292
rect 53900 33348 53956 33516
rect 54236 33506 54292 33516
rect 54348 34130 54516 34132
rect 54348 34078 54462 34130
rect 54514 34078 54516 34130
rect 54348 34076 54516 34078
rect 53900 33254 53956 33292
rect 54124 33348 54180 33358
rect 54348 33348 54404 34076
rect 54460 34066 54516 34076
rect 54460 33572 54516 33582
rect 54572 33572 54628 34300
rect 54460 33570 54628 33572
rect 54460 33518 54462 33570
rect 54514 33518 54628 33570
rect 54460 33516 54628 33518
rect 54684 34130 54740 34142
rect 54684 34078 54686 34130
rect 54738 34078 54740 34130
rect 54460 33506 54516 33516
rect 54684 33348 54740 34078
rect 54124 33346 54404 33348
rect 54124 33294 54126 33346
rect 54178 33294 54404 33346
rect 54124 33292 54404 33294
rect 54460 33292 54684 33348
rect 52780 32452 52836 33180
rect 52780 32386 52836 32396
rect 53564 33234 53620 33246
rect 53564 33182 53566 33234
rect 53618 33182 53620 33234
rect 53564 33124 53620 33182
rect 54124 33124 54180 33292
rect 53564 33068 54180 33124
rect 52668 31826 52724 31836
rect 53004 32116 53060 32126
rect 53004 31666 53060 32060
rect 53564 32004 53620 33068
rect 54460 32786 54516 33292
rect 54684 33282 54740 33292
rect 54460 32734 54462 32786
rect 54514 32734 54516 32786
rect 54460 32722 54516 32734
rect 54684 32564 54740 32574
rect 54572 32562 54740 32564
rect 54572 32510 54686 32562
rect 54738 32510 54740 32562
rect 54572 32508 54740 32510
rect 53564 31938 53620 31948
rect 53676 32452 53732 32462
rect 53004 31614 53006 31666
rect 53058 31614 53060 31666
rect 53004 31602 53060 31614
rect 53340 31892 53396 31902
rect 53340 31666 53396 31836
rect 53676 31778 53732 32396
rect 54124 32452 54180 32462
rect 54124 32358 54180 32396
rect 53676 31726 53678 31778
rect 53730 31726 53732 31778
rect 53676 31714 53732 31726
rect 54572 31892 54628 32508
rect 54684 32498 54740 32508
rect 54572 31778 54628 31836
rect 54572 31726 54574 31778
rect 54626 31726 54628 31778
rect 54572 31714 54628 31726
rect 53340 31614 53342 31666
rect 53394 31614 53396 31666
rect 53340 31602 53396 31614
rect 52668 31554 52724 31566
rect 52668 31502 52670 31554
rect 52722 31502 52724 31554
rect 52668 31332 52724 31502
rect 54460 31556 54516 31566
rect 54460 31462 54516 31500
rect 52668 31266 52724 31276
rect 52444 31106 52500 31118
rect 52444 31054 52446 31106
rect 52498 31054 52500 31106
rect 52332 29540 52388 29550
rect 52332 29446 52388 29484
rect 52220 29260 52388 29316
rect 51996 29222 52052 29260
rect 51772 28756 51828 28766
rect 51772 28642 51828 28700
rect 51772 28590 51774 28642
rect 51826 28590 51828 28642
rect 51772 28578 51828 28590
rect 52108 28756 52164 28766
rect 52108 28530 52164 28700
rect 52108 28478 52110 28530
rect 52162 28478 52164 28530
rect 52108 28466 52164 28478
rect 52108 28308 52164 28318
rect 51548 27858 51716 27860
rect 51548 27806 51550 27858
rect 51602 27806 51716 27858
rect 51548 27804 51716 27806
rect 51996 28196 52052 28206
rect 51996 27860 52052 28140
rect 52108 27970 52164 28252
rect 52108 27918 52110 27970
rect 52162 27918 52164 27970
rect 52108 27906 52164 27918
rect 51548 27794 51604 27804
rect 51996 27794 52052 27804
rect 51324 27748 51380 27758
rect 51324 27654 51380 27692
rect 51436 27636 51492 27646
rect 51436 27074 51492 27580
rect 51996 27634 52052 27646
rect 51996 27582 51998 27634
rect 52050 27582 52052 27634
rect 51436 27022 51438 27074
rect 51490 27022 51492 27074
rect 51436 26180 51492 27022
rect 51660 27300 51716 27310
rect 51996 27300 52052 27582
rect 52220 27636 52276 27646
rect 52108 27300 52164 27310
rect 51996 27298 52164 27300
rect 51996 27246 52110 27298
rect 52162 27246 52164 27298
rect 51996 27244 52164 27246
rect 51660 27074 51716 27244
rect 52108 27234 52164 27244
rect 51660 27022 51662 27074
rect 51714 27022 51716 27074
rect 51660 27010 51716 27022
rect 51884 27074 51940 27086
rect 51884 27022 51886 27074
rect 51938 27022 51940 27074
rect 51548 26962 51604 26974
rect 51548 26910 51550 26962
rect 51602 26910 51604 26962
rect 51548 26908 51604 26910
rect 51548 26852 51716 26908
rect 51660 26402 51716 26852
rect 51884 26852 51940 27022
rect 51884 26786 51940 26796
rect 51660 26350 51662 26402
rect 51714 26350 51716 26402
rect 51660 26338 51716 26350
rect 51436 26124 51716 26180
rect 51324 25396 51380 25406
rect 51324 24834 51380 25340
rect 51436 25282 51492 25294
rect 51436 25230 51438 25282
rect 51490 25230 51492 25282
rect 51436 24948 51492 25230
rect 51660 24948 51716 26124
rect 52220 26068 52276 27580
rect 52220 26002 52276 26012
rect 51772 25282 51828 25294
rect 51772 25230 51774 25282
rect 51826 25230 51828 25282
rect 51772 25060 51828 25230
rect 51772 25004 52052 25060
rect 51996 24948 52052 25004
rect 51660 24892 51828 24948
rect 51996 24892 52164 24948
rect 51436 24882 51492 24892
rect 51324 24782 51326 24834
rect 51378 24782 51380 24834
rect 51324 24770 51380 24782
rect 51548 24276 51604 24286
rect 51548 24164 51604 24220
rect 51548 24108 51716 24164
rect 51436 24052 51492 24062
rect 51436 23938 51492 23996
rect 51436 23886 51438 23938
rect 51490 23886 51492 23938
rect 51436 23874 51492 23886
rect 51660 23938 51716 24108
rect 51660 23886 51662 23938
rect 51714 23886 51716 23938
rect 51324 23716 51380 23726
rect 51324 23622 51380 23660
rect 51548 23156 51604 23166
rect 51548 22820 51604 23100
rect 51324 22764 51604 22820
rect 51660 22932 51716 23886
rect 51324 22260 51380 22764
rect 51548 22260 51604 22270
rect 51324 22204 51492 22260
rect 51212 20850 51268 20860
rect 51324 21698 51380 21710
rect 51324 21646 51326 21698
rect 51378 21646 51380 21698
rect 50988 20692 51044 20702
rect 50876 20690 51156 20692
rect 50876 20638 50990 20690
rect 51042 20638 51156 20690
rect 50876 20636 51156 20638
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50540 20244 50596 20254
rect 50876 20244 50932 20636
rect 50988 20626 51044 20636
rect 51100 20580 51156 20636
rect 51324 20580 51380 21646
rect 51436 21364 51492 22204
rect 51548 22166 51604 22204
rect 51436 21298 51492 21308
rect 51548 21924 51604 21934
rect 51100 20524 51380 20580
rect 51436 20580 51492 20590
rect 51548 20580 51604 21868
rect 51492 20524 51604 20580
rect 51436 20514 51492 20524
rect 50540 20242 50932 20244
rect 50540 20190 50542 20242
rect 50594 20190 50932 20242
rect 50540 20188 50932 20190
rect 50540 19346 50596 20188
rect 50876 20132 50932 20188
rect 50876 20066 50932 20076
rect 50988 20468 51044 20478
rect 50540 19294 50542 19346
rect 50594 19294 50596 19346
rect 50540 19282 50596 19294
rect 50876 19124 50932 19134
rect 50988 19124 51044 20412
rect 51660 20356 51716 22876
rect 51772 20468 51828 24892
rect 51884 24834 51940 24846
rect 51884 24782 51886 24834
rect 51938 24782 51940 24834
rect 51884 24612 51940 24782
rect 51884 22036 51940 24556
rect 51996 24724 52052 24734
rect 51996 23828 52052 24668
rect 51996 23380 52052 23772
rect 51996 23314 52052 23324
rect 52108 23156 52164 24892
rect 51884 21970 51940 21980
rect 51996 23100 52164 23156
rect 52220 23154 52276 23166
rect 52220 23102 52222 23154
rect 52274 23102 52276 23154
rect 51996 22708 52052 23100
rect 51996 20580 52052 22652
rect 52108 22372 52164 22382
rect 52220 22372 52276 23102
rect 52164 22316 52276 22372
rect 52108 22306 52164 22316
rect 52108 22148 52164 22158
rect 52108 22054 52164 22092
rect 51996 20578 52164 20580
rect 51996 20526 51998 20578
rect 52050 20526 52164 20578
rect 51996 20524 52164 20526
rect 51996 20514 52052 20524
rect 51772 20412 51940 20468
rect 51212 20300 51716 20356
rect 51212 19234 51268 20300
rect 51772 20244 51828 20254
rect 51660 20188 51772 20244
rect 51660 20132 51716 20188
rect 51772 20178 51828 20188
rect 51212 19182 51214 19234
rect 51266 19182 51268 19234
rect 51212 19170 51268 19182
rect 51324 20130 51716 20132
rect 51324 20078 51662 20130
rect 51714 20078 51716 20130
rect 51324 20076 51716 20078
rect 50876 19122 51044 19124
rect 50876 19070 50878 19122
rect 50930 19070 51044 19122
rect 50876 19068 51044 19070
rect 50876 19058 50932 19068
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50204 18674 50484 18676
rect 50204 18622 50206 18674
rect 50258 18622 50484 18674
rect 50204 18620 50484 18622
rect 50204 18610 50260 18620
rect 49980 18452 50036 18462
rect 49756 18398 49758 18450
rect 49810 18398 49812 18450
rect 49756 18386 49812 18398
rect 49868 18450 50036 18452
rect 49868 18398 49982 18450
rect 50034 18398 50036 18450
rect 49868 18396 50036 18398
rect 49420 17668 49476 17678
rect 49308 17666 49476 17668
rect 49308 17614 49422 17666
rect 49474 17614 49476 17666
rect 49308 17612 49476 17614
rect 48412 17554 48580 17556
rect 48412 17502 48414 17554
rect 48466 17502 48580 17554
rect 48412 17500 48580 17502
rect 49308 17556 49364 17612
rect 49420 17602 49476 17612
rect 48412 17490 48468 17500
rect 49308 17490 49364 17500
rect 49532 17556 49588 17566
rect 49532 17462 49588 17500
rect 48860 17442 48916 17454
rect 48860 17390 48862 17442
rect 48914 17390 48916 17442
rect 48860 17108 48916 17390
rect 48972 17444 49028 17454
rect 49196 17444 49252 17454
rect 49868 17444 49924 18396
rect 49980 18386 50036 18396
rect 50092 18340 50148 18350
rect 50092 18246 50148 18284
rect 50204 17892 50260 17902
rect 48972 17442 49196 17444
rect 48972 17390 48974 17442
rect 49026 17390 49196 17442
rect 48972 17388 49196 17390
rect 48972 17378 49028 17388
rect 49196 17378 49252 17388
rect 49644 17388 49924 17444
rect 49980 17442 50036 17454
rect 49980 17390 49982 17442
rect 50034 17390 50036 17442
rect 49644 17332 49700 17388
rect 49308 17276 49700 17332
rect 49980 17332 50036 17390
rect 48748 16996 48804 17006
rect 47964 16884 48020 16894
rect 47964 16882 48356 16884
rect 47964 16830 47966 16882
rect 48018 16830 48356 16882
rect 47964 16828 48356 16830
rect 47964 16818 48020 16828
rect 47740 16706 47796 16716
rect 47404 15092 47572 15148
rect 47628 16100 47684 16110
rect 47404 13972 47460 15036
rect 47516 14530 47572 14542
rect 47516 14478 47518 14530
rect 47570 14478 47572 14530
rect 47516 14308 47572 14478
rect 47516 14242 47572 14252
rect 47628 14418 47684 16044
rect 48188 16100 48244 16110
rect 48188 16006 48244 16044
rect 47852 15988 47908 15998
rect 47852 15652 47908 15932
rect 47628 14366 47630 14418
rect 47682 14366 47684 14418
rect 47516 13972 47572 13982
rect 47404 13916 47516 13972
rect 47516 13906 47572 13916
rect 47628 13748 47684 14366
rect 47740 15596 47908 15652
rect 47964 15876 48020 15886
rect 47740 14308 47796 15596
rect 47852 15428 47908 15438
rect 47852 15334 47908 15372
rect 47964 14868 48020 15820
rect 47740 14242 47796 14252
rect 47852 14812 47964 14868
rect 47852 13970 47908 14812
rect 47964 14802 48020 14812
rect 48076 15874 48132 15886
rect 48076 15822 48078 15874
rect 48130 15822 48132 15874
rect 47852 13918 47854 13970
rect 47906 13918 47908 13970
rect 47852 13906 47908 13918
rect 48076 13860 48132 15822
rect 48188 15092 48244 15102
rect 48188 14642 48244 15036
rect 48188 14590 48190 14642
rect 48242 14590 48244 14642
rect 48188 14578 48244 14590
rect 48076 13794 48132 13804
rect 48300 13860 48356 16828
rect 48748 16882 48804 16940
rect 48748 16830 48750 16882
rect 48802 16830 48804 16882
rect 48748 16818 48804 16830
rect 48636 16772 48692 16782
rect 48412 15986 48468 15998
rect 48412 15934 48414 15986
rect 48466 15934 48468 15986
rect 48412 14642 48468 15934
rect 48636 15876 48692 16716
rect 48860 15988 48916 17052
rect 48972 17220 49028 17230
rect 48972 16658 49028 17164
rect 49308 17106 49364 17276
rect 49980 17266 50036 17276
rect 49308 17054 49310 17106
rect 49362 17054 49364 17106
rect 49308 17042 49364 17054
rect 50204 17108 50260 17836
rect 50316 17780 50372 17790
rect 50428 17780 50484 18620
rect 50988 18676 51044 18686
rect 50988 18562 51044 18620
rect 50988 18510 50990 18562
rect 51042 18510 51044 18562
rect 50988 18498 51044 18510
rect 51324 18562 51380 20076
rect 51660 20066 51716 20076
rect 51884 19796 51940 20412
rect 52108 20020 52164 20524
rect 52220 20132 52276 20142
rect 52220 20038 52276 20076
rect 52108 19954 52164 19964
rect 51324 18510 51326 18562
rect 51378 18510 51380 18562
rect 51324 18498 51380 18510
rect 51436 19740 51940 19796
rect 52108 19794 52164 19806
rect 52108 19742 52110 19794
rect 52162 19742 52164 19794
rect 50316 17778 50484 17780
rect 50316 17726 50318 17778
rect 50370 17726 50484 17778
rect 50316 17724 50484 17726
rect 50316 17714 50372 17724
rect 49756 16882 49812 16894
rect 49756 16830 49758 16882
rect 49810 16830 49812 16882
rect 49756 16772 49812 16830
rect 50204 16882 50260 17052
rect 50428 16996 50484 17724
rect 50652 18450 50708 18462
rect 50652 18398 50654 18450
rect 50706 18398 50708 18450
rect 50652 17666 50708 18398
rect 50652 17614 50654 17666
rect 50706 17614 50708 17666
rect 50652 17444 50708 17614
rect 50652 17388 51044 17444
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50428 16930 50484 16940
rect 50204 16830 50206 16882
rect 50258 16830 50260 16882
rect 50204 16818 50260 16830
rect 49756 16706 49812 16716
rect 50876 16770 50932 16782
rect 50876 16718 50878 16770
rect 50930 16718 50932 16770
rect 48972 16606 48974 16658
rect 49026 16606 49028 16658
rect 48972 16212 49028 16606
rect 49084 16324 49140 16334
rect 49532 16324 49588 16334
rect 49140 16268 49476 16324
rect 49084 16230 49140 16268
rect 48972 16146 49028 16156
rect 49308 16098 49364 16110
rect 49308 16046 49310 16098
rect 49362 16046 49364 16098
rect 49308 15988 49364 16046
rect 48860 15932 49364 15988
rect 48636 15810 48692 15820
rect 49308 15652 49364 15662
rect 49308 15538 49364 15596
rect 49308 15486 49310 15538
rect 49362 15486 49364 15538
rect 49308 15474 49364 15486
rect 48748 15428 48804 15438
rect 48412 14590 48414 14642
rect 48466 14590 48468 14642
rect 48412 13972 48468 14590
rect 48524 15204 48580 15214
rect 48524 14530 48580 15148
rect 48748 15148 48804 15372
rect 48860 15316 48916 15354
rect 48860 15250 48916 15260
rect 48972 15316 49028 15326
rect 49308 15316 49364 15326
rect 48972 15314 49364 15316
rect 48972 15262 48974 15314
rect 49026 15262 49310 15314
rect 49362 15262 49364 15314
rect 48972 15260 49364 15262
rect 48972 15250 49028 15260
rect 49308 15250 49364 15260
rect 48748 15092 48916 15148
rect 48524 14478 48526 14530
rect 48578 14478 48580 14530
rect 48524 14466 48580 14478
rect 48860 14308 48916 15092
rect 48860 14252 49252 14308
rect 48860 13972 48916 13982
rect 48412 13970 48916 13972
rect 48412 13918 48862 13970
rect 48914 13918 48916 13970
rect 48412 13916 48916 13918
rect 48860 13906 48916 13916
rect 49084 13972 49140 13982
rect 48300 13804 48804 13860
rect 47628 13682 47684 13692
rect 48300 13524 48356 13804
rect 48748 13746 48804 13804
rect 49084 13858 49140 13916
rect 49084 13806 49086 13858
rect 49138 13806 49140 13858
rect 49084 13794 49140 13806
rect 48748 13694 48750 13746
rect 48802 13694 48804 13746
rect 48748 13682 48804 13694
rect 49196 13746 49252 14252
rect 49196 13694 49198 13746
rect 49250 13694 49252 13746
rect 49196 13682 49252 13694
rect 49420 13524 49476 16268
rect 49532 16210 49588 16268
rect 50204 16324 50260 16334
rect 49532 16158 49534 16210
rect 49586 16158 49588 16210
rect 49532 16146 49588 16158
rect 49868 16212 49924 16250
rect 50204 16230 50260 16268
rect 49868 16146 49924 16156
rect 50764 16212 50820 16222
rect 50876 16212 50932 16718
rect 50764 16210 50932 16212
rect 50764 16158 50766 16210
rect 50818 16158 50932 16210
rect 50764 16156 50932 16158
rect 50764 16146 50820 16156
rect 50428 16100 50484 16110
rect 50092 16098 50484 16100
rect 50092 16046 50430 16098
rect 50482 16046 50484 16098
rect 50092 16044 50484 16046
rect 49644 15988 49700 15998
rect 49644 15986 49812 15988
rect 49644 15934 49646 15986
rect 49698 15934 49812 15986
rect 49644 15932 49812 15934
rect 49644 15922 49700 15932
rect 49756 15316 49812 15932
rect 50092 15652 50148 16044
rect 50428 16034 50484 16044
rect 50876 15988 50932 15998
rect 50876 15894 50932 15932
rect 50652 15876 50708 15886
rect 50428 15874 50708 15876
rect 50428 15822 50654 15874
rect 50706 15822 50708 15874
rect 50428 15820 50708 15822
rect 50428 15764 50484 15820
rect 50652 15810 50708 15820
rect 50092 15586 50148 15596
rect 50204 15708 50484 15764
rect 50556 15708 50820 15718
rect 50092 15428 50148 15438
rect 50092 15334 50148 15372
rect 49756 15250 49812 15260
rect 49868 15314 49924 15326
rect 49868 15262 49870 15314
rect 49922 15262 49924 15314
rect 49644 15204 49700 15214
rect 49532 15202 49700 15204
rect 49532 15150 49646 15202
rect 49698 15150 49700 15202
rect 49532 15148 49700 15150
rect 49532 15092 49588 15148
rect 49644 15138 49700 15148
rect 49868 15204 49924 15262
rect 49868 15138 49924 15148
rect 49532 15026 49588 15036
rect 50204 14980 50260 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50988 15652 51044 17388
rect 51436 16996 51492 19740
rect 51660 19572 51716 19582
rect 51660 19346 51716 19516
rect 52108 19460 52164 19742
rect 52332 19684 52388 29260
rect 52444 28196 52500 31054
rect 52780 31108 52836 31118
rect 52444 28130 52500 28140
rect 52668 30212 52724 30222
rect 52668 27972 52724 30156
rect 52780 28866 52836 31052
rect 53564 31108 53620 31118
rect 53564 31014 53620 31052
rect 53900 31108 53956 31118
rect 53900 31106 54068 31108
rect 53900 31054 53902 31106
rect 53954 31054 54068 31106
rect 53900 31052 54068 31054
rect 53900 31042 53956 31052
rect 53004 30882 53060 30894
rect 53004 30830 53006 30882
rect 53058 30830 53060 30882
rect 53004 29428 53060 30830
rect 53228 30882 53284 30894
rect 53228 30830 53230 30882
rect 53282 30830 53284 30882
rect 53228 30212 53284 30830
rect 53228 30146 53284 30156
rect 53340 30100 53396 30110
rect 53340 30006 53396 30044
rect 53228 29428 53284 29438
rect 53004 29426 53396 29428
rect 53004 29374 53230 29426
rect 53282 29374 53396 29426
rect 53004 29372 53396 29374
rect 53228 29362 53284 29372
rect 52780 28814 52782 28866
rect 52834 28814 52836 28866
rect 52780 28802 52836 28814
rect 53116 28644 53172 28654
rect 53116 28642 53284 28644
rect 53116 28590 53118 28642
rect 53170 28590 53284 28642
rect 53116 28588 53284 28590
rect 53116 28578 53172 28588
rect 53004 28196 53060 28206
rect 52724 27916 52836 27972
rect 52668 27878 52724 27916
rect 52444 27858 52500 27870
rect 52444 27806 52446 27858
rect 52498 27806 52500 27858
rect 52444 26908 52500 27806
rect 52556 27746 52612 27758
rect 52556 27694 52558 27746
rect 52610 27694 52612 27746
rect 52556 27076 52612 27694
rect 52780 27076 52836 27916
rect 53004 27858 53060 28140
rect 53004 27806 53006 27858
rect 53058 27806 53060 27858
rect 53004 27794 53060 27806
rect 52892 27748 52948 27758
rect 52892 27300 52948 27692
rect 53116 27300 53172 27310
rect 52892 27298 53172 27300
rect 52892 27246 53118 27298
rect 53170 27246 53172 27298
rect 52892 27244 53172 27246
rect 53116 27234 53172 27244
rect 52892 27076 52948 27086
rect 52780 27074 52948 27076
rect 52780 27022 52894 27074
rect 52946 27022 52948 27074
rect 52780 27020 52948 27022
rect 52556 27010 52612 27020
rect 52892 27010 52948 27020
rect 52668 26962 52724 26974
rect 52668 26910 52670 26962
rect 52722 26910 52724 26962
rect 52668 26908 52724 26910
rect 53228 26908 53284 28588
rect 53340 28530 53396 29372
rect 53676 29314 53732 29326
rect 53676 29262 53678 29314
rect 53730 29262 53732 29314
rect 53676 28868 53732 29262
rect 53676 28802 53732 28812
rect 53340 28478 53342 28530
rect 53394 28478 53396 28530
rect 53340 28466 53396 28478
rect 53900 28530 53956 28542
rect 53900 28478 53902 28530
rect 53954 28478 53956 28530
rect 52444 26852 52724 26908
rect 52444 24610 52500 24622
rect 52444 24558 52446 24610
rect 52498 24558 52500 24610
rect 52444 21700 52500 24558
rect 52556 22036 52612 26852
rect 52668 26628 52724 26852
rect 52780 26852 52836 26862
rect 52780 26758 52836 26796
rect 53116 26852 53284 26908
rect 53340 28308 53396 28318
rect 53340 26908 53396 28252
rect 53676 28196 53732 28206
rect 53900 28196 53956 28478
rect 53732 28140 53844 28196
rect 53676 28130 53732 28140
rect 53564 27972 53620 27982
rect 53788 27972 53844 28140
rect 53900 28130 53956 28140
rect 53788 27916 53956 27972
rect 53564 27858 53620 27916
rect 53564 27806 53566 27858
rect 53618 27806 53620 27858
rect 53564 27794 53620 27806
rect 53900 27186 53956 27916
rect 53900 27134 53902 27186
rect 53954 27134 53956 27186
rect 53900 27122 53956 27134
rect 53452 27076 53508 27086
rect 53788 27076 53844 27086
rect 53452 27074 53844 27076
rect 53452 27022 53454 27074
rect 53506 27022 53790 27074
rect 53842 27022 53844 27074
rect 53452 27020 53844 27022
rect 53452 27010 53508 27020
rect 53788 27010 53844 27020
rect 54012 26908 54068 31052
rect 54236 31106 54292 31118
rect 54236 31054 54238 31106
rect 54290 31054 54292 31106
rect 54124 30212 54180 30222
rect 54124 28082 54180 30156
rect 54236 30100 54292 31054
rect 54572 31108 54628 31118
rect 54572 30994 54628 31052
rect 54572 30942 54574 30994
rect 54626 30942 54628 30994
rect 54460 30212 54516 30222
rect 54460 30118 54516 30156
rect 54236 30034 54292 30044
rect 54572 29652 54628 30942
rect 54460 29596 54628 29652
rect 54348 28644 54404 28654
rect 54348 28530 54404 28588
rect 54348 28478 54350 28530
rect 54402 28478 54404 28530
rect 54348 28466 54404 28478
rect 54124 28030 54126 28082
rect 54178 28030 54180 28082
rect 54124 28018 54180 28030
rect 54460 27860 54516 29596
rect 54572 29428 54628 29438
rect 54572 29334 54628 29372
rect 54796 29204 54852 35308
rect 54908 35196 55076 35308
rect 55244 35364 55300 37100
rect 55356 37090 55412 37100
rect 55580 36652 55972 36708
rect 55468 35586 55524 35598
rect 55468 35534 55470 35586
rect 55522 35534 55524 35586
rect 55468 35476 55524 35534
rect 55244 35298 55300 35308
rect 55356 35420 55524 35476
rect 55020 35140 55076 35196
rect 55020 35084 55188 35140
rect 54908 35028 54964 35038
rect 54908 34130 54964 34972
rect 54908 34078 54910 34130
rect 54962 34078 54964 34130
rect 54908 34066 54964 34078
rect 55020 34130 55076 34142
rect 55020 34078 55022 34130
rect 55074 34078 55076 34130
rect 55020 33684 55076 34078
rect 55132 34132 55188 35084
rect 55356 34916 55412 35420
rect 55580 35364 55636 36652
rect 55804 36482 55860 36494
rect 55804 36430 55806 36482
rect 55858 36430 55860 36482
rect 55804 35812 55860 36430
rect 55916 36372 55972 36652
rect 56028 36596 56084 36634
rect 56028 36530 56084 36540
rect 56028 36372 56084 36382
rect 55916 36370 56084 36372
rect 55916 36318 56030 36370
rect 56082 36318 56084 36370
rect 55916 36316 56084 36318
rect 56028 36306 56084 36316
rect 55804 35756 55972 35812
rect 55916 35588 55972 35756
rect 55804 35532 55972 35588
rect 55468 35308 55636 35364
rect 55692 35476 55748 35486
rect 55468 35252 55524 35308
rect 55468 35138 55524 35196
rect 55468 35086 55470 35138
rect 55522 35086 55524 35138
rect 55468 35074 55524 35086
rect 55580 35140 55636 35150
rect 55580 35046 55636 35084
rect 55692 35028 55748 35420
rect 55804 35252 55860 35532
rect 56028 35474 56084 35486
rect 56028 35422 56030 35474
rect 56082 35422 56084 35474
rect 55804 35186 55860 35196
rect 55916 35364 55972 35374
rect 55916 35028 55972 35308
rect 55692 34962 55748 34972
rect 55804 34972 55972 35028
rect 55356 34860 55524 34916
rect 55468 34468 55524 34860
rect 55804 34914 55860 34972
rect 55804 34862 55806 34914
rect 55858 34862 55860 34914
rect 55468 34412 55748 34468
rect 55244 34356 55300 34366
rect 55244 34354 55636 34356
rect 55244 34302 55246 34354
rect 55298 34302 55636 34354
rect 55244 34300 55636 34302
rect 55244 34290 55300 34300
rect 55132 34076 55300 34132
rect 55020 33618 55076 33628
rect 54908 33572 54964 33582
rect 54908 33348 54964 33516
rect 55020 33348 55076 33358
rect 54908 33346 55076 33348
rect 54908 33294 55022 33346
rect 55074 33294 55076 33346
rect 54908 33292 55076 33294
rect 55020 31556 55076 33292
rect 55020 31490 55076 31500
rect 55020 30884 55076 30894
rect 55020 30790 55076 30828
rect 55132 30212 55188 30222
rect 55020 29988 55076 29998
rect 55020 29894 55076 29932
rect 55132 29426 55188 30156
rect 55132 29374 55134 29426
rect 55186 29374 55188 29426
rect 55132 29362 55188 29374
rect 54908 29316 54964 29326
rect 54908 29222 54964 29260
rect 55244 29204 55300 34076
rect 55580 34130 55636 34300
rect 55580 34078 55582 34130
rect 55634 34078 55636 34130
rect 55580 34066 55636 34078
rect 55580 33908 55636 33918
rect 55356 33906 55636 33908
rect 55356 33854 55582 33906
rect 55634 33854 55636 33906
rect 55356 33852 55636 33854
rect 55356 31666 55412 33852
rect 55580 33842 55636 33852
rect 55692 33572 55748 34412
rect 55580 33516 55692 33572
rect 55468 33460 55524 33470
rect 55468 33366 55524 33404
rect 55580 32564 55636 33516
rect 55692 33506 55748 33516
rect 55804 33236 55860 34862
rect 56028 34916 56084 35422
rect 56028 34850 56084 34860
rect 55916 34802 55972 34814
rect 55916 34750 55918 34802
rect 55970 34750 55972 34802
rect 55916 34242 55972 34750
rect 55916 34190 55918 34242
rect 55970 34190 55972 34242
rect 55916 34178 55972 34190
rect 56140 33684 56196 38612
rect 56364 38500 56420 39454
rect 56252 38444 56420 38500
rect 56700 38724 56756 40460
rect 56812 38834 56868 41356
rect 56924 40628 56980 43484
rect 57036 42868 57092 44268
rect 57036 42802 57092 42812
rect 57036 42420 57092 42430
rect 57036 41970 57092 42364
rect 57036 41918 57038 41970
rect 57090 41918 57092 41970
rect 57036 41906 57092 41918
rect 56924 40562 56980 40572
rect 57036 41076 57092 41086
rect 56812 38782 56814 38834
rect 56866 38782 56868 38834
rect 56812 38770 56868 38782
rect 57036 40516 57092 41020
rect 57036 38668 57092 40460
rect 57148 39732 57204 45388
rect 57260 43540 57316 43550
rect 57260 42754 57316 43484
rect 57372 42980 57428 45500
rect 57708 45220 57764 47068
rect 57820 48130 57876 48142
rect 57820 48078 57822 48130
rect 57874 48078 57876 48130
rect 57820 46900 57876 48078
rect 58044 48132 58100 49308
rect 58156 49252 58212 52108
rect 58156 49186 58212 49196
rect 58268 49810 58324 52220
rect 58380 51492 58436 52782
rect 58940 52834 58996 52846
rect 58940 52782 58942 52834
rect 58994 52782 58996 52834
rect 58828 52164 58884 52202
rect 58828 52098 58884 52108
rect 58380 51426 58436 51436
rect 58828 51938 58884 51950
rect 58828 51886 58830 51938
rect 58882 51886 58884 51938
rect 58828 51380 58884 51886
rect 58828 51314 58884 51324
rect 58716 51044 58772 51054
rect 58716 50594 58772 50988
rect 58716 50542 58718 50594
rect 58770 50542 58772 50594
rect 58716 50530 58772 50542
rect 58492 50484 58548 50522
rect 58492 50418 58548 50428
rect 58268 49758 58270 49810
rect 58322 49758 58324 49810
rect 58156 49028 58212 49038
rect 58156 48934 58212 48972
rect 58268 48804 58324 49758
rect 58716 49810 58772 49822
rect 58716 49758 58718 49810
rect 58770 49758 58772 49810
rect 58492 49698 58548 49710
rect 58492 49646 58494 49698
rect 58546 49646 58548 49698
rect 58380 49140 58436 49150
rect 58380 49046 58436 49084
rect 58492 48916 58548 49646
rect 58716 49252 58772 49758
rect 58716 49186 58772 49196
rect 58940 49810 58996 52782
rect 58940 49758 58942 49810
rect 58994 49758 58996 49810
rect 58492 48850 58548 48860
rect 58044 48066 58100 48076
rect 58156 48748 58324 48804
rect 58716 48804 58772 48814
rect 58940 48804 58996 49758
rect 59052 52164 59108 52174
rect 59052 49812 59108 52108
rect 59612 52164 59668 52174
rect 59612 52070 59668 52108
rect 59388 51604 59444 51614
rect 59164 51268 59220 51278
rect 59164 50482 59220 51212
rect 59388 50594 59444 51548
rect 59948 51266 60004 55132
rect 61068 55094 61124 55132
rect 60732 55076 60788 55086
rect 60732 55074 61012 55076
rect 60732 55022 60734 55074
rect 60786 55022 61012 55074
rect 60732 55020 61012 55022
rect 60732 55010 60788 55020
rect 60508 54404 60564 54414
rect 60508 54402 60676 54404
rect 60508 54350 60510 54402
rect 60562 54350 60676 54402
rect 60508 54348 60676 54350
rect 60508 54338 60564 54348
rect 60284 52836 60340 52846
rect 60172 52834 60340 52836
rect 60172 52782 60286 52834
rect 60338 52782 60340 52834
rect 60172 52780 60340 52782
rect 59948 51214 59950 51266
rect 60002 51214 60004 51266
rect 59948 51202 60004 51214
rect 60060 51938 60116 51950
rect 60060 51886 60062 51938
rect 60114 51886 60116 51938
rect 60060 51268 60116 51886
rect 60060 51202 60116 51212
rect 60172 51044 60228 52780
rect 60284 52770 60340 52780
rect 59388 50542 59390 50594
rect 59442 50542 59444 50594
rect 59388 50530 59444 50542
rect 59724 50988 60228 51044
rect 60396 51268 60452 51278
rect 60396 51154 60452 51212
rect 60396 51102 60398 51154
rect 60450 51102 60452 51154
rect 59164 50430 59166 50482
rect 59218 50430 59220 50482
rect 59164 50418 59220 50430
rect 59052 49746 59108 49756
rect 59388 49698 59444 49710
rect 59388 49646 59390 49698
rect 59442 49646 59444 49698
rect 59276 49140 59332 49150
rect 59276 49046 59332 49084
rect 59052 49028 59108 49038
rect 59052 48934 59108 48972
rect 59164 48804 59220 48814
rect 58940 48748 59108 48804
rect 58044 47348 58100 47358
rect 57820 46834 57876 46844
rect 57932 47234 57988 47246
rect 57932 47182 57934 47234
rect 57986 47182 57988 47234
rect 57932 45892 57988 47182
rect 57932 45826 57988 45836
rect 57708 45154 57764 45164
rect 57372 42914 57428 42924
rect 57596 44212 57652 44222
rect 57260 42702 57262 42754
rect 57314 42702 57316 42754
rect 57260 42690 57316 42702
rect 57372 41860 57428 41870
rect 57372 41766 57428 41804
rect 57596 41636 57652 44156
rect 57820 43652 57876 43662
rect 57820 43558 57876 43596
rect 58044 43540 58100 47292
rect 58156 46674 58212 48748
rect 58716 48710 58772 48748
rect 58940 48356 58996 48366
rect 58268 48242 58324 48254
rect 58268 48190 58270 48242
rect 58322 48190 58324 48242
rect 58268 47460 58324 48190
rect 58492 48242 58548 48254
rect 58492 48190 58494 48242
rect 58546 48190 58548 48242
rect 58380 48130 58436 48142
rect 58380 48078 58382 48130
rect 58434 48078 58436 48130
rect 58380 47572 58436 48078
rect 58492 48132 58548 48190
rect 58940 48242 58996 48300
rect 58940 48190 58942 48242
rect 58994 48190 58996 48242
rect 58940 48178 58996 48190
rect 58492 48066 58548 48076
rect 58380 47506 58436 47516
rect 58492 47796 58548 47806
rect 58268 47394 58324 47404
rect 58492 47458 58548 47740
rect 58492 47406 58494 47458
rect 58546 47406 58548 47458
rect 58492 47394 58548 47406
rect 58940 47458 58996 47470
rect 58940 47406 58942 47458
rect 58994 47406 58996 47458
rect 58156 46622 58158 46674
rect 58210 46622 58212 46674
rect 58156 46610 58212 46622
rect 58380 46340 58436 46350
rect 58268 46284 58380 46340
rect 57932 43484 58100 43540
rect 58156 44772 58212 44782
rect 57820 42196 57876 42206
rect 57932 42196 57988 43484
rect 58156 42754 58212 44716
rect 58156 42702 58158 42754
rect 58210 42702 58212 42754
rect 58156 42690 58212 42702
rect 57876 42140 57988 42196
rect 58044 42308 58100 42318
rect 57820 42102 57876 42140
rect 58044 42082 58100 42252
rect 58044 42030 58046 42082
rect 58098 42030 58100 42082
rect 58044 42018 58100 42030
rect 57372 41580 57652 41636
rect 58156 41972 58212 41982
rect 58268 41972 58324 46284
rect 58380 46274 58436 46284
rect 58716 46228 58772 46238
rect 58716 45778 58772 46172
rect 58940 45892 58996 47406
rect 59052 46674 59108 48748
rect 59052 46622 59054 46674
rect 59106 46622 59108 46674
rect 59052 46610 59108 46622
rect 58940 45836 59108 45892
rect 58716 45726 58718 45778
rect 58770 45726 58772 45778
rect 58716 45714 58772 45726
rect 58940 45668 58996 45678
rect 58828 44884 58884 44894
rect 58828 44790 58884 44828
rect 58716 44098 58772 44110
rect 58716 44046 58718 44098
rect 58770 44046 58772 44098
rect 58716 43652 58772 44046
rect 58716 43586 58772 43596
rect 58940 42754 58996 45612
rect 58940 42702 58942 42754
rect 58994 42702 58996 42754
rect 58940 42690 58996 42702
rect 58156 41970 58324 41972
rect 58156 41918 58158 41970
rect 58210 41918 58324 41970
rect 58156 41916 58324 41918
rect 58604 42530 58660 42542
rect 58604 42478 58606 42530
rect 58658 42478 58660 42530
rect 57260 40292 57316 40302
rect 57260 40178 57316 40236
rect 57260 40126 57262 40178
rect 57314 40126 57316 40178
rect 57260 40114 57316 40126
rect 57260 39732 57316 39742
rect 57148 39676 57260 39732
rect 57260 39666 57316 39676
rect 56252 35140 56308 38444
rect 56588 37940 56644 37950
rect 56588 37378 56644 37884
rect 56700 37604 56756 38668
rect 56812 38612 57092 38668
rect 57148 39508 57204 39518
rect 56812 38276 56868 38612
rect 56812 38210 56868 38220
rect 57148 37938 57204 39452
rect 57148 37886 57150 37938
rect 57202 37886 57204 37938
rect 57148 37874 57204 37886
rect 57260 39396 57316 39406
rect 57260 38722 57316 39340
rect 57260 38670 57262 38722
rect 57314 38670 57316 38722
rect 56700 37548 56868 37604
rect 56588 37326 56590 37378
rect 56642 37326 56644 37378
rect 56588 37314 56644 37326
rect 56700 37380 56756 37390
rect 56700 37286 56756 37324
rect 56700 36484 56756 36494
rect 56700 36390 56756 36428
rect 56476 36370 56532 36382
rect 56476 36318 56478 36370
rect 56530 36318 56532 36370
rect 56476 36148 56532 36318
rect 56476 36082 56532 36092
rect 56700 35924 56756 35934
rect 56812 35924 56868 37548
rect 56924 37268 56980 37278
rect 56924 37174 56980 37212
rect 57260 36484 57316 38670
rect 57372 36932 57428 41580
rect 57820 40964 57876 40974
rect 57820 40962 58100 40964
rect 57820 40910 57822 40962
rect 57874 40910 58100 40962
rect 57820 40908 58100 40910
rect 57820 40898 57876 40908
rect 57596 40514 57652 40526
rect 57596 40462 57598 40514
rect 57650 40462 57652 40514
rect 57596 38668 57652 40462
rect 57820 40404 57876 40414
rect 57820 39060 57876 40348
rect 57820 38994 57876 39004
rect 57932 40180 57988 40190
rect 57932 39730 57988 40124
rect 57932 39678 57934 39730
rect 57986 39678 57988 39730
rect 57708 38836 57764 38846
rect 57932 38836 57988 39678
rect 57708 38834 57988 38836
rect 57708 38782 57710 38834
rect 57762 38782 57988 38834
rect 57708 38780 57988 38782
rect 57708 38770 57764 38780
rect 57596 38612 57764 38668
rect 57708 37940 57764 38612
rect 58044 38612 58100 40908
rect 58156 39396 58212 41916
rect 58156 39330 58212 39340
rect 58268 40628 58324 40638
rect 58268 39844 58324 40572
rect 58604 40404 58660 42478
rect 58828 41972 58884 41982
rect 58884 41916 58996 41972
rect 58828 41878 58884 41916
rect 58940 40628 58996 41916
rect 59052 40852 59108 45836
rect 59164 43314 59220 48748
rect 59276 47684 59332 47694
rect 59276 47590 59332 47628
rect 59276 47124 59332 47134
rect 59388 47124 59444 49646
rect 59612 49028 59668 49038
rect 59612 48934 59668 48972
rect 59724 48468 59780 50988
rect 59948 50820 60004 50830
rect 59948 50706 60004 50764
rect 59948 50654 59950 50706
rect 60002 50654 60004 50706
rect 59948 50642 60004 50654
rect 60396 50428 60452 51102
rect 60620 50932 60676 54348
rect 60956 53956 61012 55020
rect 61068 54404 61124 54414
rect 61516 54404 61572 54414
rect 61852 54404 61908 54414
rect 61068 54402 61908 54404
rect 61068 54350 61070 54402
rect 61122 54350 61518 54402
rect 61570 54350 61854 54402
rect 61906 54350 61908 54402
rect 61068 54348 61908 54350
rect 61068 54338 61124 54348
rect 61516 54338 61572 54348
rect 60956 53900 61348 53956
rect 60732 53508 60788 53518
rect 60732 53414 60788 53452
rect 61068 53508 61124 53518
rect 60732 53172 60788 53182
rect 60732 53078 60788 53116
rect 60732 52276 60788 52286
rect 60732 52182 60788 52220
rect 61068 52274 61124 53452
rect 61068 52222 61070 52274
rect 61122 52222 61124 52274
rect 60844 51492 60900 51502
rect 60844 51398 60900 51436
rect 60620 50866 60676 50876
rect 60060 50372 60452 50428
rect 60508 50818 60564 50830
rect 60508 50766 60510 50818
rect 60562 50766 60564 50818
rect 59836 49810 59892 49822
rect 59836 49758 59838 49810
rect 59890 49758 59892 49810
rect 59836 48804 59892 49758
rect 59948 49364 60004 49374
rect 59948 49138 60004 49308
rect 59948 49086 59950 49138
rect 60002 49086 60004 49138
rect 59948 49074 60004 49086
rect 59836 48738 59892 48748
rect 59724 48402 59780 48412
rect 59332 47068 59444 47124
rect 59612 48354 59668 48366
rect 59612 48302 59614 48354
rect 59666 48302 59668 48354
rect 59276 47058 59332 47068
rect 59612 46004 59668 48302
rect 59612 45938 59668 45948
rect 59724 47458 59780 47470
rect 59724 47406 59726 47458
rect 59778 47406 59780 47458
rect 59724 44548 59780 47406
rect 59836 45666 59892 45678
rect 59836 45614 59838 45666
rect 59890 45614 59892 45666
rect 59836 45108 59892 45614
rect 59836 45042 59892 45052
rect 59836 44548 59892 44558
rect 59724 44546 59892 44548
rect 59724 44494 59838 44546
rect 59890 44494 59892 44546
rect 59724 44492 59892 44494
rect 59612 43538 59668 43550
rect 59612 43486 59614 43538
rect 59666 43486 59668 43538
rect 59164 43262 59166 43314
rect 59218 43262 59220 43314
rect 59164 42196 59220 43262
rect 59164 42130 59220 42140
rect 59276 43316 59332 43326
rect 59052 40786 59108 40796
rect 58940 40572 59220 40628
rect 58604 40402 58884 40404
rect 58604 40350 58606 40402
rect 58658 40350 58884 40402
rect 58604 40348 58884 40350
rect 58604 40338 58660 40348
rect 58268 39618 58324 39788
rect 58268 39566 58270 39618
rect 58322 39566 58324 39618
rect 58044 38546 58100 38556
rect 58268 38388 58324 39566
rect 57820 38332 58324 38388
rect 58492 39060 58548 39070
rect 57820 38050 57876 38332
rect 58492 38274 58548 39004
rect 58492 38222 58494 38274
rect 58546 38222 58548 38274
rect 58492 38210 58548 38222
rect 57820 37998 57822 38050
rect 57874 37998 57876 38050
rect 57820 37986 57876 37998
rect 58828 38052 58884 40348
rect 58940 40402 58996 40414
rect 58940 40350 58942 40402
rect 58994 40350 58996 40402
rect 58940 38164 58996 40350
rect 59052 39618 59108 39630
rect 59052 39566 59054 39618
rect 59106 39566 59108 39618
rect 59052 39060 59108 39566
rect 59052 38994 59108 39004
rect 58940 38098 58996 38108
rect 58828 37958 58884 37996
rect 57708 37042 57764 37884
rect 59164 37492 59220 40572
rect 59276 39618 59332 43260
rect 59500 42530 59556 42542
rect 59500 42478 59502 42530
rect 59554 42478 59556 42530
rect 59500 42420 59556 42478
rect 59500 42354 59556 42364
rect 59612 42084 59668 43486
rect 59724 42754 59780 44492
rect 59836 44482 59892 44492
rect 59724 42702 59726 42754
rect 59778 42702 59780 42754
rect 59724 42690 59780 42702
rect 60060 42756 60116 50372
rect 60284 49700 60340 49710
rect 60284 49606 60340 49644
rect 60508 49138 60564 50766
rect 60620 50708 60676 50718
rect 60620 50614 60676 50652
rect 61068 50428 61124 52222
rect 61180 51604 61236 53900
rect 61292 53842 61348 53900
rect 61292 53790 61294 53842
rect 61346 53790 61348 53842
rect 61292 53778 61348 53790
rect 61292 52836 61348 52846
rect 61292 52834 61460 52836
rect 61292 52782 61294 52834
rect 61346 52782 61460 52834
rect 61292 52780 61460 52782
rect 61292 52770 61348 52780
rect 61292 51604 61348 51614
rect 61180 51602 61348 51604
rect 61180 51550 61294 51602
rect 61346 51550 61348 51602
rect 61180 51548 61348 51550
rect 61292 50818 61348 51548
rect 61404 51156 61460 52780
rect 61516 52276 61572 52286
rect 61516 52182 61572 52220
rect 61404 51090 61460 51100
rect 61292 50766 61294 50818
rect 61346 50766 61348 50818
rect 60956 50372 61124 50428
rect 61180 50482 61236 50494
rect 61180 50430 61182 50482
rect 61234 50430 61236 50482
rect 61180 50372 61236 50430
rect 61292 50428 61348 50766
rect 61516 50932 61572 50942
rect 61516 50706 61572 50876
rect 61516 50654 61518 50706
rect 61570 50654 61572 50706
rect 61516 50642 61572 50654
rect 61292 50372 61460 50428
rect 60508 49086 60510 49138
rect 60562 49086 60564 49138
rect 60508 49074 60564 49086
rect 60844 49698 60900 49710
rect 60844 49646 60846 49698
rect 60898 49646 60900 49698
rect 60732 49026 60788 49038
rect 60732 48974 60734 49026
rect 60786 48974 60788 49026
rect 60508 48916 60564 48926
rect 60284 47124 60340 47134
rect 60284 46674 60340 47068
rect 60284 46622 60286 46674
rect 60338 46622 60340 46674
rect 60284 46610 60340 46622
rect 60508 45890 60564 48860
rect 60732 48804 60788 48974
rect 60732 48738 60788 48748
rect 60844 47572 60900 49646
rect 60956 48244 61012 50372
rect 61180 50306 61236 50316
rect 61292 49810 61348 49822
rect 61292 49758 61294 49810
rect 61346 49758 61348 49810
rect 60956 48178 61012 48188
rect 61068 48802 61124 48814
rect 61068 48750 61070 48802
rect 61122 48750 61124 48802
rect 61068 47908 61124 48750
rect 61292 48132 61348 49758
rect 61404 48580 61460 50372
rect 61628 49026 61684 54348
rect 61852 54338 61908 54348
rect 61852 53506 61908 53518
rect 61852 53454 61854 53506
rect 61906 53454 61908 53506
rect 61852 52836 61908 53454
rect 62188 53508 62244 53518
rect 62188 53414 62244 53452
rect 61964 52836 62020 52846
rect 61852 52834 62132 52836
rect 61852 52782 61966 52834
rect 62018 52782 62132 52834
rect 61852 52780 62132 52782
rect 61964 52770 62020 52780
rect 61964 51940 62020 51950
rect 61852 51938 62020 51940
rect 61852 51886 61966 51938
rect 62018 51886 62020 51938
rect 61852 51884 62020 51886
rect 61740 51266 61796 51278
rect 61740 51214 61742 51266
rect 61794 51214 61796 51266
rect 61740 51156 61796 51214
rect 61740 51090 61796 51100
rect 61740 50932 61796 50942
rect 61852 50932 61908 51884
rect 61964 51874 62020 51884
rect 61796 50876 61908 50932
rect 61964 51154 62020 51166
rect 61964 51102 61966 51154
rect 62018 51102 62020 51154
rect 61740 50866 61796 50876
rect 61964 50706 62020 51102
rect 61964 50654 61966 50706
rect 62018 50654 62020 50706
rect 61964 50642 62020 50654
rect 61852 50260 61908 50270
rect 61852 50034 61908 50204
rect 61852 49982 61854 50034
rect 61906 49982 61908 50034
rect 61852 49970 61908 49982
rect 61628 48974 61630 49026
rect 61682 48974 61684 49026
rect 61628 48804 61684 48974
rect 61628 48738 61684 48748
rect 61740 48916 61796 48926
rect 62076 48916 62132 52780
rect 62636 52276 62692 52286
rect 62188 51268 62244 51278
rect 62188 51266 62580 51268
rect 62188 51214 62190 51266
rect 62242 51214 62580 51266
rect 62188 51212 62580 51214
rect 62188 51202 62244 51212
rect 61796 48860 62132 48916
rect 61740 48802 61796 48860
rect 61740 48750 61742 48802
rect 61794 48750 61796 48802
rect 61740 48738 61796 48750
rect 61404 48524 61796 48580
rect 61292 48076 61460 48132
rect 60956 47852 61124 47908
rect 60956 47796 61012 47852
rect 60956 47730 61012 47740
rect 61292 47684 61348 47694
rect 60956 47572 61012 47582
rect 60844 47570 61012 47572
rect 60844 47518 60958 47570
rect 61010 47518 61012 47570
rect 60844 47516 61012 47518
rect 60620 47460 60676 47498
rect 60620 47394 60676 47404
rect 60732 47458 60788 47470
rect 60732 47406 60734 47458
rect 60786 47406 60788 47458
rect 60732 47348 60788 47406
rect 60732 47282 60788 47292
rect 60620 47236 60676 47246
rect 60620 47142 60676 47180
rect 60732 47012 60788 47022
rect 60620 46004 60676 46014
rect 60620 45910 60676 45948
rect 60508 45838 60510 45890
rect 60562 45838 60564 45890
rect 60508 45826 60564 45838
rect 60732 45666 60788 46956
rect 60844 45892 60900 45902
rect 60844 45778 60900 45836
rect 60844 45726 60846 45778
rect 60898 45726 60900 45778
rect 60844 45714 60900 45726
rect 60732 45614 60734 45666
rect 60786 45614 60788 45666
rect 60732 45444 60788 45614
rect 60396 45388 60788 45444
rect 60396 45220 60452 45388
rect 60060 42690 60116 42700
rect 60172 45164 60452 45220
rect 60172 45106 60228 45164
rect 60172 45054 60174 45106
rect 60226 45054 60228 45106
rect 59612 42018 59668 42028
rect 59724 42308 59780 42318
rect 59500 41860 59556 41870
rect 59500 41766 59556 41804
rect 59724 41076 59780 42252
rect 59724 40982 59780 41020
rect 59612 40852 59668 40862
rect 59500 39732 59556 39742
rect 59500 39638 59556 39676
rect 59276 39566 59278 39618
rect 59330 39566 59332 39618
rect 59276 39554 59332 39566
rect 59612 39618 59668 40796
rect 59612 39566 59614 39618
rect 59666 39566 59668 39618
rect 59612 39554 59668 39566
rect 59836 39620 59892 39630
rect 59836 39526 59892 39564
rect 59724 39060 59780 39070
rect 59612 38948 59668 38958
rect 59612 38834 59668 38892
rect 59612 38782 59614 38834
rect 59666 38782 59668 38834
rect 59612 38770 59668 38782
rect 59724 38834 59780 39004
rect 59724 38782 59726 38834
rect 59778 38782 59780 38834
rect 59724 38770 59780 38782
rect 59052 37436 59220 37492
rect 59276 38612 59332 38622
rect 58492 37266 58548 37278
rect 58492 37214 58494 37266
rect 58546 37214 58548 37266
rect 57708 36990 57710 37042
rect 57762 36990 57764 37042
rect 57708 36978 57764 36990
rect 58380 37154 58436 37166
rect 58380 37102 58382 37154
rect 58434 37102 58436 37154
rect 57372 36876 57540 36932
rect 57372 36708 57428 36718
rect 57372 36614 57428 36652
rect 57260 36418 57316 36428
rect 56700 35922 56868 35924
rect 56700 35870 56702 35922
rect 56754 35870 56868 35922
rect 56700 35868 56868 35870
rect 57260 35924 57316 35934
rect 57316 35868 57428 35924
rect 56700 35858 56756 35868
rect 57260 35858 57316 35868
rect 57372 35810 57428 35868
rect 57372 35758 57374 35810
rect 57426 35758 57428 35810
rect 57372 35746 57428 35758
rect 57260 35698 57316 35710
rect 57260 35646 57262 35698
rect 57314 35646 57316 35698
rect 56252 35074 56308 35084
rect 56700 35588 56756 35598
rect 56588 34804 56644 34814
rect 56588 34710 56644 34748
rect 56252 34692 56308 34702
rect 56252 34598 56308 34636
rect 56140 33618 56196 33628
rect 56252 33348 56308 33358
rect 55804 33170 55860 33180
rect 56028 33292 56252 33348
rect 56028 32786 56084 33292
rect 56252 33282 56308 33292
rect 56476 33348 56532 33358
rect 56476 33346 56644 33348
rect 56476 33294 56478 33346
rect 56530 33294 56644 33346
rect 56476 33292 56644 33294
rect 56476 33282 56532 33292
rect 56028 32734 56030 32786
rect 56082 32734 56084 32786
rect 56028 32722 56084 32734
rect 56476 32564 56532 32574
rect 55580 32508 55860 32564
rect 55468 32452 55524 32462
rect 55580 32452 55636 32508
rect 55468 32450 55636 32452
rect 55468 32398 55470 32450
rect 55522 32398 55636 32450
rect 55468 32396 55636 32398
rect 55804 32452 55860 32508
rect 55804 32396 56084 32452
rect 55468 32386 55524 32396
rect 55692 32338 55748 32350
rect 55692 32286 55694 32338
rect 55746 32286 55748 32338
rect 55692 31892 55748 32286
rect 55748 31836 55860 31892
rect 55692 31826 55748 31836
rect 55356 31614 55358 31666
rect 55410 31614 55412 31666
rect 55356 31602 55412 31614
rect 55804 30994 55860 31836
rect 56028 31106 56084 32396
rect 56028 31054 56030 31106
rect 56082 31054 56084 31106
rect 56028 31042 56084 31054
rect 56252 31556 56308 31566
rect 55804 30942 55806 30994
rect 55858 30942 55860 30994
rect 55804 30930 55860 30942
rect 55468 30772 55524 30782
rect 55468 30770 55748 30772
rect 55468 30718 55470 30770
rect 55522 30718 55748 30770
rect 55468 30716 55748 30718
rect 55468 30706 55524 30716
rect 55468 30324 55524 30334
rect 54460 27524 54516 27804
rect 54460 27458 54516 27468
rect 54572 29148 54852 29204
rect 55132 29148 55300 29204
rect 55356 30268 55468 30324
rect 55356 30210 55412 30268
rect 55468 30258 55524 30268
rect 55356 30158 55358 30210
rect 55410 30158 55412 30210
rect 54572 27076 54628 29148
rect 55020 28756 55076 28766
rect 55020 28642 55076 28700
rect 55020 28590 55022 28642
rect 55074 28590 55076 28642
rect 55020 28578 55076 28590
rect 54684 28530 54740 28542
rect 54684 28478 54686 28530
rect 54738 28478 54740 28530
rect 54684 27636 54740 28478
rect 55020 28418 55076 28430
rect 55020 28366 55022 28418
rect 55074 28366 55076 28418
rect 55020 28084 55076 28366
rect 55020 28018 55076 28028
rect 54796 27972 54852 27982
rect 54796 27858 54852 27916
rect 54796 27806 54798 27858
rect 54850 27806 54852 27858
rect 54796 27794 54852 27806
rect 54684 27570 54740 27580
rect 53340 26852 53620 26908
rect 53116 26628 53172 26852
rect 52668 26572 53172 26628
rect 52780 25508 52836 25518
rect 52780 25414 52836 25452
rect 52892 25396 52948 25406
rect 52892 25302 52948 25340
rect 53004 25282 53060 25294
rect 53004 25230 53006 25282
rect 53058 25230 53060 25282
rect 53004 24724 53060 25230
rect 53004 24630 53060 24668
rect 53228 25282 53284 25294
rect 53228 25230 53230 25282
rect 53282 25230 53284 25282
rect 52892 24500 52948 24510
rect 52668 24164 52724 24174
rect 52668 23044 52724 24108
rect 52668 22978 52724 22988
rect 52780 24052 52836 24062
rect 52780 22930 52836 23996
rect 52892 23940 52948 24444
rect 52892 23938 53060 23940
rect 52892 23886 52894 23938
rect 52946 23886 53060 23938
rect 52892 23884 53060 23886
rect 52892 23874 52948 23884
rect 53004 23268 53060 23884
rect 53228 23828 53284 25230
rect 53340 24722 53396 24734
rect 53340 24670 53342 24722
rect 53394 24670 53396 24722
rect 53340 24612 53396 24670
rect 53340 24546 53396 24556
rect 53564 24500 53620 26852
rect 53788 26852 54068 26908
rect 54460 27074 54628 27076
rect 54460 27022 54574 27074
rect 54626 27022 54628 27074
rect 54460 27020 54628 27022
rect 53788 26178 53844 26852
rect 54348 26850 54404 26862
rect 54348 26798 54350 26850
rect 54402 26798 54404 26850
rect 54348 26404 54404 26798
rect 54348 26338 54404 26348
rect 54460 26290 54516 27020
rect 54572 27010 54628 27020
rect 54684 27076 54740 27086
rect 54684 27074 54964 27076
rect 54684 27022 54686 27074
rect 54738 27022 54964 27074
rect 54684 27020 54964 27022
rect 54684 27010 54740 27020
rect 54796 26852 54852 26862
rect 54460 26238 54462 26290
rect 54514 26238 54516 26290
rect 54460 26226 54516 26238
rect 54572 26850 54852 26852
rect 54572 26798 54798 26850
rect 54850 26798 54852 26850
rect 54572 26796 54852 26798
rect 53788 26126 53790 26178
rect 53842 26126 53844 26178
rect 53788 26114 53844 26126
rect 54236 25844 54292 25854
rect 53788 25732 53844 25742
rect 53676 25284 53732 25294
rect 53676 25190 53732 25228
rect 53788 25172 53844 25676
rect 54236 25618 54292 25788
rect 54572 25730 54628 26796
rect 54796 26786 54852 26796
rect 54684 26404 54740 26414
rect 54740 26348 54852 26404
rect 54684 26338 54740 26348
rect 54572 25678 54574 25730
rect 54626 25678 54628 25730
rect 54572 25666 54628 25678
rect 54796 26290 54852 26348
rect 54796 26238 54798 26290
rect 54850 26238 54852 26290
rect 54236 25566 54238 25618
rect 54290 25566 54292 25618
rect 54236 25554 54292 25566
rect 53788 25106 53844 25116
rect 54012 25506 54068 25518
rect 54012 25454 54014 25506
rect 54066 25454 54068 25506
rect 54012 25060 54068 25454
rect 54012 24994 54068 25004
rect 54684 24724 54740 24734
rect 53788 24612 53844 24622
rect 53564 24444 53732 24500
rect 53564 24162 53620 24174
rect 53564 24110 53566 24162
rect 53618 24110 53620 24162
rect 53452 23828 53508 23838
rect 53228 23826 53508 23828
rect 53228 23774 53454 23826
rect 53506 23774 53508 23826
rect 53228 23772 53508 23774
rect 53452 23492 53508 23772
rect 53452 23426 53508 23436
rect 53564 23268 53620 24110
rect 52892 23156 52948 23166
rect 52892 23062 52948 23100
rect 52780 22878 52782 22930
rect 52834 22878 52836 22930
rect 52780 22866 52836 22878
rect 52668 22370 52724 22382
rect 52668 22318 52670 22370
rect 52722 22318 52724 22370
rect 52668 22260 52724 22318
rect 52668 22194 52724 22204
rect 53004 22036 53060 23212
rect 53116 23266 53620 23268
rect 53116 23214 53566 23266
rect 53618 23214 53620 23266
rect 53116 23212 53620 23214
rect 53116 22258 53172 23212
rect 53564 23202 53620 23212
rect 53452 23044 53508 23054
rect 53452 22370 53508 22988
rect 53452 22318 53454 22370
rect 53506 22318 53508 22370
rect 53452 22306 53508 22318
rect 53116 22206 53118 22258
rect 53170 22206 53172 22258
rect 53116 22194 53172 22206
rect 53228 22146 53284 22158
rect 53228 22094 53230 22146
rect 53282 22094 53284 22146
rect 52556 21980 52724 22036
rect 53004 21980 53172 22036
rect 52444 21634 52500 21644
rect 52556 21362 52612 21374
rect 52556 21310 52558 21362
rect 52610 21310 52612 21362
rect 52556 20804 52612 21310
rect 52668 21028 52724 21980
rect 53004 21588 53060 21598
rect 52668 20962 52724 20972
rect 52892 21586 53060 21588
rect 52892 21534 53006 21586
rect 53058 21534 53060 21586
rect 52892 21532 53060 21534
rect 52668 20804 52724 20814
rect 52556 20802 52724 20804
rect 52556 20750 52670 20802
rect 52722 20750 52724 20802
rect 52556 20748 52724 20750
rect 52668 20738 52724 20748
rect 52892 20244 52948 21532
rect 53004 21522 53060 21532
rect 52892 20178 52948 20188
rect 53004 21252 53060 21262
rect 52780 19796 52836 19806
rect 52780 19794 52948 19796
rect 52780 19742 52782 19794
rect 52834 19742 52948 19794
rect 52780 19740 52948 19742
rect 52780 19730 52836 19740
rect 52332 19628 52724 19684
rect 52668 19460 52724 19628
rect 52780 19460 52836 19470
rect 52668 19458 52836 19460
rect 52668 19406 52782 19458
rect 52834 19406 52836 19458
rect 52668 19404 52836 19406
rect 52108 19394 52164 19404
rect 52780 19394 52836 19404
rect 51660 19294 51662 19346
rect 51714 19294 51716 19346
rect 51660 19282 51716 19294
rect 52220 19236 52276 19246
rect 52220 19234 52388 19236
rect 52220 19182 52222 19234
rect 52274 19182 52388 19234
rect 52220 19180 52388 19182
rect 52220 19170 52276 19180
rect 51548 19012 51604 19022
rect 51548 18918 51604 18956
rect 51772 19012 51828 19022
rect 51772 19010 51940 19012
rect 51772 18958 51774 19010
rect 51826 18958 51940 19010
rect 51772 18956 51940 18958
rect 51772 18946 51828 18956
rect 51772 18564 51828 18574
rect 51772 17890 51828 18508
rect 51884 18340 51940 18956
rect 51884 18274 51940 18284
rect 51996 18450 52052 18462
rect 51996 18398 51998 18450
rect 52050 18398 52052 18450
rect 51772 17838 51774 17890
rect 51826 17838 51828 17890
rect 51772 17826 51828 17838
rect 51884 18004 51940 18014
rect 51660 17780 51716 17790
rect 51660 17666 51716 17724
rect 51660 17614 51662 17666
rect 51714 17614 51716 17666
rect 51660 17602 51716 17614
rect 51884 17666 51940 17948
rect 51884 17614 51886 17666
rect 51938 17614 51940 17666
rect 51884 17602 51940 17614
rect 51436 16940 51604 16996
rect 51436 16772 51492 16782
rect 50556 15642 50820 15652
rect 50876 15596 51044 15652
rect 51212 16324 51268 16334
rect 50428 15540 50484 15550
rect 50204 14914 50260 14924
rect 50316 15538 50484 15540
rect 50316 15486 50430 15538
rect 50482 15486 50484 15538
rect 50316 15484 50484 15486
rect 49756 14868 49812 14878
rect 49812 14812 49924 14868
rect 49756 14802 49812 14812
rect 49532 14420 49588 14430
rect 49532 13746 49588 14364
rect 49756 14418 49812 14430
rect 49756 14366 49758 14418
rect 49810 14366 49812 14418
rect 49756 13970 49812 14366
rect 49756 13918 49758 13970
rect 49810 13918 49812 13970
rect 49756 13906 49812 13918
rect 49532 13694 49534 13746
rect 49586 13694 49588 13746
rect 49532 13682 49588 13694
rect 48300 13458 48356 13468
rect 49084 13468 49476 13524
rect 47292 12910 47294 12962
rect 47346 12910 47348 12962
rect 47292 12898 47348 12910
rect 47740 12962 47796 12974
rect 47740 12910 47742 12962
rect 47794 12910 47796 12962
rect 47628 12852 47684 12862
rect 47404 12850 47684 12852
rect 47404 12798 47630 12850
rect 47682 12798 47684 12850
rect 47404 12796 47684 12798
rect 47404 12404 47460 12796
rect 47628 12786 47684 12796
rect 47068 12014 47070 12066
rect 47122 12014 47124 12066
rect 47068 12002 47124 12014
rect 47180 12348 47460 12404
rect 47180 12290 47236 12348
rect 47180 12238 47182 12290
rect 47234 12238 47236 12290
rect 47180 11282 47236 12238
rect 47740 11620 47796 12910
rect 48300 12852 48356 12862
rect 47180 11230 47182 11282
rect 47234 11230 47236 11282
rect 47180 11218 47236 11230
rect 47292 11564 47796 11620
rect 47964 12796 48300 12852
rect 47964 12178 48020 12796
rect 48300 12758 48356 12796
rect 48524 12850 48580 12862
rect 48524 12798 48526 12850
rect 48578 12798 48580 12850
rect 47964 12126 47966 12178
rect 48018 12126 48020 12178
rect 46508 10782 46510 10834
rect 46562 10782 46564 10834
rect 45164 9828 45220 9838
rect 44828 9826 45220 9828
rect 44828 9774 45166 9826
rect 45218 9774 45220 9826
rect 44828 9772 45220 9774
rect 44604 9202 44660 9212
rect 44828 9602 44884 9614
rect 44828 9550 44830 9602
rect 44882 9550 44884 9602
rect 44156 9042 44324 9044
rect 44156 8990 44158 9042
rect 44210 8990 44324 9042
rect 44156 8988 44324 8990
rect 44156 8978 44212 8988
rect 44044 8754 44100 8764
rect 43932 8642 43988 8652
rect 44156 7812 44212 7822
rect 44156 7586 44212 7756
rect 44268 7700 44324 8988
rect 44492 9042 44548 9054
rect 44492 8990 44494 9042
rect 44546 8990 44548 9042
rect 44492 7812 44548 8990
rect 44492 7746 44548 7756
rect 44380 7700 44436 7710
rect 44268 7698 44436 7700
rect 44268 7646 44382 7698
rect 44434 7646 44436 7698
rect 44268 7644 44436 7646
rect 44380 7634 44436 7644
rect 44604 7700 44660 7710
rect 44828 7700 44884 9550
rect 45164 9044 45220 9772
rect 45388 9828 45444 9838
rect 46396 9828 46452 9838
rect 46508 9828 46564 10782
rect 46844 10780 47012 10836
rect 47292 10836 47348 11564
rect 47628 11396 47684 11406
rect 47964 11396 48020 12126
rect 48188 12178 48244 12190
rect 48188 12126 48190 12178
rect 48242 12126 48244 12178
rect 47628 11302 47684 11340
rect 47740 11394 48020 11396
rect 47740 11342 47966 11394
rect 48018 11342 48020 11394
rect 47740 11340 48020 11342
rect 47404 11284 47460 11294
rect 47404 11190 47460 11228
rect 47516 11172 47572 11182
rect 47516 11078 47572 11116
rect 47628 11060 47684 11070
rect 47404 10836 47460 10846
rect 47292 10780 47404 10836
rect 46732 10722 46788 10734
rect 46732 10670 46734 10722
rect 46786 10670 46788 10722
rect 45444 9772 45556 9828
rect 45388 9734 45444 9772
rect 45164 8978 45220 8988
rect 45276 9268 45332 9278
rect 44940 8932 44996 8942
rect 44940 8838 44996 8876
rect 45052 8820 45108 8830
rect 44604 7698 44884 7700
rect 44604 7646 44606 7698
rect 44658 7646 44884 7698
rect 44604 7644 44884 7646
rect 44940 8708 44996 8718
rect 44604 7634 44660 7644
rect 44156 7534 44158 7586
rect 44210 7534 44212 7586
rect 44156 7476 44212 7534
rect 44492 7588 44548 7598
rect 44492 7494 44548 7532
rect 44940 7476 44996 8652
rect 45052 8484 45108 8764
rect 45052 8258 45108 8428
rect 45052 8206 45054 8258
rect 45106 8206 45108 8258
rect 45052 8194 45108 8206
rect 45164 7700 45220 7710
rect 45276 7700 45332 9212
rect 45500 9156 45556 9772
rect 46396 9826 46564 9828
rect 46396 9774 46398 9826
rect 46450 9774 46564 9826
rect 46396 9772 46564 9774
rect 46620 10498 46676 10510
rect 46620 10446 46622 10498
rect 46674 10446 46676 10498
rect 45500 9062 45556 9100
rect 45724 9714 45780 9726
rect 45724 9662 45726 9714
rect 45778 9662 45780 9714
rect 45612 9044 45668 9054
rect 45612 8950 45668 8988
rect 45612 8372 45668 8382
rect 45164 7698 45332 7700
rect 45164 7646 45166 7698
rect 45218 7646 45332 7698
rect 45164 7644 45332 7646
rect 45388 8146 45444 8158
rect 45388 8094 45390 8146
rect 45442 8094 45444 8146
rect 45164 7634 45220 7644
rect 44940 7420 45220 7476
rect 44156 6804 44212 7420
rect 44156 6738 44212 6748
rect 45052 6802 45108 6814
rect 45052 6750 45054 6802
rect 45106 6750 45108 6802
rect 44268 6690 44324 6702
rect 44268 6638 44270 6690
rect 44322 6638 44324 6690
rect 44156 6578 44212 6590
rect 44156 6526 44158 6578
rect 44210 6526 44212 6578
rect 44156 6132 44212 6526
rect 44268 6580 44324 6638
rect 44268 6514 44324 6524
rect 44828 6578 44884 6590
rect 44828 6526 44830 6578
rect 44882 6526 44884 6578
rect 44156 6066 44212 6076
rect 44828 5908 44884 6526
rect 45052 6356 45108 6750
rect 44828 5842 44884 5852
rect 44940 6130 44996 6142
rect 44940 6078 44942 6130
rect 44994 6078 44996 6130
rect 43820 5070 43822 5122
rect 43874 5070 43876 5122
rect 43820 4788 43876 5070
rect 44156 5684 44212 5694
rect 44156 5010 44212 5628
rect 44940 5684 44996 6078
rect 45052 6020 45108 6300
rect 45052 5954 45108 5964
rect 44940 5618 44996 5628
rect 45052 5122 45108 5134
rect 45052 5070 45054 5122
rect 45106 5070 45108 5122
rect 44156 4958 44158 5010
rect 44210 4958 44212 5010
rect 44156 4946 44212 4958
rect 44940 5012 44996 5022
rect 44940 4918 44996 4956
rect 45052 4788 45108 5070
rect 43820 4732 45108 4788
rect 43820 4338 43876 4732
rect 43820 4286 43822 4338
rect 43874 4286 43876 4338
rect 43820 4274 43876 4286
rect 44604 4564 44660 4574
rect 43820 3668 43876 3678
rect 43708 3666 43876 3668
rect 43708 3614 43822 3666
rect 43874 3614 43876 3666
rect 43708 3612 43876 3614
rect 42700 3574 42756 3612
rect 43820 3602 43876 3612
rect 44268 3668 44324 3678
rect 39900 3502 39902 3554
rect 39954 3502 39956 3554
rect 39900 3490 39956 3502
rect 44268 3554 44324 3612
rect 44268 3502 44270 3554
rect 44322 3502 44324 3554
rect 44268 3490 44324 3502
rect 38332 3390 38334 3442
rect 38386 3390 38388 3442
rect 38332 3378 38388 3390
rect 44604 3442 44660 4508
rect 45164 3666 45220 7420
rect 45388 7028 45444 8094
rect 45612 7476 45668 8316
rect 45724 7924 45780 9662
rect 45836 9604 45892 9614
rect 45836 9510 45892 9548
rect 46060 9604 46116 9614
rect 46060 9602 46228 9604
rect 46060 9550 46062 9602
rect 46114 9550 46228 9602
rect 46060 9548 46228 9550
rect 46060 9538 46116 9548
rect 46060 9268 46116 9278
rect 46060 9174 46116 9212
rect 45724 7858 45780 7868
rect 46060 8596 46116 8606
rect 45612 7382 45668 7420
rect 45836 7586 45892 7598
rect 45836 7534 45838 7586
rect 45890 7534 45892 7586
rect 45388 6914 45444 6972
rect 45388 6862 45390 6914
rect 45442 6862 45444 6914
rect 45388 6850 45444 6862
rect 45500 6916 45556 6926
rect 45276 6692 45332 6702
rect 45276 6130 45332 6636
rect 45276 6078 45278 6130
rect 45330 6078 45332 6130
rect 45276 6066 45332 6078
rect 45164 3614 45166 3666
rect 45218 3614 45220 3666
rect 45164 3602 45220 3614
rect 45500 3666 45556 6860
rect 45836 6802 45892 7534
rect 45836 6750 45838 6802
rect 45890 6750 45892 6802
rect 45836 6738 45892 6750
rect 45948 6804 46004 6814
rect 45724 6692 45780 6702
rect 45724 6598 45780 6636
rect 45948 6690 46004 6748
rect 45948 6638 45950 6690
rect 46002 6638 46004 6690
rect 45948 6626 46004 6638
rect 46060 6356 46116 8540
rect 46172 7252 46228 9548
rect 46172 7186 46228 7196
rect 46284 9042 46340 9054
rect 46284 8990 46286 9042
rect 46338 8990 46340 9042
rect 46172 7028 46228 7038
rect 46172 6578 46228 6972
rect 46284 6916 46340 8990
rect 46396 7474 46452 9772
rect 46620 9604 46676 10446
rect 46620 9538 46676 9548
rect 46732 9492 46788 10670
rect 46732 9426 46788 9436
rect 46844 9268 46900 10780
rect 46956 10610 47012 10622
rect 46956 10558 46958 10610
rect 47010 10558 47012 10610
rect 46956 9716 47012 10558
rect 47292 10612 47348 10622
rect 47292 10518 47348 10556
rect 47404 10052 47460 10780
rect 47404 9958 47460 9996
rect 47516 9828 47572 9838
rect 46956 9650 47012 9660
rect 47404 9826 47572 9828
rect 47404 9774 47518 9826
rect 47570 9774 47572 9826
rect 47404 9772 47572 9774
rect 46508 9212 46900 9268
rect 46508 8484 46564 9212
rect 47180 9156 47236 9166
rect 46732 9044 46788 9054
rect 46956 9044 47012 9054
rect 46732 8950 46788 8988
rect 46844 8988 46956 9044
rect 46508 8428 46676 8484
rect 46396 7422 46398 7474
rect 46450 7422 46452 7474
rect 46396 7410 46452 7422
rect 46508 8258 46564 8270
rect 46508 8206 46510 8258
rect 46562 8206 46564 8258
rect 46284 6850 46340 6860
rect 46508 6692 46564 8206
rect 46172 6526 46174 6578
rect 46226 6526 46228 6578
rect 46172 6514 46228 6526
rect 46284 6636 46508 6692
rect 45948 6300 46116 6356
rect 45612 6020 45668 6030
rect 45612 5906 45668 5964
rect 45612 5854 45614 5906
rect 45666 5854 45668 5906
rect 45612 5842 45668 5854
rect 45836 5908 45892 5918
rect 45836 5814 45892 5852
rect 45724 5684 45780 5694
rect 45724 5346 45780 5628
rect 45724 5294 45726 5346
rect 45778 5294 45780 5346
rect 45724 5282 45780 5294
rect 45724 4564 45780 4574
rect 45724 4450 45780 4508
rect 45724 4398 45726 4450
rect 45778 4398 45780 4450
rect 45724 4386 45780 4398
rect 45500 3614 45502 3666
rect 45554 3614 45556 3666
rect 45500 3602 45556 3614
rect 45948 3778 46004 6300
rect 46284 6132 46340 6636
rect 46508 6626 46564 6636
rect 46620 7140 46676 8428
rect 46732 7700 46788 7710
rect 46844 7700 46900 8988
rect 46956 8978 47012 8988
rect 46956 8260 47012 8270
rect 46956 8258 47124 8260
rect 46956 8206 46958 8258
rect 47010 8206 47124 8258
rect 46956 8204 47124 8206
rect 46956 8194 47012 8204
rect 46732 7698 46900 7700
rect 46732 7646 46734 7698
rect 46786 7646 46900 7698
rect 46732 7644 46900 7646
rect 46732 7634 46788 7644
rect 46060 6076 46340 6132
rect 46396 6132 46452 6142
rect 46060 5346 46116 6076
rect 46172 5908 46228 5918
rect 46172 5814 46228 5852
rect 46396 5794 46452 6076
rect 46396 5742 46398 5794
rect 46450 5742 46452 5794
rect 46396 5730 46452 5742
rect 46620 5460 46676 7084
rect 47068 6692 47124 8204
rect 47180 7698 47236 9100
rect 47180 7646 47182 7698
rect 47234 7646 47236 7698
rect 47180 7634 47236 7646
rect 47404 7476 47460 9772
rect 47516 9762 47572 9772
rect 47404 7382 47460 7420
rect 46956 6636 47124 6692
rect 47516 7252 47572 7262
rect 47516 6690 47572 7196
rect 47516 6638 47518 6690
rect 47570 6638 47572 6690
rect 46956 6244 47012 6636
rect 47516 6626 47572 6638
rect 47068 6468 47124 6478
rect 47068 6466 47236 6468
rect 47068 6414 47070 6466
rect 47122 6414 47236 6466
rect 47068 6412 47236 6414
rect 47068 6402 47124 6412
rect 46956 6188 47124 6244
rect 47068 6132 47124 6188
rect 47068 6066 47124 6076
rect 47180 6130 47236 6412
rect 47292 6466 47348 6478
rect 47292 6414 47294 6466
rect 47346 6414 47348 6466
rect 47292 6244 47348 6414
rect 47292 6178 47348 6188
rect 47404 6466 47460 6478
rect 47404 6414 47406 6466
rect 47458 6414 47460 6466
rect 47180 6078 47182 6130
rect 47234 6078 47236 6130
rect 47180 6066 47236 6078
rect 46956 6018 47012 6030
rect 46956 5966 46958 6018
rect 47010 5966 47012 6018
rect 46844 5908 46900 5918
rect 46060 5294 46062 5346
rect 46114 5294 46116 5346
rect 46060 5282 46116 5294
rect 46396 5404 46676 5460
rect 46732 5906 46900 5908
rect 46732 5854 46846 5906
rect 46898 5854 46900 5906
rect 46732 5852 46900 5854
rect 45948 3726 45950 3778
rect 46002 3726 46004 3778
rect 45948 3668 46004 3726
rect 46060 3668 46116 3678
rect 45948 3666 46116 3668
rect 45948 3614 46062 3666
rect 46114 3614 46116 3666
rect 45948 3612 46116 3614
rect 46060 3602 46116 3612
rect 44604 3390 44606 3442
rect 44658 3390 44660 3442
rect 44604 3378 44660 3390
rect 46396 3220 46452 5404
rect 46732 4900 46788 5852
rect 46844 5842 46900 5852
rect 46844 5124 46900 5134
rect 46844 5030 46900 5068
rect 46732 4844 46900 4900
rect 46732 4340 46788 4350
rect 46732 4246 46788 4284
rect 46508 3668 46564 3678
rect 46508 3574 46564 3612
rect 46844 3556 46900 4844
rect 46956 4564 47012 5966
rect 46956 4498 47012 4508
rect 47292 5348 47348 5358
rect 47292 4450 47348 5292
rect 47404 5236 47460 6414
rect 47628 6130 47684 11004
rect 47740 10610 47796 11340
rect 47964 11330 48020 11340
rect 48076 11508 48132 11518
rect 47852 10948 47908 10958
rect 47852 10722 47908 10892
rect 48076 10834 48132 11452
rect 48188 11396 48244 12126
rect 48188 11330 48244 11340
rect 48300 11172 48356 11182
rect 48300 11078 48356 11116
rect 48524 10948 48580 12798
rect 48748 12178 48804 12190
rect 48972 12180 49028 12190
rect 48748 12126 48750 12178
rect 48802 12126 48804 12178
rect 48748 11508 48804 12126
rect 48748 11442 48804 11452
rect 48860 12178 49028 12180
rect 48860 12126 48974 12178
rect 49026 12126 49028 12178
rect 48860 12124 49028 12126
rect 48860 11172 48916 12124
rect 48972 12114 49028 12124
rect 49084 11506 49140 13468
rect 49196 12852 49252 12862
rect 49196 12758 49252 12796
rect 49532 12738 49588 12750
rect 49532 12686 49534 12738
rect 49586 12686 49588 12738
rect 49420 12516 49476 12526
rect 49196 12460 49420 12516
rect 49196 12402 49252 12460
rect 49420 12450 49476 12460
rect 49196 12350 49198 12402
rect 49250 12350 49252 12402
rect 49196 12338 49252 12350
rect 49084 11454 49086 11506
rect 49138 11454 49140 11506
rect 49084 11442 49140 11454
rect 49308 12178 49364 12190
rect 49308 12126 49310 12178
rect 49362 12126 49364 12178
rect 48972 11396 49028 11406
rect 48972 11302 49028 11340
rect 49308 11396 49364 12126
rect 49420 11508 49476 11518
rect 49420 11414 49476 11452
rect 49308 11330 49364 11340
rect 49084 11282 49140 11294
rect 49084 11230 49086 11282
rect 49138 11230 49140 11282
rect 49084 11172 49140 11230
rect 48916 11116 49140 11172
rect 48860 11078 48916 11116
rect 48524 10882 48580 10892
rect 48860 10948 48916 10958
rect 48076 10782 48078 10834
rect 48130 10782 48132 10834
rect 48076 10770 48132 10782
rect 48188 10836 48244 10846
rect 47852 10670 47854 10722
rect 47906 10670 47908 10722
rect 47852 10658 47908 10670
rect 47964 10724 48020 10734
rect 47740 10558 47742 10610
rect 47794 10558 47796 10610
rect 47740 10546 47796 10558
rect 47964 9268 48020 10668
rect 48188 10722 48244 10780
rect 48188 10670 48190 10722
rect 48242 10670 48244 10722
rect 48188 10658 48244 10670
rect 48860 10386 48916 10892
rect 48972 10612 49028 10622
rect 48972 10518 49028 10556
rect 48860 10334 48862 10386
rect 48914 10334 48916 10386
rect 48860 10322 48916 10334
rect 48412 9828 48468 9838
rect 48188 9826 48580 9828
rect 48188 9774 48414 9826
rect 48466 9774 48580 9826
rect 48188 9772 48580 9774
rect 47964 9212 48132 9268
rect 47964 9044 48020 9054
rect 47852 8932 47908 8942
rect 47852 8838 47908 8876
rect 47964 8818 48020 8988
rect 47964 8766 47966 8818
rect 48018 8766 48020 8818
rect 47964 8754 48020 8766
rect 47740 8484 47796 8494
rect 47740 8390 47796 8428
rect 48076 8372 48132 9212
rect 47964 8316 48132 8372
rect 48188 9154 48244 9772
rect 48412 9762 48468 9772
rect 48188 9102 48190 9154
rect 48242 9102 48244 9154
rect 47964 7588 48020 8316
rect 48076 7700 48132 7710
rect 48188 7700 48244 9102
rect 48076 7698 48244 7700
rect 48076 7646 48078 7698
rect 48130 7646 48244 7698
rect 48076 7644 48244 7646
rect 48524 8258 48580 9772
rect 48860 9716 48916 9726
rect 48748 9044 48804 9054
rect 48748 8950 48804 8988
rect 48748 8484 48804 8494
rect 48860 8484 48916 9660
rect 48804 8428 48916 8484
rect 48748 8418 48804 8428
rect 48524 8206 48526 8258
rect 48578 8206 48580 8258
rect 48076 7634 48132 7644
rect 47628 6078 47630 6130
rect 47682 6078 47684 6130
rect 47628 6066 47684 6078
rect 47740 7364 47796 7374
rect 47740 6692 47796 7308
rect 47516 5236 47572 5246
rect 47404 5234 47572 5236
rect 47404 5182 47518 5234
rect 47570 5182 47572 5234
rect 47404 5180 47572 5182
rect 47516 5170 47572 5180
rect 47628 4564 47684 4574
rect 47740 4564 47796 6636
rect 47852 6804 47908 6814
rect 47852 6578 47908 6748
rect 47852 6526 47854 6578
rect 47906 6526 47908 6578
rect 47852 6514 47908 6526
rect 47964 6018 48020 7532
rect 48188 7364 48244 7374
rect 48188 7270 48244 7308
rect 48412 6916 48468 6926
rect 48412 6690 48468 6860
rect 48412 6638 48414 6690
rect 48466 6638 48468 6690
rect 48412 6626 48468 6638
rect 48524 6580 48580 8206
rect 48860 8260 48916 8270
rect 48860 8166 48916 8204
rect 49084 8202 49140 11116
rect 49308 10722 49364 10734
rect 49308 10670 49310 10722
rect 49362 10670 49364 10722
rect 49308 10388 49364 10670
rect 49532 10612 49588 12686
rect 49756 12292 49812 12302
rect 49868 12292 49924 14812
rect 50204 13860 50260 13870
rect 50316 13860 50372 15484
rect 50428 15474 50484 15484
rect 50204 13858 50372 13860
rect 50204 13806 50206 13858
rect 50258 13806 50372 13858
rect 50204 13804 50372 13806
rect 50428 15316 50484 15326
rect 50204 13794 50260 13804
rect 49980 13748 50036 13758
rect 50092 13748 50148 13758
rect 49980 13746 50092 13748
rect 49980 13694 49982 13746
rect 50034 13694 50092 13746
rect 49980 13692 50092 13694
rect 49980 13682 50036 13692
rect 49980 13076 50036 13086
rect 49980 12982 50036 13020
rect 50092 12404 50148 13692
rect 50428 13748 50484 15260
rect 50652 15090 50708 15102
rect 50652 15038 50654 15090
rect 50706 15038 50708 15090
rect 50652 14756 50708 15038
rect 50652 14690 50708 14700
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50652 13972 50708 13982
rect 50652 13878 50708 13916
rect 50428 13682 50484 13692
rect 50092 12338 50148 12348
rect 50204 13524 50260 13534
rect 49756 12290 49924 12292
rect 49756 12238 49758 12290
rect 49810 12238 49924 12290
rect 49756 12236 49924 12238
rect 49756 12226 49812 12236
rect 49868 11394 49924 11406
rect 49868 11342 49870 11394
rect 49922 11342 49924 11394
rect 49868 11172 49924 11342
rect 49868 11106 49924 11116
rect 49532 10546 49588 10556
rect 49308 8820 49364 10332
rect 49420 10500 49476 10510
rect 49420 9044 49476 10444
rect 50092 9602 50148 9614
rect 50092 9550 50094 9602
rect 50146 9550 50148 9602
rect 49420 9042 49588 9044
rect 49420 8990 49422 9042
rect 49474 8990 49588 9042
rect 49420 8988 49588 8990
rect 49420 8978 49476 8988
rect 49308 8764 49476 8820
rect 49084 8150 49086 8202
rect 49138 8150 49140 8202
rect 49420 8260 49476 8764
rect 49420 8194 49476 8204
rect 49084 8138 49140 8150
rect 49308 8148 49364 8158
rect 49196 8036 49252 8074
rect 49196 7970 49252 7980
rect 49308 8034 49364 8092
rect 49308 7982 49310 8034
rect 49362 7982 49364 8034
rect 49196 7812 49252 7822
rect 48860 7364 48916 7374
rect 48916 7308 49140 7364
rect 48860 7270 48916 7308
rect 49084 6690 49140 7308
rect 49084 6638 49086 6690
rect 49138 6638 49140 6690
rect 49084 6626 49140 6638
rect 48636 6580 48692 6590
rect 48524 6578 48692 6580
rect 48524 6526 48638 6578
rect 48690 6526 48692 6578
rect 48524 6524 48692 6526
rect 48636 6514 48692 6524
rect 48748 6578 48804 6590
rect 48748 6526 48750 6578
rect 48802 6526 48804 6578
rect 48188 6466 48244 6478
rect 48188 6414 48190 6466
rect 48242 6414 48244 6466
rect 48188 6132 48244 6414
rect 48188 6066 48244 6076
rect 47964 5966 47966 6018
rect 48018 5966 48020 6018
rect 47964 5954 48020 5966
rect 48076 6020 48132 6030
rect 48076 5926 48132 5964
rect 48748 6020 48804 6526
rect 49084 6468 49140 6478
rect 48860 6412 49084 6468
rect 48860 6130 48916 6412
rect 49084 6402 49140 6412
rect 48860 6078 48862 6130
rect 48914 6078 48916 6130
rect 48860 6066 48916 6078
rect 49084 6132 49140 6142
rect 49196 6132 49252 7756
rect 49084 6130 49252 6132
rect 49084 6078 49086 6130
rect 49138 6078 49252 6130
rect 49084 6076 49252 6078
rect 49308 7028 49364 7982
rect 49084 6066 49140 6076
rect 48748 5926 48804 5964
rect 48524 5012 48580 5022
rect 47628 4562 47796 4564
rect 47628 4510 47630 4562
rect 47682 4510 47796 4562
rect 47628 4508 47796 4510
rect 47964 4676 48020 4686
rect 47628 4498 47684 4508
rect 47292 4398 47294 4450
rect 47346 4398 47348 4450
rect 47292 4386 47348 4398
rect 46956 3778 47012 3790
rect 46956 3726 46958 3778
rect 47010 3726 47012 3778
rect 46956 3666 47012 3726
rect 46956 3614 46958 3666
rect 47010 3614 47012 3666
rect 46956 3602 47012 3614
rect 47964 3666 48020 4620
rect 48076 4452 48132 4462
rect 48076 4358 48132 4396
rect 47964 3614 47966 3666
rect 48018 3614 48020 3666
rect 47964 3602 48020 3614
rect 48524 3668 48580 4956
rect 48972 4564 49028 4574
rect 49308 4564 49364 6972
rect 49532 6802 49588 8988
rect 49644 8932 49700 8942
rect 50092 8932 50148 9550
rect 49700 8876 50148 8932
rect 49644 8838 49700 8876
rect 49532 6750 49534 6802
rect 49586 6750 49588 6802
rect 49532 6468 49588 6750
rect 49980 7588 50036 7598
rect 49980 6578 50036 7532
rect 50204 7364 50260 13468
rect 50876 13076 50932 15596
rect 51212 15540 51268 16268
rect 51436 16210 51492 16716
rect 51436 16158 51438 16210
rect 51490 16158 51492 16210
rect 51436 16146 51492 16158
rect 51548 16548 51604 16940
rect 51548 15988 51604 16492
rect 51996 16884 52052 18398
rect 52332 18450 52388 19180
rect 52556 19234 52612 19246
rect 52556 19182 52558 19234
rect 52610 19182 52612 19234
rect 52556 18564 52612 19182
rect 52556 18498 52612 18508
rect 52332 18398 52334 18450
rect 52386 18398 52388 18450
rect 52220 18228 52276 18238
rect 52220 18134 52276 18172
rect 52108 17892 52164 17902
rect 52108 17554 52164 17836
rect 52332 17780 52388 18398
rect 52892 18452 52948 19740
rect 52892 18386 52948 18396
rect 52556 17780 52612 17790
rect 52332 17778 52612 17780
rect 52332 17726 52558 17778
rect 52610 17726 52612 17778
rect 52332 17724 52612 17726
rect 52556 17714 52612 17724
rect 52108 17502 52110 17554
rect 52162 17502 52164 17554
rect 52108 17490 52164 17502
rect 53004 17332 53060 21196
rect 53116 20914 53172 21980
rect 53228 21924 53284 22094
rect 53228 21858 53284 21868
rect 53340 22146 53396 22158
rect 53340 22094 53342 22146
rect 53394 22094 53396 22146
rect 53340 21812 53396 22094
rect 53340 21746 53396 21756
rect 53452 21474 53508 21486
rect 53452 21422 53454 21474
rect 53506 21422 53508 21474
rect 53452 21364 53508 21422
rect 53676 21364 53732 24444
rect 53788 23716 53844 24556
rect 54684 23940 54740 24668
rect 54796 24276 54852 26238
rect 54908 25732 54964 27020
rect 55132 26908 55188 29148
rect 55356 28866 55412 30158
rect 55580 30100 55636 30110
rect 55468 29428 55524 29438
rect 55468 29334 55524 29372
rect 55356 28814 55358 28866
rect 55410 28814 55412 28866
rect 55356 28802 55412 28814
rect 55468 29092 55524 29102
rect 55244 28420 55300 28430
rect 55244 27746 55300 28364
rect 55244 27694 55246 27746
rect 55298 27694 55300 27746
rect 55244 27074 55300 27694
rect 55356 27748 55412 27758
rect 55356 27654 55412 27692
rect 55468 27636 55524 29036
rect 55580 28642 55636 30044
rect 55692 28868 55748 30716
rect 56028 30212 56084 30250
rect 56028 30146 56084 30156
rect 55804 29988 55860 29998
rect 55804 29894 55860 29932
rect 56028 29988 56084 29998
rect 55916 29540 55972 29550
rect 55916 29446 55972 29484
rect 55804 29426 55860 29438
rect 55804 29374 55806 29426
rect 55858 29374 55860 29426
rect 55804 29204 55860 29374
rect 55804 29138 55860 29148
rect 55916 29204 55972 29214
rect 56028 29204 56084 29932
rect 55916 29202 56084 29204
rect 55916 29150 55918 29202
rect 55970 29150 56084 29202
rect 55916 29148 56084 29150
rect 55916 29138 55972 29148
rect 56252 28980 56308 31500
rect 56476 30884 56532 32508
rect 56588 31556 56644 33292
rect 56588 31490 56644 31500
rect 56588 31332 56644 31342
rect 56588 31106 56644 31276
rect 56588 31054 56590 31106
rect 56642 31054 56644 31106
rect 56588 31042 56644 31054
rect 56476 30828 56644 30884
rect 56252 28914 56308 28924
rect 56476 30212 56532 30222
rect 55692 28812 55972 28868
rect 55580 28590 55582 28642
rect 55634 28590 55636 28642
rect 55580 28578 55636 28590
rect 55804 28532 55860 28542
rect 55804 28438 55860 28476
rect 55468 27412 55524 27580
rect 55356 27356 55524 27412
rect 55580 28196 55636 28206
rect 55356 27300 55412 27356
rect 55356 27234 55412 27244
rect 55244 27022 55246 27074
rect 55298 27022 55300 27074
rect 55244 27010 55300 27022
rect 55468 27074 55524 27086
rect 55468 27022 55470 27074
rect 55522 27022 55524 27074
rect 55468 26908 55524 27022
rect 55580 27074 55636 28140
rect 55580 27022 55582 27074
rect 55634 27022 55636 27074
rect 55580 27010 55636 27022
rect 55692 27970 55748 27982
rect 55692 27918 55694 27970
rect 55746 27918 55748 27970
rect 55692 26908 55748 27918
rect 55804 27858 55860 27870
rect 55804 27806 55806 27858
rect 55858 27806 55860 27858
rect 55804 27300 55860 27806
rect 55804 27074 55860 27244
rect 55804 27022 55806 27074
rect 55858 27022 55860 27074
rect 55804 27010 55860 27022
rect 55132 26852 55300 26908
rect 55468 26852 55748 26908
rect 55132 26292 55188 26302
rect 54908 25666 54964 25676
rect 55020 26236 55132 26292
rect 54908 25508 54964 25518
rect 55020 25508 55076 26236
rect 55132 26226 55188 26236
rect 55132 25620 55188 25630
rect 55132 25526 55188 25564
rect 54908 25506 55076 25508
rect 54908 25454 54910 25506
rect 54962 25454 55076 25506
rect 54908 25452 55076 25454
rect 54908 25442 54964 25452
rect 55132 25396 55188 25406
rect 55132 24724 55188 25340
rect 55244 24834 55300 26852
rect 55580 26628 55636 26852
rect 55580 26562 55636 26572
rect 55804 26404 55860 26414
rect 55692 26348 55804 26404
rect 55244 24782 55246 24834
rect 55298 24782 55300 24834
rect 55244 24770 55300 24782
rect 55356 26178 55412 26190
rect 55356 26126 55358 26178
rect 55410 26126 55412 26178
rect 54796 24210 54852 24220
rect 54908 24722 55188 24724
rect 54908 24670 55134 24722
rect 55186 24670 55188 24722
rect 54908 24668 55188 24670
rect 54908 24050 54964 24668
rect 55132 24658 55188 24668
rect 54908 23998 54910 24050
rect 54962 23998 54964 24050
rect 54908 23986 54964 23998
rect 54796 23940 54852 23950
rect 54684 23884 54796 23940
rect 54796 23846 54852 23884
rect 53788 22370 53844 23660
rect 54236 23716 54292 23726
rect 54236 22482 54292 23660
rect 54236 22430 54238 22482
rect 54290 22430 54292 22482
rect 54236 22418 54292 22430
rect 54348 23380 54404 23390
rect 53788 22318 53790 22370
rect 53842 22318 53844 22370
rect 53788 22306 53844 22318
rect 54348 22370 54404 23324
rect 54572 23268 54628 23278
rect 54572 23154 54628 23212
rect 54572 23102 54574 23154
rect 54626 23102 54628 23154
rect 54572 23090 54628 23102
rect 54796 23044 54852 23054
rect 54796 22950 54852 22988
rect 54348 22318 54350 22370
rect 54402 22318 54404 22370
rect 54348 22306 54404 22318
rect 54012 22258 54068 22270
rect 55132 22260 55188 22270
rect 54012 22206 54014 22258
rect 54066 22206 54068 22258
rect 54012 21924 54068 22206
rect 54012 21858 54068 21868
rect 54460 22258 55188 22260
rect 54460 22206 55134 22258
rect 55186 22206 55188 22258
rect 54460 22204 55188 22206
rect 54460 21588 54516 22204
rect 55132 22194 55188 22204
rect 55356 22036 55412 26126
rect 55692 25620 55748 26348
rect 55804 26310 55860 26348
rect 55692 25554 55748 25564
rect 55804 25506 55860 25518
rect 55804 25454 55806 25506
rect 55858 25454 55860 25506
rect 55468 25282 55524 25294
rect 55468 25230 55470 25282
rect 55522 25230 55524 25282
rect 55468 24722 55524 25230
rect 55468 24670 55470 24722
rect 55522 24670 55524 24722
rect 55468 24658 55524 24670
rect 55692 24276 55748 24286
rect 55020 21980 55412 22036
rect 55468 23940 55524 23950
rect 54236 21532 54516 21588
rect 54684 21586 54740 21598
rect 54684 21534 54686 21586
rect 54738 21534 54740 21586
rect 53452 21298 53508 21308
rect 53564 21308 53676 21364
rect 53116 20862 53118 20914
rect 53170 20862 53172 20914
rect 53116 20850 53172 20862
rect 53116 19794 53172 19806
rect 53116 19742 53118 19794
rect 53170 19742 53172 19794
rect 53116 19124 53172 19742
rect 53564 19460 53620 21308
rect 53676 21298 53732 21308
rect 53900 21476 53956 21486
rect 53900 20802 53956 21420
rect 53900 20750 53902 20802
rect 53954 20750 53956 20802
rect 53900 20738 53956 20750
rect 54012 21474 54068 21486
rect 54012 21422 54014 21474
rect 54066 21422 54068 21474
rect 54012 21252 54068 21422
rect 54012 20802 54068 21196
rect 54012 20750 54014 20802
rect 54066 20750 54068 20802
rect 54012 20738 54068 20750
rect 54124 21362 54180 21374
rect 54124 21310 54126 21362
rect 54178 21310 54180 21362
rect 54124 20804 54180 21310
rect 54236 20914 54292 21532
rect 54460 21364 54516 21374
rect 54460 21270 54516 21308
rect 54684 21252 54740 21534
rect 55020 21588 55076 21980
rect 55356 21812 55412 21822
rect 55356 21718 55412 21756
rect 55020 21494 55076 21532
rect 55244 21700 55300 21710
rect 55244 21586 55300 21644
rect 55244 21534 55246 21586
rect 55298 21534 55300 21586
rect 55244 21522 55300 21534
rect 54684 21186 54740 21196
rect 54236 20862 54238 20914
rect 54290 20862 54292 20914
rect 54236 20850 54292 20862
rect 54348 20916 54404 20926
rect 54124 20738 54180 20748
rect 53900 20130 53956 20142
rect 53900 20078 53902 20130
rect 53954 20078 53956 20130
rect 53676 20020 53732 20030
rect 53676 19926 53732 19964
rect 53900 19796 53956 20078
rect 54348 20130 54404 20860
rect 54348 20078 54350 20130
rect 54402 20078 54404 20130
rect 54348 20066 54404 20078
rect 54460 20802 54516 20814
rect 54460 20750 54462 20802
rect 54514 20750 54516 20802
rect 54460 20132 54516 20750
rect 54460 20066 54516 20076
rect 54572 20692 54628 20702
rect 54572 20130 54628 20636
rect 54572 20078 54574 20130
rect 54626 20078 54628 20130
rect 54572 20066 54628 20078
rect 55020 20244 55076 20254
rect 55020 20018 55076 20188
rect 55020 19966 55022 20018
rect 55074 19966 55076 20018
rect 55020 19954 55076 19966
rect 54460 19906 54516 19918
rect 54460 19854 54462 19906
rect 54514 19854 54516 19906
rect 54460 19796 54516 19854
rect 53900 19740 54516 19796
rect 54572 19908 54628 19918
rect 53452 19404 53620 19460
rect 53116 19058 53172 19068
rect 53228 19346 53284 19358
rect 53228 19294 53230 19346
rect 53282 19294 53284 19346
rect 53228 19012 53284 19294
rect 53116 18450 53172 18462
rect 53116 18398 53118 18450
rect 53170 18398 53172 18450
rect 53116 18340 53172 18398
rect 53228 18452 53284 18956
rect 53340 18452 53396 18462
rect 53228 18450 53396 18452
rect 53228 18398 53342 18450
rect 53394 18398 53396 18450
rect 53228 18396 53396 18398
rect 53116 17556 53172 18284
rect 53340 18228 53396 18396
rect 53340 18162 53396 18172
rect 53228 17556 53284 17566
rect 53116 17500 53228 17556
rect 53228 17462 53284 17500
rect 53004 17276 53284 17332
rect 51884 16436 51940 16446
rect 51548 15922 51604 15932
rect 51772 16324 51828 16334
rect 50988 15428 51044 15438
rect 50988 15334 51044 15372
rect 51212 15426 51268 15484
rect 51212 15374 51214 15426
rect 51266 15374 51268 15426
rect 51212 15362 51268 15374
rect 51548 15428 51604 15438
rect 51548 15334 51604 15372
rect 51660 14306 51716 14318
rect 51660 14254 51662 14306
rect 51714 14254 51716 14306
rect 51660 14196 51716 14254
rect 51548 14140 51660 14196
rect 50540 13020 50932 13076
rect 50540 12850 50596 13020
rect 50540 12798 50542 12850
rect 50594 12798 50596 12850
rect 50540 12786 50596 12798
rect 50652 12852 50708 12862
rect 50652 12758 50708 12796
rect 50316 12738 50372 12750
rect 50316 12686 50318 12738
rect 50370 12686 50372 12738
rect 50316 12516 50372 12686
rect 50428 12740 50484 12750
rect 50428 12646 50484 12684
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50316 12450 50372 12460
rect 50540 12178 50596 12190
rect 50540 12126 50542 12178
rect 50594 12126 50596 12178
rect 50540 11618 50596 12126
rect 50540 11566 50542 11618
rect 50594 11566 50596 11618
rect 50540 11554 50596 11566
rect 50876 11394 50932 13020
rect 50988 13746 51044 13758
rect 50988 13694 50990 13746
rect 51042 13694 51044 13746
rect 50988 12962 51044 13694
rect 51212 13748 51268 13758
rect 51436 13748 51492 13758
rect 51212 13746 51492 13748
rect 51212 13694 51214 13746
rect 51266 13694 51438 13746
rect 51490 13694 51492 13746
rect 51212 13692 51492 13694
rect 51212 13682 51268 13692
rect 51436 13682 51492 13692
rect 50988 12910 50990 12962
rect 51042 12910 51044 12962
rect 50988 12898 51044 12910
rect 51436 13076 51492 13086
rect 51548 13076 51604 14140
rect 51660 14130 51716 14140
rect 51772 13746 51828 16268
rect 51884 16210 51940 16380
rect 51884 16158 51886 16210
rect 51938 16158 51940 16210
rect 51884 16146 51940 16158
rect 51884 15314 51940 15326
rect 51884 15262 51886 15314
rect 51938 15262 51940 15314
rect 51884 15204 51940 15262
rect 51884 15138 51940 15148
rect 51996 15148 52052 16828
rect 53004 16770 53060 16782
rect 53004 16718 53006 16770
rect 53058 16718 53060 16770
rect 53004 15988 53060 16718
rect 53116 15988 53172 15998
rect 53004 15986 53172 15988
rect 53004 15934 53118 15986
rect 53170 15934 53172 15986
rect 53004 15932 53172 15934
rect 52780 15874 52836 15886
rect 52780 15822 52782 15874
rect 52834 15822 52836 15874
rect 52780 15540 52836 15822
rect 53116 15876 53172 15932
rect 53116 15810 53172 15820
rect 52780 15474 52836 15484
rect 53116 15428 53172 15438
rect 52332 15204 52388 15242
rect 51996 15092 52164 15148
rect 52332 15138 52388 15148
rect 51996 14308 52052 14318
rect 51772 13694 51774 13746
rect 51826 13694 51828 13746
rect 51772 13682 51828 13694
rect 51884 14306 52052 14308
rect 51884 14254 51998 14306
rect 52050 14254 52052 14306
rect 51884 14252 52052 14254
rect 51436 13074 51604 13076
rect 51436 13022 51438 13074
rect 51490 13022 51604 13074
rect 51436 13020 51604 13022
rect 51212 12292 51268 12302
rect 51212 12198 51268 12236
rect 51436 11508 51492 13020
rect 51660 12964 51716 12974
rect 51660 12962 51828 12964
rect 51660 12910 51662 12962
rect 51714 12910 51828 12962
rect 51660 12908 51828 12910
rect 51660 12898 51716 12908
rect 51100 11452 51492 11508
rect 50876 11342 50878 11394
rect 50930 11342 50932 11394
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50428 10610 50484 10622
rect 50428 10558 50430 10610
rect 50482 10558 50484 10610
rect 50428 10164 50484 10558
rect 50428 10050 50484 10108
rect 50428 9998 50430 10050
rect 50482 9998 50484 10050
rect 50428 8148 50484 9998
rect 50652 10612 50708 10622
rect 50652 9714 50708 10556
rect 50652 9662 50654 9714
rect 50706 9662 50708 9714
rect 50652 9650 50708 9662
rect 50876 9716 50932 11342
rect 50876 9650 50932 9660
rect 50988 11396 51044 11406
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50988 9156 51044 11340
rect 51100 11394 51156 11452
rect 51100 11342 51102 11394
rect 51154 11342 51156 11394
rect 51100 11330 51156 11342
rect 51772 11394 51828 12908
rect 51772 11342 51774 11394
rect 51826 11342 51828 11394
rect 51212 11172 51268 11182
rect 51212 9714 51268 11116
rect 51436 11170 51492 11182
rect 51436 11118 51438 11170
rect 51490 11118 51492 11170
rect 51436 11060 51492 11118
rect 51436 10994 51492 11004
rect 51772 9828 51828 11342
rect 51772 9762 51828 9772
rect 51212 9662 51214 9714
rect 51266 9662 51268 9714
rect 51212 9650 51268 9662
rect 51660 9716 51716 9726
rect 51660 9622 51716 9660
rect 51436 9156 51492 9166
rect 50988 9154 51492 9156
rect 50988 9102 51438 9154
rect 51490 9102 51492 9154
rect 50988 9100 51492 9102
rect 51436 9090 51492 9100
rect 51548 9044 51604 9054
rect 51548 8428 51604 8988
rect 51436 8372 51604 8428
rect 51660 9042 51716 9054
rect 51660 8990 51662 9042
rect 51714 8990 51716 9042
rect 51436 8370 51492 8372
rect 51436 8318 51438 8370
rect 51490 8318 51492 8370
rect 51436 8306 51492 8318
rect 50428 8082 50484 8092
rect 49980 6526 49982 6578
rect 50034 6526 50036 6578
rect 49980 6514 50036 6526
rect 50092 7308 50204 7364
rect 49532 6402 49588 6412
rect 49420 6244 49476 6254
rect 49420 6130 49476 6188
rect 49420 6078 49422 6130
rect 49474 6078 49476 6130
rect 49420 6066 49476 6078
rect 49980 6132 50036 6142
rect 50092 6132 50148 7308
rect 50204 7298 50260 7308
rect 50316 8034 50372 8046
rect 50316 7982 50318 8034
rect 50370 7982 50372 8034
rect 50316 6692 50372 7982
rect 51660 8036 51716 8990
rect 51884 8428 51940 14252
rect 51996 14242 52052 14252
rect 52108 13972 52164 15092
rect 53116 14754 53172 15372
rect 53116 14702 53118 14754
rect 53170 14702 53172 14754
rect 53116 14690 53172 14702
rect 52892 14418 52948 14430
rect 52892 14366 52894 14418
rect 52946 14366 52948 14418
rect 52892 14196 52948 14366
rect 52892 14130 52948 14140
rect 51996 12738 52052 12750
rect 51996 12686 51998 12738
rect 52050 12686 52052 12738
rect 51996 11396 52052 12686
rect 51996 11330 52052 11340
rect 51996 9828 52052 9838
rect 51996 9734 52052 9772
rect 51660 7970 51716 7980
rect 51772 8372 51940 8428
rect 51996 8372 52052 8382
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 51660 7700 51716 7710
rect 51660 7606 51716 7644
rect 51100 7476 51156 7486
rect 51100 7362 51156 7420
rect 51100 7310 51102 7362
rect 51154 7310 51156 7362
rect 49980 6130 50148 6132
rect 49980 6078 49982 6130
rect 50034 6078 50148 6130
rect 49980 6076 50148 6078
rect 50204 6690 50372 6692
rect 50204 6638 50318 6690
rect 50370 6638 50372 6690
rect 50204 6636 50372 6638
rect 49980 6066 50036 6076
rect 49644 5682 49700 5694
rect 49644 5630 49646 5682
rect 49698 5630 49700 5682
rect 49644 5234 49700 5630
rect 50204 5682 50260 6636
rect 50316 6626 50372 6636
rect 50764 6692 50820 6702
rect 50764 6598 50820 6636
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50316 6132 50372 6142
rect 50316 6038 50372 6076
rect 50204 5630 50206 5682
rect 50258 5630 50260 5682
rect 50204 5618 50260 5630
rect 50764 5794 50820 5806
rect 50764 5742 50766 5794
rect 50818 5742 50820 5794
rect 49644 5182 49646 5234
rect 49698 5182 49700 5234
rect 49644 5170 49700 5182
rect 50764 5236 50820 5742
rect 50764 5170 50820 5180
rect 50204 5124 50260 5134
rect 50204 5030 50260 5068
rect 51100 5124 51156 7310
rect 51212 7140 51268 7150
rect 51212 6690 51268 7084
rect 51212 6638 51214 6690
rect 51266 6638 51268 6690
rect 51212 6626 51268 6638
rect 51660 7028 51716 7038
rect 51660 6690 51716 6972
rect 51660 6638 51662 6690
rect 51714 6638 51716 6690
rect 51660 6626 51716 6638
rect 51100 5058 51156 5068
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 48972 4562 49364 4564
rect 48972 4510 48974 4562
rect 49026 4510 49364 4562
rect 48972 4508 49364 4510
rect 48972 4498 49028 4508
rect 48524 3574 48580 3612
rect 49308 4228 49364 4238
rect 46844 3490 46900 3500
rect 47516 3556 47572 3566
rect 47516 3462 47572 3500
rect 49308 3556 49364 4172
rect 49308 3490 49364 3500
rect 51772 3332 51828 8372
rect 51996 8278 52052 8316
rect 52108 7698 52164 13916
rect 52332 13860 52388 13870
rect 52332 13766 52388 13804
rect 52556 13748 52612 13758
rect 52556 13654 52612 13692
rect 53004 12738 53060 12750
rect 53004 12686 53006 12738
rect 53058 12686 53060 12738
rect 52668 12292 52724 12302
rect 53004 12292 53060 12686
rect 52668 12290 53060 12292
rect 52668 12238 52670 12290
rect 52722 12238 53060 12290
rect 52668 12236 53060 12238
rect 52220 12178 52276 12190
rect 52220 12126 52222 12178
rect 52274 12126 52276 12178
rect 52220 11060 52276 12126
rect 52220 10994 52276 11004
rect 52668 11170 52724 12236
rect 53004 12068 53060 12078
rect 52668 11118 52670 11170
rect 52722 11118 52724 11170
rect 52668 10948 52724 11118
rect 52780 11172 52836 11182
rect 52780 11078 52836 11116
rect 52892 11170 52948 11182
rect 52892 11118 52894 11170
rect 52946 11118 52948 11170
rect 52892 11060 52948 11118
rect 52892 10994 52948 11004
rect 52668 10892 52836 10948
rect 52444 10612 52500 10622
rect 52668 10612 52724 10622
rect 52500 10610 52724 10612
rect 52500 10558 52670 10610
rect 52722 10558 52724 10610
rect 52500 10556 52724 10558
rect 52444 10546 52500 10556
rect 52556 10388 52612 10398
rect 52556 10294 52612 10332
rect 52668 9268 52724 10556
rect 52780 10612 52836 10892
rect 52780 10546 52836 10556
rect 53004 10052 53060 12012
rect 53116 11396 53172 11406
rect 53116 11282 53172 11340
rect 53116 11230 53118 11282
rect 53170 11230 53172 11282
rect 53116 10722 53172 11230
rect 53116 10670 53118 10722
rect 53170 10670 53172 10722
rect 53116 10658 53172 10670
rect 52892 9996 53060 10052
rect 52780 9828 52836 9838
rect 52780 9734 52836 9772
rect 52780 9268 52836 9278
rect 52668 9266 52836 9268
rect 52668 9214 52782 9266
rect 52834 9214 52836 9266
rect 52668 9212 52836 9214
rect 52780 9202 52836 9212
rect 52668 9044 52724 9054
rect 52668 8950 52724 8988
rect 52892 8370 52948 9996
rect 53228 8428 53284 17276
rect 53340 16996 53396 17006
rect 53340 14308 53396 16940
rect 53452 16212 53508 19404
rect 53564 19234 53620 19246
rect 53564 19182 53566 19234
rect 53618 19182 53620 19234
rect 53564 18340 53620 19182
rect 54348 19234 54404 19246
rect 54348 19182 54350 19234
rect 54402 19182 54404 19234
rect 54348 19124 54404 19182
rect 54236 19068 54348 19124
rect 53676 18900 53732 18910
rect 53676 18562 53732 18844
rect 53788 18676 53844 18686
rect 53788 18582 53844 18620
rect 53676 18510 53678 18562
rect 53730 18510 53732 18562
rect 53676 18498 53732 18510
rect 54012 18562 54068 18574
rect 54012 18510 54014 18562
rect 54066 18510 54068 18562
rect 54012 18452 54068 18510
rect 54124 18452 54180 18462
rect 54012 18450 54180 18452
rect 54012 18398 54126 18450
rect 54178 18398 54180 18450
rect 54012 18396 54180 18398
rect 54124 18386 54180 18396
rect 53564 17892 53620 18284
rect 53564 17826 53620 17836
rect 53676 18004 53732 18014
rect 53676 17554 53732 17948
rect 53788 17780 53844 17790
rect 53788 17668 53844 17724
rect 53788 17666 53956 17668
rect 53788 17614 53790 17666
rect 53842 17614 53956 17666
rect 53788 17612 53956 17614
rect 53788 17602 53844 17612
rect 53676 17502 53678 17554
rect 53730 17502 53732 17554
rect 53676 17490 53732 17502
rect 53788 17108 53844 17118
rect 53452 16146 53508 16156
rect 53676 16882 53732 16894
rect 53676 16830 53678 16882
rect 53730 16830 53732 16882
rect 53452 15988 53508 15998
rect 53452 14754 53508 15932
rect 53564 15428 53620 15438
rect 53564 15334 53620 15372
rect 53676 15204 53732 16830
rect 53676 15138 53732 15148
rect 53452 14702 53454 14754
rect 53506 14702 53508 14754
rect 53452 14690 53508 14702
rect 53340 14242 53396 14252
rect 53340 13748 53396 13758
rect 53788 13748 53844 17052
rect 53900 14754 53956 17612
rect 54236 17666 54292 19068
rect 54348 19058 54404 19068
rect 54348 18228 54404 18238
rect 54348 18134 54404 18172
rect 54236 17614 54238 17666
rect 54290 17614 54292 17666
rect 53900 14702 53902 14754
rect 53954 14702 53956 14754
rect 53900 14690 53956 14702
rect 54012 16100 54068 16110
rect 53396 13692 53844 13748
rect 53900 14420 53956 14430
rect 53340 13654 53396 13692
rect 53900 13634 53956 14364
rect 53900 13582 53902 13634
rect 53954 13582 53956 13634
rect 53900 13570 53956 13582
rect 54012 14084 54068 16044
rect 53788 13524 53844 13534
rect 53340 13076 53396 13086
rect 53340 12982 53396 13020
rect 53340 12740 53396 12750
rect 53340 12290 53396 12684
rect 53340 12238 53342 12290
rect 53394 12238 53396 12290
rect 53340 12226 53396 12238
rect 52892 8318 52894 8370
rect 52946 8318 52948 8370
rect 52892 8306 52948 8318
rect 53004 8372 53284 8428
rect 53340 9268 53396 9278
rect 53004 8306 53060 8316
rect 53340 8370 53396 9212
rect 53676 8930 53732 8942
rect 53676 8878 53678 8930
rect 53730 8878 53732 8930
rect 53676 8820 53732 8878
rect 53676 8754 53732 8764
rect 53340 8318 53342 8370
rect 53394 8318 53396 8370
rect 53340 8306 53396 8318
rect 53788 8370 53844 13468
rect 54012 13412 54068 14028
rect 53900 13356 54068 13412
rect 54236 13412 54292 17614
rect 54460 17556 54516 17566
rect 54572 17556 54628 19852
rect 55468 19906 55524 23884
rect 55468 19854 55470 19906
rect 55522 19854 55524 19906
rect 55468 19842 55524 19854
rect 55580 23044 55636 23054
rect 54684 19236 54740 19246
rect 54684 17666 54740 19180
rect 54908 18452 54964 18462
rect 54908 18358 54964 18396
rect 55580 18116 55636 22988
rect 55692 21810 55748 24220
rect 55692 21758 55694 21810
rect 55746 21758 55748 21810
rect 55692 21746 55748 21758
rect 55804 22372 55860 25454
rect 55916 22484 55972 28812
rect 56252 28756 56308 28766
rect 56252 28662 56308 28700
rect 56476 28532 56532 30156
rect 56588 29426 56644 30828
rect 56700 30434 56756 35532
rect 57260 35364 57316 35646
rect 57260 35298 57316 35308
rect 56812 35252 56868 35262
rect 56812 34692 56868 35196
rect 57484 35252 57540 36876
rect 58380 36260 58436 37102
rect 58380 35924 58436 36204
rect 58156 35922 58436 35924
rect 58156 35870 58382 35922
rect 58434 35870 58436 35922
rect 58156 35868 58436 35870
rect 57484 35186 57540 35196
rect 58044 35474 58100 35486
rect 58044 35422 58046 35474
rect 58098 35422 58100 35474
rect 58044 35140 58100 35422
rect 58044 35074 58100 35084
rect 56924 34916 56980 34926
rect 56924 34822 56980 34860
rect 58044 34916 58100 34926
rect 58156 34916 58212 35868
rect 58380 35858 58436 35868
rect 58492 36036 58548 37214
rect 58044 34914 58212 34916
rect 58044 34862 58046 34914
rect 58098 34862 58212 34914
rect 58044 34860 58212 34862
rect 58268 34916 58324 34926
rect 58492 34916 58548 35980
rect 58828 35700 58884 35710
rect 58828 35606 58884 35644
rect 58268 34914 58548 34916
rect 58268 34862 58270 34914
rect 58322 34862 58548 34914
rect 58268 34860 58548 34862
rect 58716 35140 58772 35150
rect 58044 34850 58100 34860
rect 57148 34802 57204 34814
rect 57148 34750 57150 34802
rect 57202 34750 57204 34802
rect 56924 34692 56980 34702
rect 56812 34636 56924 34692
rect 56812 33348 56868 33358
rect 56812 33254 56868 33292
rect 56812 32788 56868 32798
rect 56812 32116 56868 32732
rect 56924 32450 56980 34636
rect 57036 34580 57092 34590
rect 57036 34242 57092 34524
rect 57148 34356 57204 34750
rect 58268 34692 58324 34860
rect 58268 34626 58324 34636
rect 57148 34290 57204 34300
rect 57036 34190 57038 34242
rect 57090 34190 57092 34242
rect 57036 34178 57092 34190
rect 57036 33908 57092 33918
rect 57036 32562 57092 33852
rect 58716 33908 58772 35084
rect 59052 34356 59108 37436
rect 59276 36820 59332 38556
rect 59500 38164 59556 38174
rect 59500 38050 59556 38108
rect 59500 37998 59502 38050
rect 59554 37998 59556 38050
rect 59500 37492 59556 37998
rect 59500 37426 59556 37436
rect 59612 37938 59668 37950
rect 59612 37886 59614 37938
rect 59666 37886 59668 37938
rect 59276 36370 59332 36764
rect 59276 36318 59278 36370
rect 59330 36318 59332 36370
rect 59276 36306 59332 36318
rect 59500 37156 59556 37166
rect 59500 35812 59556 37100
rect 59612 37044 59668 37886
rect 59612 36978 59668 36988
rect 60060 37378 60116 37390
rect 60060 37326 60062 37378
rect 60114 37326 60116 37378
rect 60060 36484 60116 37326
rect 60060 36418 60116 36428
rect 59612 35812 59668 35822
rect 59500 35810 59668 35812
rect 59500 35758 59614 35810
rect 59666 35758 59668 35810
rect 59500 35756 59668 35758
rect 59612 35746 59668 35756
rect 59612 34916 59668 34926
rect 59612 34802 59668 34860
rect 59612 34750 59614 34802
rect 59666 34750 59668 34802
rect 59612 34738 59668 34750
rect 59836 34914 59892 34926
rect 59836 34862 59838 34914
rect 59890 34862 59892 34914
rect 59164 34356 59220 34366
rect 59052 34354 59220 34356
rect 59052 34302 59166 34354
rect 59218 34302 59220 34354
rect 59052 34300 59220 34302
rect 59164 34290 59220 34300
rect 59388 34244 59444 34254
rect 58828 33908 58884 33918
rect 58716 33906 58884 33908
rect 58716 33854 58830 33906
rect 58882 33854 58884 33906
rect 58716 33852 58884 33854
rect 57036 32510 57038 32562
rect 57090 32510 57092 32562
rect 57036 32498 57092 32510
rect 57148 33572 57204 33582
rect 56924 32398 56926 32450
rect 56978 32398 56980 32450
rect 56924 32386 56980 32398
rect 56812 31220 56868 32060
rect 57148 32002 57204 33516
rect 58156 33348 58212 33358
rect 57484 32788 57540 32798
rect 57484 32694 57540 32732
rect 57596 32732 57876 32788
rect 57596 32564 57652 32732
rect 57820 32676 57876 32732
rect 57932 32676 57988 32686
rect 57820 32674 57988 32676
rect 57820 32622 57934 32674
rect 57986 32622 57988 32674
rect 57820 32620 57988 32622
rect 57932 32610 57988 32620
rect 57148 31950 57150 32002
rect 57202 31950 57204 32002
rect 57148 31938 57204 31950
rect 57260 32508 57652 32564
rect 57708 32562 57764 32574
rect 57708 32510 57710 32562
rect 57762 32510 57764 32562
rect 57148 31556 57204 31566
rect 56812 31164 56980 31220
rect 56700 30382 56702 30434
rect 56754 30382 56756 30434
rect 56700 30370 56756 30382
rect 56812 30994 56868 31006
rect 56812 30942 56814 30994
rect 56866 30942 56868 30994
rect 56812 30436 56868 30942
rect 56812 30370 56868 30380
rect 56924 30210 56980 31164
rect 57036 30882 57092 30894
rect 57036 30830 57038 30882
rect 57090 30830 57092 30882
rect 57036 30324 57092 30830
rect 57036 30258 57092 30268
rect 56924 30158 56926 30210
rect 56978 30158 56980 30210
rect 56924 30100 56980 30158
rect 57148 30100 57204 31500
rect 56924 30034 56980 30044
rect 57036 30044 57204 30100
rect 57260 30994 57316 32508
rect 57260 30942 57262 30994
rect 57314 30942 57316 30994
rect 56588 29374 56590 29426
rect 56642 29374 56644 29426
rect 56588 29092 56644 29374
rect 56700 29538 56756 29550
rect 56700 29486 56702 29538
rect 56754 29486 56756 29538
rect 56700 29428 56756 29486
rect 56700 29362 56756 29372
rect 56924 29540 56980 29550
rect 56700 29204 56756 29214
rect 56700 29202 56868 29204
rect 56700 29150 56702 29202
rect 56754 29150 56868 29202
rect 56700 29148 56868 29150
rect 56700 29138 56756 29148
rect 56588 29026 56644 29036
rect 56588 28868 56644 28878
rect 56644 28812 56756 28868
rect 56588 28802 56644 28812
rect 56476 28466 56532 28476
rect 56588 28642 56644 28654
rect 56588 28590 56590 28642
rect 56642 28590 56644 28642
rect 56476 28308 56532 28318
rect 56252 28252 56476 28308
rect 56028 26292 56084 26302
rect 56028 26068 56084 26236
rect 56028 26002 56084 26012
rect 56028 25844 56084 25854
rect 56028 25506 56084 25788
rect 56028 25454 56030 25506
rect 56082 25454 56084 25506
rect 56028 23044 56084 25454
rect 56028 22978 56084 22988
rect 55916 22428 56196 22484
rect 55804 21588 55860 22316
rect 56028 22260 56084 22270
rect 55916 21588 55972 21598
rect 55804 21586 55972 21588
rect 55804 21534 55918 21586
rect 55970 21534 55972 21586
rect 55804 21532 55972 21534
rect 55804 21028 55860 21038
rect 55692 20802 55748 20814
rect 55692 20750 55694 20802
rect 55746 20750 55748 20802
rect 55692 20020 55748 20750
rect 55692 19234 55748 19964
rect 55692 19182 55694 19234
rect 55746 19182 55748 19234
rect 55692 18228 55748 19182
rect 55804 19124 55860 20972
rect 55916 20018 55972 21532
rect 55916 19966 55918 20018
rect 55970 19966 55972 20018
rect 55916 19954 55972 19966
rect 55804 19058 55860 19068
rect 56028 18676 56084 22204
rect 56140 20802 56196 22428
rect 56252 20916 56308 28252
rect 56476 28242 56532 28252
rect 56364 28084 56420 28094
rect 56364 23940 56420 28028
rect 56588 27524 56644 28590
rect 56700 28420 56756 28812
rect 56812 28644 56868 29148
rect 56812 28578 56868 28588
rect 56700 28364 56868 28420
rect 56812 28082 56868 28364
rect 56812 28030 56814 28082
rect 56866 28030 56868 28082
rect 56812 27860 56868 28030
rect 56924 28082 56980 29484
rect 57036 28308 57092 30044
rect 57260 29764 57316 30942
rect 57372 32338 57428 32350
rect 57372 32286 57374 32338
rect 57426 32286 57428 32338
rect 57372 30210 57428 32286
rect 57484 31892 57540 31902
rect 57484 31798 57540 31836
rect 57596 31556 57652 31566
rect 57596 31218 57652 31500
rect 57596 31166 57598 31218
rect 57650 31166 57652 31218
rect 57596 31154 57652 31166
rect 57372 30158 57374 30210
rect 57426 30158 57428 30210
rect 57372 30146 57428 30158
rect 57708 30436 57764 32510
rect 57820 31780 57876 31790
rect 57820 30996 57876 31724
rect 57932 31332 57988 31342
rect 57988 31276 58100 31332
rect 57932 31266 57988 31276
rect 57932 30996 57988 31006
rect 57820 30994 57988 30996
rect 57820 30942 57934 30994
rect 57986 30942 57988 30994
rect 57820 30940 57988 30942
rect 57932 30930 57988 30940
rect 58044 30660 58100 31276
rect 58156 31106 58212 33292
rect 58380 32788 58436 32798
rect 58380 32786 58660 32788
rect 58380 32734 58382 32786
rect 58434 32734 58660 32786
rect 58380 32732 58660 32734
rect 58380 32722 58436 32732
rect 58492 32564 58548 32574
rect 58492 32470 58548 32508
rect 58380 32340 58436 32350
rect 58156 31054 58158 31106
rect 58210 31054 58212 31106
rect 58156 31042 58212 31054
rect 58268 32338 58436 32340
rect 58268 32286 58382 32338
rect 58434 32286 58436 32338
rect 58268 32284 58436 32286
rect 58044 30604 58212 30660
rect 57260 29708 57428 29764
rect 57260 29204 57316 29214
rect 57260 29110 57316 29148
rect 57148 28754 57204 28766
rect 57148 28702 57150 28754
rect 57202 28702 57204 28754
rect 57148 28420 57204 28702
rect 57148 28354 57204 28364
rect 57372 28642 57428 29708
rect 57596 29428 57652 29438
rect 57596 29334 57652 29372
rect 57372 28590 57374 28642
rect 57426 28590 57428 28642
rect 57036 28242 57092 28252
rect 56924 28030 56926 28082
rect 56978 28030 56980 28082
rect 56924 28018 56980 28030
rect 57036 27970 57092 27982
rect 57036 27918 57038 27970
rect 57090 27918 57092 27970
rect 56812 27804 56980 27860
rect 56476 27468 56644 27524
rect 56476 26964 56532 27468
rect 56812 27300 56868 27310
rect 56812 27186 56868 27244
rect 56812 27134 56814 27186
rect 56866 27134 56868 27186
rect 56812 27122 56868 27134
rect 56700 27074 56756 27086
rect 56700 27022 56702 27074
rect 56754 27022 56756 27074
rect 56476 26898 56532 26908
rect 56588 26962 56644 26974
rect 56588 26910 56590 26962
rect 56642 26910 56644 26962
rect 56588 25844 56644 26910
rect 56700 26628 56756 27022
rect 56700 26178 56756 26572
rect 56700 26126 56702 26178
rect 56754 26126 56756 26178
rect 56700 26114 56756 26126
rect 56924 25844 56980 27804
rect 57036 27188 57092 27918
rect 57260 27858 57316 27870
rect 57260 27806 57262 27858
rect 57314 27806 57316 27858
rect 57036 27132 57204 27188
rect 57036 26964 57092 26974
rect 57036 26290 57092 26908
rect 57036 26238 57038 26290
rect 57090 26238 57092 26290
rect 57036 26226 57092 26238
rect 57148 26852 57204 27132
rect 56588 25788 56868 25844
rect 56476 25732 56532 25742
rect 56532 25676 56644 25732
rect 56476 25666 56532 25676
rect 56588 25284 56644 25676
rect 56812 25508 56868 25788
rect 56924 25778 56980 25788
rect 56812 25452 56980 25508
rect 56812 25284 56868 25294
rect 56588 25228 56756 25284
rect 56588 24276 56644 24286
rect 56364 23884 56532 23940
rect 56364 23716 56420 23726
rect 56364 23622 56420 23660
rect 56476 22596 56532 23884
rect 56588 23826 56644 24220
rect 56588 23774 56590 23826
rect 56642 23774 56644 23826
rect 56588 23762 56644 23774
rect 56700 23826 56756 25228
rect 56812 24946 56868 25228
rect 56812 24894 56814 24946
rect 56866 24894 56868 24946
rect 56812 24882 56868 24894
rect 56924 24500 56980 25452
rect 57148 25506 57204 26796
rect 57260 26404 57316 27806
rect 57260 26338 57316 26348
rect 57372 26292 57428 28590
rect 57708 28530 57764 30380
rect 58044 29428 58100 29438
rect 58044 29334 58100 29372
rect 58156 28866 58212 30604
rect 58156 28814 58158 28866
rect 58210 28814 58212 28866
rect 58156 28802 58212 28814
rect 57708 28478 57710 28530
rect 57762 28478 57764 28530
rect 57708 28196 57764 28478
rect 57708 28130 57764 28140
rect 57932 28644 57988 28654
rect 57596 27972 57652 27982
rect 57596 27858 57652 27916
rect 57596 27806 57598 27858
rect 57650 27806 57652 27858
rect 57596 27794 57652 27806
rect 57596 27524 57652 27534
rect 57484 27074 57540 27086
rect 57484 27022 57486 27074
rect 57538 27022 57540 27074
rect 57484 26516 57540 27022
rect 57484 26450 57540 26460
rect 57372 26226 57428 26236
rect 57148 25454 57150 25506
rect 57202 25454 57204 25506
rect 57148 25442 57204 25454
rect 57260 25394 57316 25406
rect 57260 25342 57262 25394
rect 57314 25342 57316 25394
rect 57260 25284 57316 25342
rect 57260 25218 57316 25228
rect 57260 25060 57316 25070
rect 57316 25004 57428 25060
rect 57260 24994 57316 25004
rect 57036 24948 57092 24958
rect 57036 24854 57092 24892
rect 57148 24836 57204 24846
rect 57148 24742 57204 24780
rect 56924 24434 56980 24444
rect 57260 24722 57316 24734
rect 57260 24670 57262 24722
rect 57314 24670 57316 24722
rect 56700 23774 56702 23826
rect 56754 23774 56756 23826
rect 56700 23762 56756 23774
rect 56924 24276 56980 24286
rect 56588 23492 56644 23502
rect 56588 23378 56644 23436
rect 56588 23326 56590 23378
rect 56642 23326 56644 23378
rect 56588 23314 56644 23326
rect 56924 23154 56980 24220
rect 57148 24052 57204 24062
rect 57148 23958 57204 23996
rect 57036 23938 57092 23950
rect 57036 23886 57038 23938
rect 57090 23886 57092 23938
rect 57036 23828 57092 23886
rect 57036 23762 57092 23772
rect 57260 23492 57316 24670
rect 57260 23426 57316 23436
rect 56924 23102 56926 23154
rect 56978 23102 56980 23154
rect 56924 23090 56980 23102
rect 57036 23044 57092 23054
rect 57148 23044 57204 23054
rect 57092 23042 57204 23044
rect 57092 22990 57150 23042
rect 57202 22990 57204 23042
rect 57092 22988 57204 22990
rect 56476 22540 56644 22596
rect 56308 20860 56420 20916
rect 56252 20822 56308 20860
rect 56140 20750 56142 20802
rect 56194 20750 56196 20802
rect 56140 20244 56196 20750
rect 56364 20802 56420 20860
rect 56364 20750 56366 20802
rect 56418 20750 56420 20802
rect 56364 20738 56420 20750
rect 56588 20802 56644 22540
rect 57036 22146 57092 22988
rect 57148 22978 57204 22988
rect 57260 22932 57316 22942
rect 57260 22258 57316 22876
rect 57260 22206 57262 22258
rect 57314 22206 57316 22258
rect 57260 22194 57316 22206
rect 57036 22094 57038 22146
rect 57090 22094 57092 22146
rect 57036 22036 57092 22094
rect 57036 21970 57092 21980
rect 57148 22148 57204 22158
rect 56588 20750 56590 20802
rect 56642 20750 56644 20802
rect 56140 20178 56196 20188
rect 56252 20690 56308 20702
rect 56252 20638 56254 20690
rect 56306 20638 56308 20690
rect 56252 19236 56308 20638
rect 56588 20692 56644 20750
rect 56588 20626 56644 20636
rect 57036 20020 57092 20030
rect 57036 19926 57092 19964
rect 56588 19908 56644 19918
rect 56588 19814 56644 19852
rect 56812 19460 56868 19470
rect 56812 19458 56980 19460
rect 56812 19406 56814 19458
rect 56866 19406 56980 19458
rect 56812 19404 56980 19406
rect 56812 19394 56868 19404
rect 56252 19142 56308 19180
rect 56476 19234 56532 19246
rect 56476 19182 56478 19234
rect 56530 19182 56532 19234
rect 55916 18620 56084 18676
rect 56252 18676 56308 18686
rect 56476 18676 56532 19182
rect 56308 18620 56532 18676
rect 56700 19236 56756 19246
rect 55692 18162 55748 18172
rect 55804 18226 55860 18238
rect 55804 18174 55806 18226
rect 55858 18174 55860 18226
rect 55580 18050 55636 18060
rect 55804 17892 55860 18174
rect 55692 17890 55860 17892
rect 55692 17838 55806 17890
rect 55858 17838 55860 17890
rect 55692 17836 55860 17838
rect 54684 17614 54686 17666
rect 54738 17614 54740 17666
rect 54684 17602 54740 17614
rect 55020 17666 55076 17678
rect 55020 17614 55022 17666
rect 55074 17614 55076 17666
rect 54516 17500 54628 17556
rect 55020 17556 55076 17614
rect 55356 17556 55412 17566
rect 55020 17554 55412 17556
rect 55020 17502 55358 17554
rect 55410 17502 55412 17554
rect 55020 17500 55412 17502
rect 54460 17462 54516 17500
rect 54348 17444 54404 17454
rect 54348 17350 54404 17388
rect 54572 17108 54628 17118
rect 54628 17052 54740 17108
rect 54572 17014 54628 17052
rect 54348 16882 54404 16894
rect 54348 16830 54350 16882
rect 54402 16830 54404 16882
rect 54348 16212 54404 16830
rect 54460 16772 54516 16782
rect 54460 16678 54516 16716
rect 54572 16212 54628 16222
rect 54348 16210 54628 16212
rect 54348 16158 54574 16210
rect 54626 16158 54628 16210
rect 54348 16156 54628 16158
rect 54348 13748 54404 16156
rect 54572 16146 54628 16156
rect 54684 16098 54740 17052
rect 54684 16046 54686 16098
rect 54738 16046 54740 16098
rect 54684 16034 54740 16046
rect 54796 16994 54852 17006
rect 54796 16942 54798 16994
rect 54850 16942 54852 16994
rect 54796 16100 54852 16942
rect 54796 16034 54852 16044
rect 54908 16772 54964 16782
rect 54908 15426 54964 16716
rect 54908 15374 54910 15426
rect 54962 15374 54964 15426
rect 54908 15362 54964 15374
rect 55020 14530 55076 17500
rect 55356 17490 55412 17500
rect 55468 16994 55524 17006
rect 55468 16942 55470 16994
rect 55522 16942 55524 16994
rect 55468 16772 55524 16942
rect 55468 16706 55524 16716
rect 55580 16882 55636 16894
rect 55580 16830 55582 16882
rect 55634 16830 55636 16882
rect 55468 16324 55524 16334
rect 55580 16324 55636 16830
rect 55468 16322 55636 16324
rect 55468 16270 55470 16322
rect 55522 16270 55636 16322
rect 55468 16268 55636 16270
rect 55356 16098 55412 16110
rect 55356 16046 55358 16098
rect 55410 16046 55412 16098
rect 55356 15988 55412 16046
rect 55356 15922 55412 15932
rect 55356 15426 55412 15438
rect 55356 15374 55358 15426
rect 55410 15374 55412 15426
rect 55356 15316 55412 15374
rect 55356 15250 55412 15260
rect 55468 15148 55524 16268
rect 55692 15764 55748 17836
rect 55804 17826 55860 17836
rect 55916 17556 55972 18620
rect 56028 18452 56084 18462
rect 56252 18452 56308 18620
rect 56028 18450 56308 18452
rect 56028 18398 56030 18450
rect 56082 18398 56308 18450
rect 56028 18396 56308 18398
rect 56364 18452 56420 18462
rect 56028 18386 56084 18396
rect 55916 17500 56084 17556
rect 56028 17106 56084 17500
rect 56028 17054 56030 17106
rect 56082 17054 56084 17106
rect 55804 16994 55860 17006
rect 55804 16942 55806 16994
rect 55858 16942 55860 16994
rect 55804 16212 55860 16942
rect 55916 16996 55972 17006
rect 55916 16902 55972 16940
rect 55804 16146 55860 16156
rect 55692 15708 55972 15764
rect 55916 15538 55972 15708
rect 55916 15486 55918 15538
rect 55970 15486 55972 15538
rect 55916 15474 55972 15486
rect 55020 14478 55022 14530
rect 55074 14478 55076 14530
rect 55020 14420 55076 14478
rect 55244 15092 55524 15148
rect 55580 15202 55636 15214
rect 55580 15150 55582 15202
rect 55634 15150 55636 15202
rect 55580 15148 55636 15150
rect 56028 15148 56084 17054
rect 56140 16772 56196 18396
rect 56140 16706 56196 16716
rect 56252 18116 56308 18126
rect 55580 15092 56084 15148
rect 56140 16212 56196 16222
rect 56140 15316 56196 16156
rect 55244 14530 55300 15092
rect 55804 14642 55860 15092
rect 55804 14590 55806 14642
rect 55858 14590 55860 14642
rect 55804 14578 55860 14590
rect 55244 14478 55246 14530
rect 55298 14478 55300 14530
rect 55244 14466 55300 14478
rect 55916 14532 55972 14542
rect 56140 14532 56196 15260
rect 56252 14756 56308 18060
rect 56364 17666 56420 18396
rect 56364 17614 56366 17666
rect 56418 17614 56420 17666
rect 56364 17602 56420 17614
rect 56588 18228 56644 18238
rect 56476 17220 56532 17230
rect 56252 14690 56308 14700
rect 56364 15428 56420 15438
rect 55916 14530 56196 14532
rect 55916 14478 55918 14530
rect 55970 14478 56196 14530
rect 55916 14476 56196 14478
rect 55916 14466 55972 14476
rect 55020 14354 55076 14364
rect 55916 14308 55972 14318
rect 54572 13748 54628 13758
rect 55356 13748 55412 13758
rect 54348 13746 54740 13748
rect 54348 13694 54574 13746
rect 54626 13694 54740 13746
rect 54348 13692 54740 13694
rect 54572 13682 54628 13692
rect 54236 13356 54516 13412
rect 53900 9492 53956 13356
rect 54236 13076 54292 13086
rect 54124 12964 54180 12974
rect 54124 12870 54180 12908
rect 54012 12850 54068 12862
rect 54012 12798 54014 12850
rect 54066 12798 54068 12850
rect 54012 12740 54068 12798
rect 54124 12740 54180 12750
rect 54012 12684 54124 12740
rect 54124 12674 54180 12684
rect 54236 11284 54292 13020
rect 54012 11282 54292 11284
rect 54012 11230 54238 11282
rect 54290 11230 54292 11282
rect 54012 11228 54292 11230
rect 54012 9714 54068 11228
rect 54236 11218 54292 11228
rect 54348 11060 54404 11070
rect 54124 10612 54180 10622
rect 54124 10518 54180 10556
rect 54348 10610 54404 11004
rect 54348 10558 54350 10610
rect 54402 10558 54404 10610
rect 54348 10546 54404 10558
rect 54012 9662 54014 9714
rect 54066 9662 54068 9714
rect 54012 9650 54068 9662
rect 53900 9436 54180 9492
rect 53788 8318 53790 8370
rect 53842 8318 53844 8370
rect 53788 8306 53844 8318
rect 52108 7646 52110 7698
rect 52162 7646 52164 7698
rect 52108 7634 52164 7646
rect 54012 7700 54068 9436
rect 54124 9266 54180 9436
rect 54124 9214 54126 9266
rect 54178 9214 54180 9266
rect 54124 9202 54180 9214
rect 54460 9268 54516 13356
rect 54684 13186 54740 13692
rect 55356 13654 55412 13692
rect 54684 13134 54686 13186
rect 54738 13134 54740 13186
rect 54684 13122 54740 13134
rect 55804 13076 55860 13086
rect 55020 12962 55076 12974
rect 55020 12910 55022 12962
rect 55074 12910 55076 12962
rect 55020 12740 55076 12910
rect 55244 12964 55300 12974
rect 55244 12850 55300 12908
rect 55244 12798 55246 12850
rect 55298 12798 55300 12850
rect 55244 12786 55300 12798
rect 55692 12964 55748 12974
rect 55020 12404 55076 12684
rect 55132 12404 55188 12414
rect 55020 12402 55188 12404
rect 55020 12350 55134 12402
rect 55186 12350 55188 12402
rect 55020 12348 55188 12350
rect 55132 12338 55188 12348
rect 55468 12404 55524 12414
rect 55468 12310 55524 12348
rect 55692 12180 55748 12908
rect 55804 12850 55860 13020
rect 55804 12798 55806 12850
rect 55858 12798 55860 12850
rect 55804 12404 55860 12798
rect 55804 12338 55860 12348
rect 55580 12178 55748 12180
rect 55580 12126 55694 12178
rect 55746 12126 55748 12178
rect 55580 12124 55748 12126
rect 55580 11618 55636 12124
rect 55692 12114 55748 12124
rect 55580 11566 55582 11618
rect 55634 11566 55636 11618
rect 55580 11554 55636 11566
rect 55916 11396 55972 14252
rect 56252 12852 56308 12862
rect 55580 11340 55972 11396
rect 56140 12796 56252 12852
rect 55580 9938 55636 11340
rect 56140 11284 56196 12796
rect 56252 12758 56308 12796
rect 56364 12850 56420 15372
rect 56364 12798 56366 12850
rect 56418 12798 56420 12850
rect 56364 12786 56420 12798
rect 56476 15316 56532 17164
rect 56588 17106 56644 18172
rect 56700 17780 56756 19180
rect 56812 19124 56868 19134
rect 56812 18452 56868 19068
rect 56924 18564 56980 19404
rect 57036 18564 57092 18574
rect 56924 18562 57092 18564
rect 56924 18510 57038 18562
rect 57090 18510 57092 18562
rect 56924 18508 57092 18510
rect 56812 18396 56980 18452
rect 56812 17780 56868 17790
rect 56700 17778 56868 17780
rect 56700 17726 56814 17778
rect 56866 17726 56868 17778
rect 56700 17724 56868 17726
rect 56812 17714 56868 17724
rect 56924 17556 56980 18396
rect 57036 18004 57092 18508
rect 57148 18452 57204 22092
rect 57372 21924 57428 25004
rect 57484 23268 57540 23278
rect 57484 22370 57540 23212
rect 57484 22318 57486 22370
rect 57538 22318 57540 22370
rect 57484 22306 57540 22318
rect 57260 21868 57428 21924
rect 57260 21586 57316 21868
rect 57596 21812 57652 27468
rect 57708 27412 57764 27422
rect 57708 27188 57764 27356
rect 57820 27188 57876 27198
rect 57708 27186 57876 27188
rect 57708 27134 57822 27186
rect 57874 27134 57876 27186
rect 57708 27132 57876 27134
rect 57708 26514 57764 27132
rect 57820 27122 57876 27132
rect 57932 27076 57988 28588
rect 58044 28532 58100 28542
rect 58044 27634 58100 28476
rect 58156 27860 58212 27870
rect 58268 27860 58324 32284
rect 58380 32274 58436 32284
rect 58380 31556 58436 31566
rect 58380 29538 58436 31500
rect 58380 29486 58382 29538
rect 58434 29486 58436 29538
rect 58380 29474 58436 29486
rect 58604 27972 58660 32732
rect 58716 31106 58772 33852
rect 58828 33842 58884 33852
rect 59388 33234 59444 34188
rect 59612 33908 59668 33918
rect 59836 33908 59892 34862
rect 59668 33852 59892 33908
rect 59612 33814 59668 33852
rect 59388 33182 59390 33234
rect 59442 33182 59444 33234
rect 59388 33170 59444 33182
rect 60172 32562 60228 45054
rect 60732 45106 60788 45118
rect 60732 45054 60734 45106
rect 60786 45054 60788 45106
rect 60284 44996 60340 45006
rect 60340 44940 60452 44996
rect 60284 44930 60340 44940
rect 60396 42756 60452 44940
rect 60620 44772 60676 44782
rect 60620 44546 60676 44716
rect 60620 44494 60622 44546
rect 60674 44494 60676 44546
rect 60620 44482 60676 44494
rect 60620 42980 60676 42990
rect 60732 42980 60788 45054
rect 60956 44772 61012 47516
rect 60844 44716 61012 44772
rect 61068 47572 61124 47582
rect 60844 44324 60900 44716
rect 60956 44548 61012 44558
rect 61068 44548 61124 47516
rect 61292 47068 61348 47628
rect 61180 47012 61348 47068
rect 61180 45106 61236 47012
rect 61404 46676 61460 48076
rect 61516 48018 61572 48030
rect 61516 47966 61518 48018
rect 61570 47966 61572 48018
rect 61516 47684 61572 47966
rect 61516 47618 61572 47628
rect 61628 47234 61684 47246
rect 61628 47182 61630 47234
rect 61682 47182 61684 47234
rect 61628 47068 61684 47182
rect 61516 47012 61684 47068
rect 61516 46946 61572 46956
rect 61740 46900 61796 48524
rect 62076 48356 62132 48366
rect 62076 48262 62132 48300
rect 61852 48242 61908 48254
rect 61852 48190 61854 48242
rect 61906 48190 61908 48242
rect 61852 46900 61908 48190
rect 61964 48244 62020 48254
rect 61964 47682 62020 48188
rect 61964 47630 61966 47682
rect 62018 47630 62020 47682
rect 61964 47618 62020 47630
rect 62076 47908 62132 47918
rect 61964 47012 62020 47022
rect 61964 46900 62020 46956
rect 61852 46844 62020 46900
rect 61740 46834 61796 46844
rect 61404 46610 61460 46620
rect 61516 46674 61572 46686
rect 61964 46676 62020 46686
rect 61516 46622 61518 46674
rect 61570 46622 61572 46674
rect 61292 46564 61348 46574
rect 61292 46470 61348 46508
rect 61516 46340 61572 46622
rect 61852 46674 62020 46676
rect 61852 46622 61966 46674
rect 62018 46622 62020 46674
rect 61852 46620 62020 46622
rect 61516 46274 61572 46284
rect 61740 46562 61796 46574
rect 61740 46510 61742 46562
rect 61794 46510 61796 46562
rect 61740 46340 61796 46510
rect 61740 46274 61796 46284
rect 61292 45892 61348 45902
rect 61292 45798 61348 45836
rect 61628 45668 61684 45678
rect 61628 45574 61684 45612
rect 61628 45220 61684 45230
rect 61628 45126 61684 45164
rect 61180 45054 61182 45106
rect 61234 45054 61236 45106
rect 61180 45042 61236 45054
rect 61404 45108 61460 45118
rect 60956 44546 61348 44548
rect 60956 44494 60958 44546
rect 61010 44494 61348 44546
rect 60956 44492 61348 44494
rect 60956 44482 61012 44492
rect 60900 44268 61236 44324
rect 60844 44230 60900 44268
rect 61180 44210 61236 44268
rect 61180 44158 61182 44210
rect 61234 44158 61236 44210
rect 61180 44146 61236 44158
rect 60620 42978 60900 42980
rect 60620 42926 60622 42978
rect 60674 42926 60900 42978
rect 60620 42924 60900 42926
rect 60620 42914 60676 42924
rect 60396 42700 60788 42756
rect 60732 41298 60788 42700
rect 60732 41246 60734 41298
rect 60786 41246 60788 41298
rect 60732 41234 60788 41246
rect 60508 41188 60564 41198
rect 60508 41094 60564 41132
rect 60620 40516 60676 40526
rect 60508 40402 60564 40414
rect 60508 40350 60510 40402
rect 60562 40350 60564 40402
rect 60396 40292 60452 40302
rect 60396 38668 60452 40236
rect 60508 40180 60564 40350
rect 60508 39618 60564 40124
rect 60508 39566 60510 39618
rect 60562 39566 60564 39618
rect 60508 39554 60564 39566
rect 60620 39506 60676 40460
rect 60844 40068 60900 42924
rect 60956 42868 61012 42878
rect 60956 42754 61012 42812
rect 60956 42702 60958 42754
rect 61010 42702 61012 42754
rect 60956 41412 61012 42702
rect 61292 42756 61348 44492
rect 61292 42690 61348 42700
rect 61404 42754 61460 45052
rect 61516 44210 61572 44222
rect 61516 44158 61518 44210
rect 61570 44158 61572 44210
rect 61516 43652 61572 44158
rect 61516 42868 61572 43596
rect 61852 43204 61908 46620
rect 61964 46610 62020 46620
rect 62076 46004 62132 47852
rect 62188 47348 62244 47358
rect 62188 47254 62244 47292
rect 62188 46676 62244 46686
rect 62188 46674 62356 46676
rect 62188 46622 62190 46674
rect 62242 46622 62356 46674
rect 62188 46620 62356 46622
rect 62188 46610 62244 46620
rect 61964 45948 62132 46004
rect 61964 45890 62020 45948
rect 62188 45892 62244 45902
rect 61964 45838 61966 45890
rect 62018 45838 62020 45890
rect 61964 43540 62020 45838
rect 61964 43474 62020 43484
rect 62076 45836 62188 45892
rect 62076 44884 62132 45836
rect 62188 45798 62244 45836
rect 61964 43316 62020 43326
rect 61964 43222 62020 43260
rect 61516 42802 61572 42812
rect 61740 43148 61908 43204
rect 61404 42702 61406 42754
rect 61458 42702 61460 42754
rect 61404 42690 61460 42702
rect 61628 42756 61684 42766
rect 61628 42642 61684 42700
rect 61628 42590 61630 42642
rect 61682 42590 61684 42642
rect 61628 42578 61684 42590
rect 61292 42420 61348 42430
rect 61180 41972 61236 41982
rect 60956 41346 61012 41356
rect 61068 41860 61124 41870
rect 61068 41298 61124 41804
rect 61180 41524 61236 41916
rect 61180 41458 61236 41468
rect 61068 41246 61070 41298
rect 61122 41246 61124 41298
rect 61068 41234 61124 41246
rect 61180 41076 61236 41086
rect 61068 41074 61236 41076
rect 61068 41022 61182 41074
rect 61234 41022 61236 41074
rect 61068 41020 61236 41022
rect 60956 40964 61012 40974
rect 60956 40870 61012 40908
rect 61068 40852 61124 41020
rect 61180 41010 61236 41020
rect 61068 40404 61124 40796
rect 61068 40338 61124 40348
rect 61180 40628 61236 40638
rect 61180 40290 61236 40572
rect 61180 40238 61182 40290
rect 61234 40238 61236 40290
rect 61180 40226 61236 40238
rect 60844 40012 61236 40068
rect 60620 39454 60622 39506
rect 60674 39454 60676 39506
rect 60620 39442 60676 39454
rect 60956 39844 61012 39854
rect 60508 38948 60564 38958
rect 60508 38854 60564 38892
rect 60956 38948 61012 39788
rect 60732 38836 60788 38846
rect 60732 38742 60788 38780
rect 60172 32510 60174 32562
rect 60226 32510 60228 32562
rect 59724 32340 59780 32350
rect 58828 31780 58884 31790
rect 58828 31666 58884 31724
rect 58828 31614 58830 31666
rect 58882 31614 58884 31666
rect 58828 31602 58884 31614
rect 58716 31054 58718 31106
rect 58770 31054 58772 31106
rect 58716 31042 58772 31054
rect 59612 30996 59668 31006
rect 59612 30902 59668 30940
rect 59276 30882 59332 30894
rect 59276 30830 59278 30882
rect 59330 30830 59332 30882
rect 59276 30548 59332 30830
rect 59276 30482 59332 30492
rect 59724 30100 59780 32284
rect 60172 31780 60228 32510
rect 60172 31714 60228 31724
rect 60284 38612 60452 38668
rect 59948 31554 60004 31566
rect 59948 31502 59950 31554
rect 60002 31502 60004 31554
rect 59948 30548 60004 31502
rect 60284 30772 60340 38612
rect 60508 38052 60564 38062
rect 60508 37958 60564 37996
rect 60956 38052 61012 38892
rect 60956 37986 61012 37996
rect 61068 39730 61124 39742
rect 61068 39678 61070 39730
rect 61122 39678 61124 39730
rect 60844 37940 60900 37950
rect 60844 37846 60900 37884
rect 60620 37826 60676 37838
rect 60620 37774 60622 37826
rect 60674 37774 60676 37826
rect 60396 37492 60452 37502
rect 60396 37266 60452 37436
rect 60620 37380 60676 37774
rect 60620 37314 60676 37324
rect 60732 37826 60788 37838
rect 61068 37828 61124 39678
rect 60732 37774 60734 37826
rect 60786 37774 60788 37826
rect 60396 37214 60398 37266
rect 60450 37214 60452 37266
rect 60396 37202 60452 37214
rect 60732 37268 60788 37774
rect 60956 37772 61124 37828
rect 60732 37212 60900 37268
rect 60620 37044 60676 37054
rect 60620 36594 60676 36988
rect 60620 36542 60622 36594
rect 60674 36542 60676 36594
rect 60620 36530 60676 36542
rect 60508 36260 60564 36270
rect 60508 36166 60564 36204
rect 60732 36258 60788 36270
rect 60732 36206 60734 36258
rect 60786 36206 60788 36258
rect 60732 36036 60788 36206
rect 60844 36148 60900 37212
rect 60956 37044 61012 37772
rect 61068 37492 61124 37502
rect 61068 37266 61124 37436
rect 61068 37214 61070 37266
rect 61122 37214 61124 37266
rect 61068 37202 61124 37214
rect 60956 36988 61124 37044
rect 61068 36596 61124 36988
rect 61068 36530 61124 36540
rect 60956 36484 61012 36494
rect 60956 36372 61012 36428
rect 60956 36370 61124 36372
rect 60956 36318 60958 36370
rect 61010 36318 61124 36370
rect 60956 36316 61124 36318
rect 60956 36306 61012 36316
rect 60844 36082 60900 36092
rect 60732 35970 60788 35980
rect 61068 35138 61124 36316
rect 61068 35086 61070 35138
rect 61122 35086 61124 35138
rect 61068 35074 61124 35086
rect 60732 34916 60788 34926
rect 60732 34822 60788 34860
rect 60508 34802 60564 34814
rect 60508 34750 60510 34802
rect 60562 34750 60564 34802
rect 60508 33572 60564 34750
rect 60732 34244 60788 34254
rect 60732 34150 60788 34188
rect 60508 33506 60564 33516
rect 60732 33348 60788 33358
rect 60732 33254 60788 33292
rect 60508 33236 60564 33246
rect 60508 33142 60564 33180
rect 60508 32564 60564 32574
rect 60508 32470 60564 32508
rect 61068 32562 61124 32574
rect 61068 32510 61070 32562
rect 61122 32510 61124 32562
rect 61068 32002 61124 32510
rect 61180 32564 61236 40012
rect 61292 38668 61348 42364
rect 61628 41860 61684 41870
rect 61628 41766 61684 41804
rect 61740 41636 61796 43148
rect 62076 43092 62132 44828
rect 61404 41580 61796 41636
rect 61852 43036 62132 43092
rect 62188 44994 62244 45006
rect 62188 44942 62190 44994
rect 62242 44942 62244 44994
rect 61404 41076 61460 41580
rect 61404 40516 61460 41020
rect 61404 40402 61460 40460
rect 61628 41412 61684 41422
rect 61404 40350 61406 40402
rect 61458 40350 61460 40402
rect 61404 40338 61460 40350
rect 61516 40404 61572 40414
rect 61516 40180 61572 40348
rect 61404 40124 61572 40180
rect 61404 39284 61460 40124
rect 61404 39218 61460 39228
rect 61516 39618 61572 39630
rect 61516 39566 61518 39618
rect 61570 39566 61572 39618
rect 61404 38836 61460 38846
rect 61404 38742 61460 38780
rect 61292 38612 61460 38668
rect 61292 38052 61348 38062
rect 61292 37958 61348 37996
rect 61292 36484 61348 36494
rect 61292 36390 61348 36428
rect 61292 35252 61348 35262
rect 61292 34692 61348 35196
rect 61404 35140 61460 38612
rect 61516 37156 61572 39566
rect 61628 39396 61684 41356
rect 61740 41300 61796 41310
rect 61740 41186 61796 41244
rect 61740 41134 61742 41186
rect 61794 41134 61796 41186
rect 61740 41122 61796 41134
rect 61740 40962 61796 40974
rect 61740 40910 61742 40962
rect 61794 40910 61796 40962
rect 61740 40740 61796 40910
rect 61740 40674 61796 40684
rect 61740 40516 61796 40526
rect 61740 39508 61796 40460
rect 61852 39620 61908 43036
rect 62076 41972 62132 41982
rect 62076 41878 62132 41916
rect 62076 40404 62132 40414
rect 62076 40310 62132 40348
rect 62188 40292 62244 44942
rect 62300 41748 62356 46620
rect 62300 40628 62356 41692
rect 62300 40562 62356 40572
rect 62412 42196 62468 42206
rect 62188 40226 62244 40236
rect 61964 40180 62020 40190
rect 62020 40124 62132 40180
rect 61964 40114 62020 40124
rect 62076 39842 62132 40124
rect 62076 39790 62078 39842
rect 62130 39790 62132 39842
rect 62076 39778 62132 39790
rect 61852 39564 62132 39620
rect 61740 39452 62020 39508
rect 61628 39340 61796 39396
rect 61628 37826 61684 37838
rect 61628 37774 61630 37826
rect 61682 37774 61684 37826
rect 61628 37492 61684 37774
rect 61740 37492 61796 39340
rect 61852 38948 61908 38958
rect 61852 38722 61908 38892
rect 61852 38670 61854 38722
rect 61906 38670 61908 38722
rect 61852 38658 61908 38670
rect 61964 38050 62020 39452
rect 61964 37998 61966 38050
rect 62018 37998 62020 38050
rect 61964 37986 62020 37998
rect 62076 37828 62132 39564
rect 61964 37772 62132 37828
rect 62188 39506 62244 39518
rect 62188 39454 62190 39506
rect 62242 39454 62244 39506
rect 61852 37492 61908 37502
rect 61740 37490 61908 37492
rect 61740 37438 61854 37490
rect 61906 37438 61908 37490
rect 61740 37436 61908 37438
rect 61628 37426 61684 37436
rect 61852 37426 61908 37436
rect 61964 37268 62020 37772
rect 61852 37212 62020 37268
rect 62076 37268 62132 37278
rect 61516 37154 61684 37156
rect 61516 37102 61518 37154
rect 61570 37102 61684 37154
rect 61516 37100 61684 37102
rect 61516 37090 61572 37100
rect 61628 36482 61684 37100
rect 61628 36430 61630 36482
rect 61682 36430 61684 36482
rect 61516 36372 61572 36382
rect 61516 36278 61572 36316
rect 61628 36148 61684 36430
rect 61628 36082 61684 36092
rect 61740 36820 61796 36830
rect 61740 35586 61796 36764
rect 61740 35534 61742 35586
rect 61794 35534 61796 35586
rect 61740 35522 61796 35534
rect 61740 35140 61796 35150
rect 61404 35138 61796 35140
rect 61404 35086 61742 35138
rect 61794 35086 61796 35138
rect 61404 35084 61796 35086
rect 61740 35074 61796 35084
rect 61852 34804 61908 37212
rect 62076 37174 62132 37212
rect 62188 36932 62244 39454
rect 61964 36876 62244 36932
rect 61964 36820 62020 36876
rect 61964 36754 62020 36764
rect 61964 36596 62020 36606
rect 61964 36482 62020 36540
rect 61964 36430 61966 36482
rect 62018 36430 62020 36482
rect 61964 36418 62020 36430
rect 62188 35924 62244 35934
rect 62188 35830 62244 35868
rect 61964 34804 62020 34814
rect 61852 34802 62020 34804
rect 61852 34750 61966 34802
rect 62018 34750 62020 34802
rect 61852 34748 62020 34750
rect 61404 34692 61460 34702
rect 61292 34690 61460 34692
rect 61292 34638 61406 34690
rect 61458 34638 61460 34690
rect 61292 34636 61460 34638
rect 61404 34626 61460 34636
rect 61740 34244 61796 34254
rect 61740 34150 61796 34188
rect 61740 33348 61796 33358
rect 61740 33254 61796 33292
rect 61964 33234 62020 34748
rect 61964 33182 61966 33234
rect 62018 33182 62020 33234
rect 61404 33122 61460 33134
rect 61404 33070 61406 33122
rect 61458 33070 61460 33122
rect 61404 32676 61460 33070
rect 61628 32676 61684 32686
rect 61404 32674 61796 32676
rect 61404 32622 61630 32674
rect 61682 32622 61796 32674
rect 61404 32620 61796 32622
rect 61628 32610 61684 32620
rect 61236 32508 61460 32564
rect 61180 32498 61236 32508
rect 61068 31950 61070 32002
rect 61122 31950 61124 32002
rect 60508 31778 60564 31790
rect 60508 31726 60510 31778
rect 60562 31726 60564 31778
rect 60508 31332 60564 31726
rect 60508 31266 60564 31276
rect 60284 30706 60340 30716
rect 59948 30482 60004 30492
rect 59724 30034 59780 30044
rect 60284 30212 60340 30222
rect 58716 29986 58772 29998
rect 58716 29934 58718 29986
rect 58770 29934 58772 29986
rect 58716 28532 58772 29934
rect 59836 29986 59892 29998
rect 59836 29934 59838 29986
rect 59890 29934 59892 29986
rect 59612 29652 59668 29662
rect 58828 29540 58884 29550
rect 58828 29426 58884 29484
rect 58828 29374 58830 29426
rect 58882 29374 58884 29426
rect 58828 29362 58884 29374
rect 58716 28466 58772 28476
rect 58828 29204 58884 29214
rect 58604 27906 58660 27916
rect 58156 27858 58324 27860
rect 58156 27806 58158 27858
rect 58210 27806 58324 27858
rect 58156 27804 58324 27806
rect 58716 27860 58772 27870
rect 58828 27860 58884 29148
rect 59276 28532 59332 28542
rect 59276 28438 59332 28476
rect 58716 27858 58884 27860
rect 58716 27806 58718 27858
rect 58770 27806 58884 27858
rect 58716 27804 58884 27806
rect 58156 27794 58212 27804
rect 58716 27794 58772 27804
rect 58044 27582 58046 27634
rect 58098 27582 58100 27634
rect 58044 27570 58100 27582
rect 58268 27300 58324 27310
rect 58268 27206 58324 27244
rect 58044 27076 58100 27086
rect 57932 27074 58100 27076
rect 57932 27022 58046 27074
rect 58098 27022 58100 27074
rect 57932 27020 58100 27022
rect 58044 27010 58100 27020
rect 58828 27074 58884 27804
rect 59388 27634 59444 27646
rect 59388 27582 59390 27634
rect 59442 27582 59444 27634
rect 59388 27298 59444 27582
rect 59388 27246 59390 27298
rect 59442 27246 59444 27298
rect 58828 27022 58830 27074
rect 58882 27022 58884 27074
rect 58828 27010 58884 27022
rect 59052 27188 59108 27198
rect 57708 26462 57710 26514
rect 57762 26462 57764 26514
rect 57708 26450 57764 26462
rect 58268 26852 58324 26862
rect 58044 26068 58100 26078
rect 57708 25956 57764 25966
rect 57708 22148 57764 25900
rect 57820 24836 57876 24846
rect 57820 24742 57876 24780
rect 57820 23042 57876 23054
rect 57820 22990 57822 23042
rect 57874 22990 57876 23042
rect 57820 22260 57876 22990
rect 57820 22194 57876 22204
rect 57708 22082 57764 22092
rect 57596 21756 57876 21812
rect 57260 21534 57262 21586
rect 57314 21534 57316 21586
rect 57260 21364 57316 21534
rect 57260 21298 57316 21308
rect 57372 21700 57428 21710
rect 57372 19796 57428 21644
rect 57708 21588 57764 21598
rect 57596 21476 57652 21486
rect 57484 21474 57652 21476
rect 57484 21422 57598 21474
rect 57650 21422 57652 21474
rect 57484 21420 57652 21422
rect 57484 20020 57540 21420
rect 57596 21410 57652 21420
rect 57596 20244 57652 20282
rect 57596 20178 57652 20188
rect 57708 20130 57764 21532
rect 57708 20078 57710 20130
rect 57762 20078 57764 20130
rect 57708 20066 57764 20078
rect 57484 19964 57652 20020
rect 57596 19908 57652 19964
rect 57484 19796 57540 19806
rect 57372 19794 57540 19796
rect 57372 19742 57486 19794
rect 57538 19742 57540 19794
rect 57372 19740 57540 19742
rect 57484 19730 57540 19740
rect 57596 18676 57652 19852
rect 57708 18676 57764 18686
rect 57596 18674 57764 18676
rect 57596 18622 57710 18674
rect 57762 18622 57764 18674
rect 57596 18620 57764 18622
rect 57708 18610 57764 18620
rect 57148 18386 57204 18396
rect 57372 18450 57428 18462
rect 57372 18398 57374 18450
rect 57426 18398 57428 18450
rect 57036 17938 57092 17948
rect 57148 18228 57204 18238
rect 57036 17668 57092 17678
rect 57036 17574 57092 17612
rect 56588 17054 56590 17106
rect 56642 17054 56644 17106
rect 56588 17042 56644 17054
rect 56700 17500 56980 17556
rect 56588 16212 56644 16222
rect 56588 16098 56644 16156
rect 56588 16046 56590 16098
rect 56642 16046 56644 16098
rect 56588 16034 56644 16046
rect 56588 15316 56644 15326
rect 56476 15314 56644 15316
rect 56476 15262 56590 15314
rect 56642 15262 56644 15314
rect 56476 15260 56644 15262
rect 56252 11618 56308 11630
rect 56252 11566 56254 11618
rect 56306 11566 56308 11618
rect 56252 11506 56308 11566
rect 56252 11454 56254 11506
rect 56306 11454 56308 11506
rect 56252 11442 56308 11454
rect 56476 11284 56532 15260
rect 56588 15250 56644 15260
rect 56588 14196 56644 14206
rect 56588 13746 56644 14140
rect 56588 13694 56590 13746
rect 56642 13694 56644 13746
rect 56588 13682 56644 13694
rect 56588 13524 56644 13534
rect 56588 12962 56644 13468
rect 56588 12910 56590 12962
rect 56642 12910 56644 12962
rect 56588 12898 56644 12910
rect 56700 13412 56756 17500
rect 57148 16882 57204 18172
rect 57372 17780 57428 18398
rect 57372 17714 57428 17724
rect 57708 17444 57764 17454
rect 57596 16996 57652 17006
rect 57596 16902 57652 16940
rect 57708 16994 57764 17388
rect 57708 16942 57710 16994
rect 57762 16942 57764 16994
rect 57708 16930 57764 16942
rect 57372 16884 57428 16894
rect 57148 16830 57150 16882
rect 57202 16830 57204 16882
rect 57148 16818 57204 16830
rect 57260 16882 57428 16884
rect 57260 16830 57374 16882
rect 57426 16830 57428 16882
rect 57260 16828 57428 16830
rect 57036 15876 57092 15886
rect 56812 15204 56868 15214
rect 56812 13746 56868 15148
rect 56812 13694 56814 13746
rect 56866 13694 56868 13746
rect 56812 13682 56868 13694
rect 56588 12404 56644 12414
rect 56588 12310 56644 12348
rect 56700 11618 56756 13356
rect 56924 13188 56980 13198
rect 56924 13074 56980 13132
rect 56924 13022 56926 13074
rect 56978 13022 56980 13074
rect 56924 13010 56980 13022
rect 56924 12292 56980 12302
rect 57036 12292 57092 15820
rect 57260 14532 57316 16828
rect 57372 16818 57428 16828
rect 57820 16548 57876 21756
rect 57932 21588 57988 21598
rect 57932 21252 57988 21532
rect 57932 21186 57988 21196
rect 58044 21028 58100 26012
rect 58268 24834 58324 26796
rect 58604 26404 58660 26414
rect 58268 24782 58270 24834
rect 58322 24782 58324 24834
rect 58268 24770 58324 24782
rect 58492 25844 58548 25854
rect 58156 24724 58212 24734
rect 58156 24276 58212 24668
rect 58492 24722 58548 25788
rect 58604 25730 58660 26348
rect 59052 26290 59108 27132
rect 59388 26908 59444 27246
rect 59052 26238 59054 26290
rect 59106 26238 59108 26290
rect 59052 26226 59108 26238
rect 59164 26852 59444 26908
rect 59164 25732 59220 26852
rect 58604 25678 58606 25730
rect 58658 25678 58660 25730
rect 58604 25666 58660 25678
rect 58828 25676 59220 25732
rect 58716 25618 58772 25630
rect 58716 25566 58718 25618
rect 58770 25566 58772 25618
rect 58492 24670 58494 24722
rect 58546 24670 58548 24722
rect 58492 24658 58548 24670
rect 58604 25506 58660 25518
rect 58604 25454 58606 25506
rect 58658 25454 58660 25506
rect 58604 24948 58660 25454
rect 58156 24220 58324 24276
rect 58156 24052 58212 24062
rect 58156 23826 58212 23996
rect 58156 23774 58158 23826
rect 58210 23774 58212 23826
rect 58156 23762 58212 23774
rect 58156 22372 58212 22382
rect 58156 22278 58212 22316
rect 58268 21812 58324 24220
rect 58604 23156 58660 24892
rect 58716 23492 58772 25566
rect 58828 24946 58884 25676
rect 58828 24894 58830 24946
rect 58882 24894 58884 24946
rect 58828 24882 58884 24894
rect 59276 25172 59332 25182
rect 59276 24722 59332 25116
rect 59276 24670 59278 24722
rect 59330 24670 59332 24722
rect 59276 24658 59332 24670
rect 58716 23156 58772 23436
rect 59500 24500 59556 24510
rect 59052 23156 59108 23166
rect 58716 23154 59108 23156
rect 58716 23102 59054 23154
rect 59106 23102 59108 23154
rect 58716 23100 59108 23102
rect 58604 23062 58660 23100
rect 58828 22820 58884 22830
rect 58884 22764 58996 22820
rect 58828 22754 58884 22764
rect 57932 20972 58100 21028
rect 58156 21756 58324 21812
rect 57932 19012 57988 20972
rect 58156 20244 58212 21756
rect 58380 21700 58436 21710
rect 58380 21698 58548 21700
rect 58380 21646 58382 21698
rect 58434 21646 58548 21698
rect 58380 21644 58548 21646
rect 58380 21634 58436 21644
rect 58044 20188 58212 20244
rect 58268 21586 58324 21598
rect 58268 21534 58270 21586
rect 58322 21534 58324 21586
rect 58044 19572 58100 20188
rect 58156 20018 58212 20030
rect 58156 19966 58158 20018
rect 58210 19966 58212 20018
rect 58156 19796 58212 19966
rect 58156 19730 58212 19740
rect 58268 20020 58324 21534
rect 58380 21474 58436 21486
rect 58380 21422 58382 21474
rect 58434 21422 58436 21474
rect 58380 21028 58436 21422
rect 58380 20962 58436 20972
rect 58380 20804 58436 20814
rect 58380 20710 58436 20748
rect 58044 19506 58100 19516
rect 58156 19236 58212 19246
rect 58268 19236 58324 19964
rect 58212 19180 58324 19236
rect 58492 19234 58548 21644
rect 58828 21140 58884 21150
rect 58604 21028 58660 21038
rect 58604 20934 58660 20972
rect 58828 20802 58884 21084
rect 58828 20750 58830 20802
rect 58882 20750 58884 20802
rect 58828 20738 58884 20750
rect 58940 20356 58996 22764
rect 59052 22596 59108 23100
rect 59052 22530 59108 22540
rect 59388 22258 59444 22270
rect 59388 22206 59390 22258
rect 59442 22206 59444 22258
rect 59388 22148 59444 22206
rect 59388 22082 59444 22092
rect 59500 21812 59556 24444
rect 59612 23604 59668 29596
rect 59724 28980 59780 28990
rect 59724 28084 59780 28924
rect 59836 28644 59892 29934
rect 60284 29428 60340 30156
rect 61068 30212 61124 31950
rect 61068 30146 61124 30156
rect 61292 32338 61348 32350
rect 61292 32286 61294 32338
rect 61346 32286 61348 32338
rect 60508 29988 60564 29998
rect 60508 29894 60564 29932
rect 60620 29986 60676 29998
rect 60620 29934 60622 29986
rect 60674 29934 60676 29986
rect 59836 28578 59892 28588
rect 60060 28868 60116 28878
rect 59724 28028 60004 28084
rect 59724 27860 59780 27870
rect 59724 27766 59780 27804
rect 59724 27524 59780 27534
rect 59724 26516 59780 27468
rect 59836 27188 59892 27198
rect 59836 26962 59892 27132
rect 59836 26910 59838 26962
rect 59890 26910 59892 26962
rect 59836 26898 59892 26910
rect 59724 26460 59892 26516
rect 59724 26290 59780 26302
rect 59724 26238 59726 26290
rect 59778 26238 59780 26290
rect 59724 25844 59780 26238
rect 59724 25778 59780 25788
rect 59612 23548 59780 23604
rect 59164 21756 59556 21812
rect 59052 21588 59108 21626
rect 59052 21522 59108 21532
rect 59052 21362 59108 21374
rect 59052 21310 59054 21362
rect 59106 21310 59108 21362
rect 59052 21028 59108 21310
rect 59052 20962 59108 20972
rect 59052 20804 59108 20842
rect 59052 20738 59108 20748
rect 59164 20802 59220 21756
rect 59500 21700 59556 21756
rect 59612 21700 59668 21710
rect 59500 21698 59668 21700
rect 59500 21646 59614 21698
rect 59666 21646 59668 21698
rect 59500 21644 59668 21646
rect 59612 21634 59668 21644
rect 59276 21586 59332 21598
rect 59276 21534 59278 21586
rect 59330 21534 59332 21586
rect 59276 21364 59332 21534
rect 59500 21476 59556 21486
rect 59500 21382 59556 21420
rect 59332 21308 59444 21364
rect 59276 21298 59332 21308
rect 59164 20750 59166 20802
rect 59218 20750 59220 20802
rect 59164 20738 59220 20750
rect 59388 20692 59444 21308
rect 59500 20692 59556 20702
rect 59388 20690 59556 20692
rect 59388 20638 59502 20690
rect 59554 20638 59556 20690
rect 59388 20636 59556 20638
rect 59500 20626 59556 20636
rect 58828 20300 58996 20356
rect 59052 20580 59108 20590
rect 58492 19182 58494 19234
rect 58546 19182 58548 19234
rect 58156 19142 58212 19180
rect 57932 18956 58212 19012
rect 58044 18788 58100 18798
rect 57820 16482 57876 16492
rect 57932 18450 57988 18462
rect 57932 18398 57934 18450
rect 57986 18398 57988 18450
rect 57932 17442 57988 18398
rect 57932 17390 57934 17442
rect 57986 17390 57988 17442
rect 57596 16098 57652 16110
rect 57596 16046 57598 16098
rect 57650 16046 57652 16098
rect 57596 15988 57652 16046
rect 57596 15922 57652 15932
rect 57932 15988 57988 17390
rect 58044 16210 58100 18732
rect 58156 18340 58212 18956
rect 58492 18788 58548 19182
rect 58716 19796 58772 19806
rect 58492 18722 58548 18732
rect 58604 19122 58660 19134
rect 58604 19070 58606 19122
rect 58658 19070 58660 19122
rect 58156 18284 58324 18340
rect 58044 16158 58046 16210
rect 58098 16158 58100 16210
rect 58044 16146 58100 16158
rect 58156 16658 58212 16670
rect 58156 16606 58158 16658
rect 58210 16606 58212 16658
rect 58156 16100 58212 16606
rect 58156 16034 58212 16044
rect 57932 15922 57988 15932
rect 58044 15876 58100 15886
rect 57372 15202 57428 15214
rect 57372 15150 57374 15202
rect 57426 15150 57428 15202
rect 57372 15148 57428 15150
rect 57372 15092 57652 15148
rect 57596 14642 57652 15092
rect 57596 14590 57598 14642
rect 57650 14590 57652 14642
rect 57596 14578 57652 14590
rect 57484 14532 57540 14542
rect 57260 14530 57540 14532
rect 57260 14478 57486 14530
rect 57538 14478 57540 14530
rect 57260 14476 57540 14478
rect 57484 14466 57540 14476
rect 57708 14420 57764 14430
rect 57148 13748 57204 13758
rect 57148 13654 57204 13692
rect 57596 13636 57652 13646
rect 57372 13580 57596 13636
rect 57372 13074 57428 13580
rect 57596 13542 57652 13580
rect 57372 13022 57374 13074
rect 57426 13022 57428 13074
rect 57372 13010 57428 13022
rect 57596 13076 57652 13086
rect 56924 12290 57092 12292
rect 56924 12238 56926 12290
rect 56978 12238 57092 12290
rect 56924 12236 57092 12238
rect 57148 12628 57204 12638
rect 56924 12226 56980 12236
rect 56700 11566 56702 11618
rect 56754 11566 56756 11618
rect 56700 11506 56756 11566
rect 56700 11454 56702 11506
rect 56754 11454 56756 11506
rect 56700 11442 56756 11454
rect 57148 12180 57204 12572
rect 57148 11506 57204 12124
rect 57372 12068 57428 12078
rect 57372 11974 57428 12012
rect 57148 11454 57150 11506
rect 57202 11454 57204 11506
rect 57148 11442 57204 11454
rect 57596 11506 57652 13020
rect 57596 11454 57598 11506
rect 57650 11454 57652 11506
rect 57596 11442 57652 11454
rect 56140 11228 56420 11284
rect 56476 11228 56756 11284
rect 55580 9886 55582 9938
rect 55634 9886 55636 9938
rect 55580 9874 55636 9886
rect 56364 9938 56420 11228
rect 56364 9886 56366 9938
rect 56418 9886 56420 9938
rect 55020 9602 55076 9614
rect 55020 9550 55022 9602
rect 55074 9550 55076 9602
rect 54572 9268 54628 9278
rect 54516 9266 54628 9268
rect 54516 9214 54574 9266
rect 54626 9214 54628 9266
rect 54516 9212 54628 9214
rect 54460 9174 54516 9212
rect 54572 8596 54628 9212
rect 55020 8708 55076 9550
rect 55020 8642 55076 8652
rect 55916 9602 55972 9614
rect 55916 9550 55918 9602
rect 55970 9550 55972 9602
rect 54572 8530 54628 8540
rect 55916 8596 55972 9550
rect 55916 8530 55972 8540
rect 54012 7634 54068 7644
rect 54124 8036 54180 8046
rect 54124 7476 54180 7980
rect 54124 7410 54180 7420
rect 52444 7364 52500 7374
rect 52444 7270 52500 7308
rect 52892 7362 52948 7374
rect 52892 7310 52894 7362
rect 52946 7310 52948 7362
rect 52892 7028 52948 7310
rect 52892 6962 52948 6972
rect 52108 6466 52164 6478
rect 52108 6414 52110 6466
rect 52162 6414 52164 6466
rect 52108 6132 52164 6414
rect 52108 6066 52164 6076
rect 56364 4564 56420 9886
rect 56700 10834 56756 11228
rect 57708 11060 57764 14364
rect 57932 14306 57988 14318
rect 57932 14254 57934 14306
rect 57986 14254 57988 14306
rect 57932 13524 57988 14254
rect 57932 13458 57988 13468
rect 58044 13970 58100 15820
rect 58044 13918 58046 13970
rect 58098 13918 58100 13970
rect 57820 13412 57876 13422
rect 57820 13074 57876 13356
rect 58044 13300 58100 13918
rect 58044 13234 58100 13244
rect 58156 14756 58212 14766
rect 58156 13748 58212 14700
rect 57820 13022 57822 13074
rect 57874 13022 57876 13074
rect 57820 13010 57876 13022
rect 58156 12852 58212 13692
rect 58268 13076 58324 18284
rect 58492 18228 58548 18238
rect 58492 18134 58548 18172
rect 58380 16772 58436 16782
rect 58380 16210 58436 16716
rect 58604 16324 58660 19070
rect 58604 16258 58660 16268
rect 58380 16158 58382 16210
rect 58434 16158 58436 16210
rect 58380 16146 58436 16158
rect 58716 16100 58772 19740
rect 58828 18340 58884 20300
rect 58940 20132 58996 20142
rect 59052 20132 59108 20524
rect 59724 20356 59780 23548
rect 59836 21140 59892 26460
rect 59948 23380 60004 28028
rect 60060 24834 60116 28812
rect 60284 28532 60340 29372
rect 60396 29540 60452 29550
rect 60396 28868 60452 29484
rect 60620 28868 60676 29934
rect 60732 29986 60788 29998
rect 60732 29934 60734 29986
rect 60786 29934 60788 29986
rect 60732 29428 60788 29934
rect 60956 29988 61012 29998
rect 60956 29894 61012 29932
rect 61292 29540 61348 32286
rect 61404 31778 61460 32508
rect 61404 31726 61406 31778
rect 61458 31726 61460 31778
rect 61404 31714 61460 31726
rect 61628 31780 61684 31790
rect 61516 31556 61572 31566
rect 61516 31462 61572 31500
rect 61628 30324 61684 31724
rect 61740 31668 61796 32620
rect 61852 31668 61908 31678
rect 61740 31666 61908 31668
rect 61740 31614 61854 31666
rect 61906 31614 61908 31666
rect 61740 31612 61908 31614
rect 61852 31602 61908 31612
rect 61964 31444 62020 33182
rect 62076 34130 62132 34142
rect 62076 34078 62078 34130
rect 62130 34078 62132 34130
rect 62076 32452 62132 34078
rect 62412 33348 62468 42140
rect 62524 40852 62580 51212
rect 62636 46452 62692 52220
rect 62636 46386 62692 46396
rect 62636 45220 62692 45230
rect 62748 45220 62804 55244
rect 62972 52164 63028 52174
rect 62692 45164 62804 45220
rect 62860 46564 62916 46574
rect 62636 45154 62692 45164
rect 62524 40786 62580 40796
rect 62860 34244 62916 46508
rect 62860 34178 62916 34188
rect 62972 34692 63028 52108
rect 62412 33282 62468 33292
rect 62076 32386 62132 32396
rect 61628 30258 61684 30268
rect 61740 31388 62020 31444
rect 62076 31668 62132 31678
rect 61516 30210 61572 30222
rect 61516 30158 61518 30210
rect 61570 30158 61572 30210
rect 61404 30100 61460 30110
rect 61516 30100 61572 30158
rect 61460 30044 61572 30100
rect 61404 30034 61460 30044
rect 60732 29362 60788 29372
rect 61068 29538 61348 29540
rect 61068 29486 61294 29538
rect 61346 29486 61348 29538
rect 61068 29484 61348 29486
rect 61068 29204 61124 29484
rect 61292 29474 61348 29484
rect 61404 29426 61460 29438
rect 61404 29374 61406 29426
rect 61458 29374 61460 29426
rect 60844 29148 61124 29204
rect 61180 29316 61236 29326
rect 60396 28812 60564 28868
rect 60508 28642 60564 28812
rect 60620 28802 60676 28812
rect 60732 29092 60788 29102
rect 60732 28754 60788 29036
rect 60732 28702 60734 28754
rect 60786 28702 60788 28754
rect 60732 28690 60788 28702
rect 60508 28590 60510 28642
rect 60562 28590 60564 28642
rect 60508 28578 60564 28590
rect 60284 28476 60452 28532
rect 60396 28420 60452 28476
rect 60844 28530 60900 29148
rect 60844 28478 60846 28530
rect 60898 28478 60900 28530
rect 60844 28466 60900 28478
rect 61068 28644 61124 28654
rect 60732 28420 60788 28430
rect 60396 28418 60788 28420
rect 60396 28366 60734 28418
rect 60786 28366 60788 28418
rect 60396 28364 60788 28366
rect 60732 28354 60788 28364
rect 60284 28308 60340 28318
rect 60172 27634 60228 27646
rect 60172 27582 60174 27634
rect 60226 27582 60228 27634
rect 60172 27076 60228 27582
rect 60284 27524 60340 28252
rect 61068 27748 61124 28588
rect 60284 27458 60340 27468
rect 60844 27692 61124 27748
rect 61180 28642 61236 29260
rect 61180 28590 61182 28642
rect 61234 28590 61236 28642
rect 60620 27188 60676 27198
rect 60620 27094 60676 27132
rect 60844 27186 60900 27692
rect 60844 27134 60846 27186
rect 60898 27134 60900 27186
rect 60844 27122 60900 27134
rect 61180 27188 61236 28590
rect 61404 28420 61460 29374
rect 61628 28644 61684 28654
rect 61628 28550 61684 28588
rect 61292 27972 61348 27982
rect 61404 27972 61460 28364
rect 61348 27916 61460 27972
rect 61516 28532 61572 28542
rect 61516 28082 61572 28476
rect 61516 28030 61518 28082
rect 61570 28030 61572 28082
rect 61292 27906 61348 27916
rect 61180 27122 61236 27132
rect 61516 27188 61572 28030
rect 61516 27122 61572 27132
rect 60172 27010 60228 27020
rect 61404 27076 61460 27086
rect 61404 26982 61460 27020
rect 61740 26908 61796 31388
rect 61964 30884 62020 30894
rect 61964 30790 62020 30828
rect 62076 30660 62132 31612
rect 61852 30604 62132 30660
rect 61852 30098 61908 30604
rect 62636 30324 62692 30334
rect 61852 30046 61854 30098
rect 61906 30046 61908 30098
rect 61852 30034 61908 30046
rect 62188 30100 62244 30110
rect 62188 30006 62244 30044
rect 62412 29428 62468 29438
rect 61964 29202 62020 29214
rect 61964 29150 61966 29202
rect 62018 29150 62020 29202
rect 61964 28196 62020 29150
rect 62188 28642 62244 28654
rect 62188 28590 62190 28642
rect 62242 28590 62244 28642
rect 62188 28420 62244 28590
rect 62188 28354 62244 28364
rect 60172 26852 60228 26862
rect 60172 26290 60228 26796
rect 61180 26852 61236 26862
rect 61740 26852 61908 26908
rect 61180 26758 61236 26796
rect 61740 26628 61796 26638
rect 61628 26516 61684 26526
rect 61628 26422 61684 26460
rect 61740 26514 61796 26572
rect 61740 26462 61742 26514
rect 61794 26462 61796 26514
rect 61740 26450 61796 26462
rect 60172 26238 60174 26290
rect 60226 26238 60228 26290
rect 60172 26226 60228 26238
rect 60396 26404 60452 26414
rect 60396 26066 60452 26348
rect 60396 26014 60398 26066
rect 60450 26014 60452 26066
rect 60396 26002 60452 26014
rect 60956 25620 61012 25630
rect 60956 25618 61460 25620
rect 60956 25566 60958 25618
rect 61010 25566 61460 25618
rect 60956 25564 61460 25566
rect 60956 25554 61012 25564
rect 60620 25396 60676 25406
rect 60620 25302 60676 25340
rect 61292 25394 61348 25406
rect 61292 25342 61294 25394
rect 61346 25342 61348 25394
rect 60060 24782 60062 24834
rect 60114 24782 60116 24834
rect 60060 24770 60116 24782
rect 60956 24500 61012 24510
rect 61012 24444 61124 24500
rect 60956 24434 61012 24444
rect 60060 24164 60116 24174
rect 60956 24164 61012 24174
rect 60060 24070 60116 24108
rect 60844 24108 60956 24164
rect 60620 23828 60676 23838
rect 60620 23734 60676 23772
rect 59948 23324 60116 23380
rect 59836 21074 59892 21084
rect 59948 23154 60004 23166
rect 59948 23102 59950 23154
rect 60002 23102 60004 23154
rect 59948 21028 60004 23102
rect 59948 20962 60004 20972
rect 59836 20916 59892 20926
rect 59836 20802 59892 20860
rect 59836 20750 59838 20802
rect 59890 20750 59892 20802
rect 59836 20738 59892 20750
rect 59836 20356 59892 20366
rect 59724 20300 59836 20356
rect 59836 20290 59892 20300
rect 58940 20130 59108 20132
rect 58940 20078 58942 20130
rect 58994 20078 59108 20130
rect 58940 20076 59108 20078
rect 58940 20066 58996 20076
rect 58828 18274 58884 18284
rect 59052 19684 59108 19694
rect 58940 17556 58996 17566
rect 58604 16044 58772 16100
rect 58828 16100 58884 16110
rect 58604 14980 58660 16044
rect 58828 15148 58884 16044
rect 58268 13010 58324 13020
rect 58380 14924 58604 14980
rect 58268 12852 58324 12862
rect 57932 12850 58324 12852
rect 57932 12798 58270 12850
rect 58322 12798 58324 12850
rect 57932 12796 58324 12798
rect 57932 12402 57988 12796
rect 58268 12786 58324 12796
rect 58380 12628 58436 14924
rect 58604 14914 58660 14924
rect 58716 15092 58884 15148
rect 58604 14644 58660 14654
rect 58604 14306 58660 14588
rect 58716 14642 58772 15092
rect 58940 14980 58996 17500
rect 59052 15540 59108 19628
rect 59836 19460 59892 19470
rect 59836 19366 59892 19404
rect 59500 19234 59556 19246
rect 59500 19182 59502 19234
rect 59554 19182 59556 19234
rect 59388 18564 59444 18574
rect 59388 17554 59444 18508
rect 59500 17892 59556 19182
rect 59500 17826 59556 17836
rect 59724 19122 59780 19134
rect 59724 19070 59726 19122
rect 59778 19070 59780 19122
rect 59388 17502 59390 17554
rect 59442 17502 59444 17554
rect 59388 16994 59444 17502
rect 59388 16942 59390 16994
rect 59442 16942 59444 16994
rect 59276 16212 59332 16222
rect 59276 16118 59332 16156
rect 59052 15474 59108 15484
rect 59388 15204 59444 16942
rect 59500 16098 59556 16110
rect 59500 16046 59502 16098
rect 59554 16046 59556 16098
rect 59500 15988 59556 16046
rect 59500 15922 59556 15932
rect 59500 15204 59556 15214
rect 59388 15202 59556 15204
rect 59388 15150 59502 15202
rect 59554 15150 59556 15202
rect 59388 15148 59556 15150
rect 59500 15138 59556 15148
rect 58716 14590 58718 14642
rect 58770 14590 58772 14642
rect 58716 14578 58772 14590
rect 58828 14924 58996 14980
rect 59388 14980 59444 14990
rect 58604 14254 58606 14306
rect 58658 14254 58660 14306
rect 58604 14242 58660 14254
rect 58828 14532 58884 14924
rect 58492 14084 58548 14094
rect 58492 13970 58548 14028
rect 58492 13918 58494 13970
rect 58546 13918 58548 13970
rect 58492 13906 58548 13918
rect 58828 13074 58884 14476
rect 59276 14306 59332 14318
rect 59276 14254 59278 14306
rect 59330 14254 59332 14306
rect 58828 13022 58830 13074
rect 58882 13022 58884 13074
rect 58828 13010 58884 13022
rect 58940 13634 58996 13646
rect 58940 13582 58942 13634
rect 58994 13582 58996 13634
rect 57932 12350 57934 12402
rect 57986 12350 57988 12402
rect 57932 12338 57988 12350
rect 58044 12572 58436 12628
rect 58044 11506 58100 12572
rect 58828 12404 58884 12414
rect 58828 12310 58884 12348
rect 58268 12180 58324 12190
rect 58268 12086 58324 12124
rect 58940 12068 58996 13582
rect 59164 13076 59220 13086
rect 59164 12982 59220 13020
rect 59164 12068 59220 12078
rect 58940 12012 59164 12068
rect 59164 11974 59220 12012
rect 59276 11732 59332 14254
rect 59388 13970 59444 14924
rect 59724 14532 59780 19070
rect 59948 19124 60004 19134
rect 59836 19012 59892 19022
rect 59836 18918 59892 18956
rect 59948 18564 60004 19068
rect 59948 18470 60004 18508
rect 59836 18452 59892 18462
rect 59836 18340 59892 18396
rect 60060 18452 60116 23324
rect 60620 22596 60676 22606
rect 60844 22596 60900 24108
rect 60956 24098 61012 24108
rect 60956 23940 61012 23950
rect 61068 23940 61124 24444
rect 60956 23938 61124 23940
rect 60956 23886 60958 23938
rect 61010 23886 61124 23938
rect 60956 23884 61124 23886
rect 60956 23874 61012 23884
rect 61180 23826 61236 23838
rect 61180 23774 61182 23826
rect 61234 23774 61236 23826
rect 60956 23268 61012 23278
rect 60956 23174 61012 23212
rect 61180 23156 61236 23774
rect 60956 22596 61012 22606
rect 60844 22594 61012 22596
rect 60844 22542 60958 22594
rect 61010 22542 61012 22594
rect 60844 22540 61012 22542
rect 60620 22502 60676 22540
rect 60956 22530 61012 22540
rect 60508 21812 60564 21822
rect 60396 21588 60452 21598
rect 60172 21364 60228 21402
rect 60172 21298 60228 21308
rect 60060 18386 60116 18396
rect 60172 21140 60228 21150
rect 59836 18284 60004 18340
rect 59388 13918 59390 13970
rect 59442 13918 59444 13970
rect 59388 13906 59444 13918
rect 59500 14476 59780 14532
rect 59836 16548 59892 16558
rect 59500 12852 59556 14476
rect 59724 14308 59780 14318
rect 59836 14308 59892 16492
rect 59948 15538 60004 18284
rect 60172 17108 60228 21084
rect 60284 20132 60340 20142
rect 60284 19012 60340 20076
rect 60284 18946 60340 18956
rect 60396 17108 60452 21532
rect 60508 21026 60564 21756
rect 60508 20974 60510 21026
rect 60562 20974 60564 21026
rect 60508 20962 60564 20974
rect 60620 20916 60676 20926
rect 60508 20692 60564 20702
rect 60508 19458 60564 20636
rect 60508 19406 60510 19458
rect 60562 19406 60564 19458
rect 60508 19394 60564 19406
rect 60508 19236 60564 19246
rect 60620 19236 60676 20860
rect 60732 20804 60788 20814
rect 60732 20710 60788 20748
rect 60956 20804 61012 20814
rect 61180 20804 61236 23100
rect 61292 22258 61348 25342
rect 61292 22206 61294 22258
rect 61346 22206 61348 22258
rect 61292 21364 61348 22206
rect 61404 22260 61460 25564
rect 61516 25394 61572 25406
rect 61516 25342 61518 25394
rect 61570 25342 61572 25394
rect 61516 24164 61572 25342
rect 61516 24098 61572 24108
rect 61628 23826 61684 23838
rect 61628 23774 61630 23826
rect 61682 23774 61684 23826
rect 61516 22260 61572 22270
rect 61404 22258 61572 22260
rect 61404 22206 61518 22258
rect 61570 22206 61572 22258
rect 61404 22204 61572 22206
rect 61516 21812 61572 22204
rect 61292 21298 61348 21308
rect 61404 21810 61572 21812
rect 61404 21758 61518 21810
rect 61570 21758 61572 21810
rect 61404 21756 61572 21758
rect 61012 20748 61236 20804
rect 60956 20738 61012 20748
rect 60956 20578 61012 20590
rect 60956 20526 60958 20578
rect 61010 20526 61012 20578
rect 60956 20244 61012 20526
rect 61068 20580 61124 20590
rect 61068 20486 61124 20524
rect 61180 20578 61236 20590
rect 61180 20526 61182 20578
rect 61234 20526 61236 20578
rect 61180 20468 61236 20526
rect 61180 20402 61236 20412
rect 61404 20244 61460 21756
rect 61516 21746 61572 21756
rect 61628 21476 61684 23774
rect 60956 20188 61348 20244
rect 61068 19906 61124 19918
rect 61068 19854 61070 19906
rect 61122 19854 61124 19906
rect 60732 19236 60788 19246
rect 60620 19234 60788 19236
rect 60620 19182 60734 19234
rect 60786 19182 60788 19234
rect 60620 19180 60788 19182
rect 60508 18788 60564 19180
rect 60732 19170 60788 19180
rect 60564 18732 60676 18788
rect 60508 18722 60564 18732
rect 60620 18116 60676 18732
rect 60844 18676 60900 18686
rect 60844 18582 60900 18620
rect 61068 18452 61124 19854
rect 61292 18900 61348 20188
rect 61404 20178 61460 20188
rect 61516 21420 61684 21476
rect 61516 20130 61572 21420
rect 61628 21028 61684 21038
rect 61628 20934 61684 20972
rect 61516 20078 61518 20130
rect 61570 20078 61572 20130
rect 61516 20066 61572 20078
rect 61404 20020 61460 20030
rect 61404 19926 61460 19964
rect 61628 20018 61684 20030
rect 61628 19966 61630 20018
rect 61682 19966 61684 20018
rect 61628 19236 61684 19966
rect 61852 19796 61908 26852
rect 61964 26514 62020 28140
rect 62076 27636 62132 27646
rect 62076 27298 62132 27580
rect 62076 27246 62078 27298
rect 62130 27246 62132 27298
rect 62076 27234 62132 27246
rect 62188 27188 62244 27198
rect 62244 27132 62356 27188
rect 62188 27094 62244 27132
rect 61964 26462 61966 26514
rect 62018 26462 62020 26514
rect 61964 26450 62020 26462
rect 62188 26404 62244 26414
rect 62188 26310 62244 26348
rect 62188 24612 62244 24622
rect 62300 24612 62356 27132
rect 62188 24610 62356 24612
rect 62188 24558 62190 24610
rect 62242 24558 62356 24610
rect 62188 24556 62356 24558
rect 62188 24546 62244 24556
rect 62076 22930 62132 22942
rect 62076 22878 62078 22930
rect 62130 22878 62132 22930
rect 61964 21028 62020 21038
rect 62076 21028 62132 22878
rect 61964 21026 62132 21028
rect 61964 20974 61966 21026
rect 62018 20974 62132 21026
rect 61964 20972 62132 20974
rect 62188 22036 62244 22046
rect 61964 20916 62020 20972
rect 61964 20850 62020 20860
rect 62188 20914 62244 21980
rect 62188 20862 62190 20914
rect 62242 20862 62244 20914
rect 62188 20850 62244 20862
rect 62076 20356 62132 20366
rect 62132 20300 62244 20356
rect 62076 20290 62132 20300
rect 61964 20018 62020 20030
rect 61964 19966 61966 20018
rect 62018 19966 62020 20018
rect 61964 19908 62020 19966
rect 61964 19842 62020 19852
rect 61628 19170 61684 19180
rect 61740 19740 61908 19796
rect 61404 19124 61460 19134
rect 61404 19030 61460 19068
rect 61516 19010 61572 19022
rect 61516 18958 61518 19010
rect 61570 18958 61572 19010
rect 61404 18900 61460 18910
rect 61516 18900 61572 18958
rect 61292 18844 61404 18900
rect 61460 18844 61572 18900
rect 61628 19012 61684 19022
rect 61404 18834 61460 18844
rect 61628 18788 61684 18956
rect 61516 18732 61684 18788
rect 61180 18452 61236 18462
rect 61068 18450 61236 18452
rect 61068 18398 61182 18450
rect 61234 18398 61236 18450
rect 61068 18396 61236 18398
rect 60620 18060 61012 18116
rect 60620 17892 60676 17902
rect 60620 17798 60676 17836
rect 60508 17780 60564 17790
rect 60508 17666 60564 17724
rect 60508 17614 60510 17666
rect 60562 17614 60564 17666
rect 60508 17602 60564 17614
rect 60732 17780 60788 17790
rect 60732 17666 60788 17724
rect 60732 17614 60734 17666
rect 60786 17614 60788 17666
rect 60732 17602 60788 17614
rect 60844 17556 60900 17566
rect 60508 17108 60564 17118
rect 60396 17106 60564 17108
rect 60396 17054 60510 17106
rect 60562 17054 60564 17106
rect 60396 17052 60564 17054
rect 60172 17042 60228 17052
rect 60508 17042 60564 17052
rect 60844 17106 60900 17500
rect 60956 17554 61012 18060
rect 60956 17502 60958 17554
rect 61010 17502 61012 17554
rect 60956 17490 61012 17502
rect 60844 17054 60846 17106
rect 60898 17054 60900 17106
rect 60844 17042 60900 17054
rect 61180 17106 61236 18396
rect 61292 18340 61348 18350
rect 61292 17554 61348 18284
rect 61292 17502 61294 17554
rect 61346 17502 61348 17554
rect 61292 17490 61348 17502
rect 61180 17054 61182 17106
rect 61234 17054 61236 17106
rect 61180 17042 61236 17054
rect 61404 17444 61460 17454
rect 60620 16772 60676 16782
rect 60620 16210 60676 16716
rect 60620 16158 60622 16210
rect 60674 16158 60676 16210
rect 60620 16146 60676 16158
rect 61180 16436 61236 16446
rect 61068 15876 61124 15886
rect 61068 15782 61124 15820
rect 59948 15486 59950 15538
rect 60002 15486 60004 15538
rect 59948 15474 60004 15486
rect 60396 15540 60452 15550
rect 60396 15446 60452 15484
rect 60844 15540 60900 15550
rect 60844 15446 60900 15484
rect 61068 14756 61124 14766
rect 61068 14642 61124 14700
rect 61068 14590 61070 14642
rect 61122 14590 61124 14642
rect 60620 14532 60676 14542
rect 60620 14438 60676 14476
rect 61068 14420 61124 14590
rect 61068 14354 61124 14364
rect 59724 14306 59892 14308
rect 59724 14254 59726 14306
rect 59778 14254 59892 14306
rect 59724 14252 59892 14254
rect 59724 14242 59780 14252
rect 59612 13972 59668 13982
rect 59612 13074 59668 13916
rect 60284 13972 60340 13982
rect 60284 13878 60340 13916
rect 61180 13970 61236 16380
rect 61404 16324 61460 17388
rect 61516 17106 61572 18732
rect 61516 17054 61518 17106
rect 61570 17054 61572 17106
rect 61516 17042 61572 17054
rect 61628 17780 61684 17790
rect 61628 17666 61684 17724
rect 61628 17614 61630 17666
rect 61682 17614 61684 17666
rect 61292 16268 61460 16324
rect 61516 16548 61572 16558
rect 61292 14644 61348 16268
rect 61516 16210 61572 16492
rect 61516 16158 61518 16210
rect 61570 16158 61572 16210
rect 61516 16146 61572 16158
rect 61404 15540 61460 15550
rect 61404 15446 61460 15484
rect 61628 15148 61684 17614
rect 61740 15538 61796 19740
rect 61852 19572 61908 19582
rect 61852 19122 61908 19516
rect 61852 19070 61854 19122
rect 61906 19070 61908 19122
rect 61852 19058 61908 19070
rect 62188 19012 62244 20300
rect 62188 19010 62356 19012
rect 62188 18958 62190 19010
rect 62242 18958 62356 19010
rect 62188 18956 62356 18958
rect 62188 18946 62244 18956
rect 62188 18788 62244 18798
rect 61852 18562 61908 18574
rect 61852 18510 61854 18562
rect 61906 18510 61908 18562
rect 61852 18340 61908 18510
rect 62076 18452 62132 18462
rect 61852 18274 61908 18284
rect 61964 18396 62076 18452
rect 61852 17668 61908 17678
rect 61852 17574 61908 17612
rect 61964 17220 62020 18396
rect 62076 18358 62132 18396
rect 62188 17666 62244 18732
rect 62188 17614 62190 17666
rect 62242 17614 62244 17666
rect 62188 17602 62244 17614
rect 62076 17444 62132 17454
rect 62076 17350 62132 17388
rect 61964 17164 62132 17220
rect 61852 16994 61908 17006
rect 61852 16942 61854 16994
rect 61906 16942 61908 16994
rect 61852 16660 61908 16942
rect 61852 16594 61908 16604
rect 61964 16996 62020 17006
rect 61964 16436 62020 16940
rect 61740 15486 61742 15538
rect 61794 15486 61796 15538
rect 61740 15474 61796 15486
rect 61852 16380 62020 16436
rect 61628 15092 61796 15148
rect 61292 14578 61348 14588
rect 61628 14644 61684 14654
rect 61628 14550 61684 14588
rect 61180 13918 61182 13970
rect 61234 13918 61236 13970
rect 60732 13860 60788 13870
rect 60732 13766 60788 13804
rect 59836 13748 59892 13758
rect 59836 13654 59892 13692
rect 59612 13022 59614 13074
rect 59666 13022 59668 13074
rect 59612 13010 59668 13022
rect 59500 12404 59556 12796
rect 59612 12404 59668 12414
rect 59500 12402 59668 12404
rect 59500 12350 59614 12402
rect 59666 12350 59668 12402
rect 59500 12348 59668 12350
rect 59612 12338 59668 12348
rect 61180 12404 61236 13918
rect 61740 13970 61796 15092
rect 61740 13918 61742 13970
rect 61794 13918 61796 13970
rect 61740 13906 61796 13918
rect 61852 13074 61908 16380
rect 61964 16212 62020 16222
rect 61964 16118 62020 16156
rect 62076 14420 62132 17164
rect 62188 17108 62244 17118
rect 62188 17014 62244 17052
rect 62188 15540 62244 15550
rect 62188 14642 62244 15484
rect 62188 14590 62190 14642
rect 62242 14590 62244 14642
rect 62188 14578 62244 14590
rect 62076 14364 62244 14420
rect 62188 13970 62244 14364
rect 62188 13918 62190 13970
rect 62242 13918 62244 13970
rect 62188 13906 62244 13918
rect 61852 13022 61854 13074
rect 61906 13022 61908 13074
rect 61852 13010 61908 13022
rect 62300 13074 62356 18956
rect 62412 14756 62468 29372
rect 62524 25956 62580 25966
rect 62524 16772 62580 25900
rect 62524 16706 62580 16716
rect 62636 15540 62692 30268
rect 62972 30324 63028 34636
rect 62972 30258 63028 30268
rect 62860 29988 62916 29998
rect 62860 19460 62916 29932
rect 62860 19394 62916 19404
rect 62972 27636 63028 27646
rect 62972 17780 63028 27580
rect 62972 17714 63028 17724
rect 62636 15474 62692 15484
rect 62412 14690 62468 14700
rect 62300 13022 62302 13074
rect 62354 13022 62356 13074
rect 62300 13010 62356 13022
rect 61180 12338 61236 12348
rect 59276 11666 59332 11676
rect 58044 11454 58046 11506
rect 58098 11454 58100 11506
rect 58044 11442 58100 11454
rect 56700 10782 56702 10834
rect 56754 10782 56756 10834
rect 56700 8036 56756 10782
rect 57148 11004 57764 11060
rect 57148 10836 57204 11004
rect 57148 10742 57204 10780
rect 56700 7970 56756 7980
rect 56364 4498 56420 4508
rect 51772 3266 51828 3276
rect 46396 3154 46452 3164
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 38220 1708 38388 1764
rect 38332 800 38388 1708
rect 34636 700 35028 756
rect 38304 0 38416 800
<< via2 >>
rect 11452 60508 11508 60564
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 10108 57148 10164 57204
rect 5740 56924 5796 56980
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 1708 55020 1764 55076
rect 1708 54460 1764 54516
rect 1596 53900 1652 53956
rect 1484 53452 1540 53508
rect 1260 48188 1316 48244
rect 1148 45500 1204 45556
rect 1148 38892 1204 38948
rect 1148 30380 1204 30436
rect 924 23660 980 23716
rect 924 17724 980 17780
rect 2492 55074 2548 55076
rect 2492 55022 2494 55074
rect 2494 55022 2546 55074
rect 2546 55022 2548 55074
rect 2492 55020 2548 55022
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4844 51602 4900 51604
rect 4844 51550 4846 51602
rect 4846 51550 4898 51602
rect 4898 51550 4900 51602
rect 4844 51548 4900 51550
rect 2828 50540 2884 50596
rect 1484 46956 1540 47012
rect 1596 49532 1652 49588
rect 1484 39452 1540 39508
rect 1932 49196 1988 49252
rect 1708 48802 1764 48804
rect 1708 48750 1710 48802
rect 1710 48750 1762 48802
rect 1762 48750 1764 48802
rect 1708 48748 1764 48750
rect 2044 48914 2100 48916
rect 2044 48862 2046 48914
rect 2046 48862 2098 48914
rect 2098 48862 2100 48914
rect 2044 48860 2100 48862
rect 1932 48242 1988 48244
rect 1932 48190 1934 48242
rect 1934 48190 1986 48242
rect 1986 48190 1988 48242
rect 1932 48188 1988 48190
rect 1708 48076 1764 48132
rect 2716 49810 2772 49812
rect 2716 49758 2718 49810
rect 2718 49758 2770 49810
rect 2770 49758 2772 49810
rect 2716 49756 2772 49758
rect 2492 49196 2548 49252
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4172 50652 4228 50708
rect 4396 50482 4452 50484
rect 4396 50430 4398 50482
rect 4398 50430 4450 50482
rect 4450 50430 4452 50482
rect 4396 50428 4452 50430
rect 5180 50594 5236 50596
rect 5180 50542 5182 50594
rect 5182 50542 5234 50594
rect 5234 50542 5236 50594
rect 5180 50540 5236 50542
rect 3388 49756 3444 49812
rect 3948 49532 4004 49588
rect 3836 49084 3892 49140
rect 2716 48914 2772 48916
rect 2716 48862 2718 48914
rect 2718 48862 2770 48914
rect 2770 48862 2772 48914
rect 2716 48860 2772 48862
rect 2380 48188 2436 48244
rect 2492 46844 2548 46900
rect 2268 46786 2324 46788
rect 2268 46734 2270 46786
rect 2270 46734 2322 46786
rect 2322 46734 2324 46786
rect 2268 46732 2324 46734
rect 2380 45948 2436 46004
rect 1708 45052 1764 45108
rect 1820 44322 1876 44324
rect 1820 44270 1822 44322
rect 1822 44270 1874 44322
rect 1874 44270 1876 44322
rect 1820 44268 1876 44270
rect 2044 44210 2100 44212
rect 2044 44158 2046 44210
rect 2046 44158 2098 44210
rect 2098 44158 2100 44210
rect 2044 44156 2100 44158
rect 2716 46060 2772 46116
rect 2604 45724 2660 45780
rect 2716 45388 2772 45444
rect 2268 44268 2324 44324
rect 2604 44268 2660 44324
rect 2380 44210 2436 44212
rect 2380 44158 2382 44210
rect 2382 44158 2434 44210
rect 2434 44158 2436 44210
rect 2380 44156 2436 44158
rect 3500 48914 3556 48916
rect 3500 48862 3502 48914
rect 3502 48862 3554 48914
rect 3554 48862 3556 48914
rect 3500 48860 3556 48862
rect 3612 46844 3668 46900
rect 3164 45218 3220 45220
rect 3164 45166 3166 45218
rect 3166 45166 3218 45218
rect 3218 45166 3220 45218
rect 3164 45164 3220 45166
rect 3052 45106 3108 45108
rect 3052 45054 3054 45106
rect 3054 45054 3106 45106
rect 3106 45054 3108 45106
rect 3052 45052 3108 45054
rect 3052 44210 3108 44212
rect 3052 44158 3054 44210
rect 3054 44158 3106 44210
rect 3106 44158 3108 44210
rect 3052 44156 3108 44158
rect 2156 42924 2212 42980
rect 2156 42642 2212 42644
rect 2156 42590 2158 42642
rect 2158 42590 2210 42642
rect 2210 42590 2212 42642
rect 2156 42588 2212 42590
rect 2044 41916 2100 41972
rect 1596 39116 1652 39172
rect 2156 41858 2212 41860
rect 2156 41806 2158 41858
rect 2158 41806 2210 41858
rect 2210 41806 2212 41858
rect 2156 41804 2212 41806
rect 1596 38892 1652 38948
rect 1596 37884 1652 37940
rect 1484 36092 1540 36148
rect 3612 46060 3668 46116
rect 3612 45836 3668 45892
rect 3388 45052 3444 45108
rect 3948 48748 4004 48804
rect 4060 49026 4116 49028
rect 4060 48974 4062 49026
rect 4062 48974 4114 49026
rect 4114 48974 4116 49026
rect 4060 48972 4116 48974
rect 4172 48636 4228 48692
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4508 49138 4564 49140
rect 4508 49086 4510 49138
rect 4510 49086 4562 49138
rect 4562 49086 4564 49138
rect 4508 49084 4564 49086
rect 4732 49026 4788 49028
rect 4732 48974 4734 49026
rect 4734 48974 4786 49026
rect 4786 48974 4788 49026
rect 4732 48972 4788 48974
rect 3948 46956 4004 47012
rect 3836 46674 3892 46676
rect 3836 46622 3838 46674
rect 3838 46622 3890 46674
rect 3890 46622 3892 46674
rect 3836 46620 3892 46622
rect 4060 46620 4116 46676
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4732 47628 4788 47684
rect 5516 49532 5572 49588
rect 5628 49138 5684 49140
rect 5628 49086 5630 49138
rect 5630 49086 5682 49138
rect 5682 49086 5684 49138
rect 5628 49084 5684 49086
rect 4956 48860 5012 48916
rect 8652 55020 8708 55076
rect 9548 54796 9604 54852
rect 8652 53506 8708 53508
rect 8652 53454 8654 53506
rect 8654 53454 8706 53506
rect 8706 53454 8708 53506
rect 8652 53452 8708 53454
rect 9100 53506 9156 53508
rect 9100 53454 9102 53506
rect 9102 53454 9154 53506
rect 9154 53454 9156 53506
rect 9100 53452 9156 53454
rect 8540 53228 8596 53284
rect 6860 52892 6916 52948
rect 7756 52946 7812 52948
rect 7756 52894 7758 52946
rect 7758 52894 7810 52946
rect 7810 52894 7812 52946
rect 7756 52892 7812 52894
rect 6188 52108 6244 52164
rect 5852 51602 5908 51604
rect 5852 51550 5854 51602
rect 5854 51550 5906 51602
rect 5906 51550 5908 51602
rect 5852 51548 5908 51550
rect 6524 51660 6580 51716
rect 6412 51100 6468 51156
rect 5964 50034 6020 50036
rect 5964 49982 5966 50034
rect 5966 49982 6018 50034
rect 6018 49982 6020 50034
rect 5964 49980 6020 49982
rect 5852 49026 5908 49028
rect 5852 48974 5854 49026
rect 5854 48974 5906 49026
rect 5906 48974 5908 49026
rect 5852 48972 5908 48974
rect 6076 48636 6132 48692
rect 4956 47740 5012 47796
rect 4956 47346 5012 47348
rect 4956 47294 4958 47346
rect 4958 47294 5010 47346
rect 5010 47294 5012 47346
rect 4956 47292 5012 47294
rect 5404 47292 5460 47348
rect 5068 47234 5124 47236
rect 5068 47182 5070 47234
rect 5070 47182 5122 47234
rect 5122 47182 5124 47234
rect 5068 47180 5124 47182
rect 4508 46396 4564 46452
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4172 45836 4228 45892
rect 4284 45500 4340 45556
rect 4508 45388 4564 45444
rect 4060 45164 4116 45220
rect 3500 44434 3556 44436
rect 3500 44382 3502 44434
rect 3502 44382 3554 44434
rect 3554 44382 3556 44434
rect 3500 44380 3556 44382
rect 3388 44322 3444 44324
rect 3388 44270 3390 44322
rect 3390 44270 3442 44322
rect 3442 44270 3444 44322
rect 3388 44268 3444 44270
rect 3276 44044 3332 44100
rect 2492 42978 2548 42980
rect 2492 42926 2494 42978
rect 2494 42926 2546 42978
rect 2546 42926 2548 42978
rect 2492 42924 2548 42926
rect 1932 40962 1988 40964
rect 1932 40910 1934 40962
rect 1934 40910 1986 40962
rect 1986 40910 1988 40962
rect 1932 40908 1988 40910
rect 2268 40684 2324 40740
rect 2492 42588 2548 42644
rect 3836 43820 3892 43876
rect 4172 45052 4228 45108
rect 4620 45052 4676 45108
rect 4844 45666 4900 45668
rect 4844 45614 4846 45666
rect 4846 45614 4898 45666
rect 4898 45614 4900 45666
rect 4844 45612 4900 45614
rect 4844 44994 4900 44996
rect 4844 44942 4846 44994
rect 4846 44942 4898 44994
rect 4898 44942 4900 44994
rect 4844 44940 4900 44942
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4620 44434 4676 44436
rect 4620 44382 4622 44434
rect 4622 44382 4674 44434
rect 4674 44382 4676 44434
rect 4620 44380 4676 44382
rect 4396 44322 4452 44324
rect 4396 44270 4398 44322
rect 4398 44270 4450 44322
rect 4450 44270 4452 44322
rect 4396 44268 4452 44270
rect 4172 44210 4228 44212
rect 4172 44158 4174 44210
rect 4174 44158 4226 44210
rect 4226 44158 4228 44210
rect 4172 44156 4228 44158
rect 4060 44044 4116 44100
rect 3724 43260 3780 43316
rect 3388 42588 3444 42644
rect 3724 42924 3780 42980
rect 3164 42252 3220 42308
rect 3276 42476 3332 42532
rect 3388 42364 3444 42420
rect 2940 41970 2996 41972
rect 2940 41918 2942 41970
rect 2942 41918 2994 41970
rect 2994 41918 2996 41970
rect 2940 41916 2996 41918
rect 2716 40514 2772 40516
rect 2716 40462 2718 40514
rect 2718 40462 2770 40514
rect 2770 40462 2772 40514
rect 2716 40460 2772 40462
rect 2268 39452 2324 39508
rect 2380 40236 2436 40292
rect 2940 41468 2996 41524
rect 3164 41916 3220 41972
rect 2940 41298 2996 41300
rect 2940 41246 2942 41298
rect 2942 41246 2994 41298
rect 2994 41246 2996 41298
rect 2940 41244 2996 41246
rect 3164 40460 3220 40516
rect 3388 40290 3444 40292
rect 3388 40238 3390 40290
rect 3390 40238 3442 40290
rect 3442 40238 3444 40290
rect 3388 40236 3444 40238
rect 2044 38556 2100 38612
rect 2268 38220 2324 38276
rect 2492 37436 2548 37492
rect 2716 37938 2772 37940
rect 2716 37886 2718 37938
rect 2718 37886 2770 37938
rect 2770 37886 2772 37938
rect 2716 37884 2772 37886
rect 2716 37660 2772 37716
rect 2828 37378 2884 37380
rect 2828 37326 2830 37378
rect 2830 37326 2882 37378
rect 2882 37326 2884 37378
rect 2828 37324 2884 37326
rect 3052 38108 3108 38164
rect 4172 43372 4228 43428
rect 4508 43260 4564 43316
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4172 42978 4228 42980
rect 4172 42926 4174 42978
rect 4174 42926 4226 42978
rect 4226 42926 4228 42978
rect 4172 42924 4228 42926
rect 4620 42866 4676 42868
rect 4620 42814 4622 42866
rect 4622 42814 4674 42866
rect 4674 42814 4676 42866
rect 4620 42812 4676 42814
rect 4060 42642 4116 42644
rect 4060 42590 4062 42642
rect 4062 42590 4114 42642
rect 4114 42590 4116 42642
rect 4060 42588 4116 42590
rect 4844 42588 4900 42644
rect 3948 42082 4004 42084
rect 3948 42030 3950 42082
rect 3950 42030 4002 42082
rect 4002 42030 4004 42082
rect 3948 42028 4004 42030
rect 3948 41244 4004 41300
rect 3836 40460 3892 40516
rect 3724 39394 3780 39396
rect 3724 39342 3726 39394
rect 3726 39342 3778 39394
rect 3778 39342 3780 39394
rect 3724 39340 3780 39342
rect 4172 39730 4228 39732
rect 4172 39678 4174 39730
rect 4174 39678 4226 39730
rect 4226 39678 4228 39730
rect 4172 39676 4228 39678
rect 4284 42252 4340 42308
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 3388 37660 3444 37716
rect 3276 37436 3332 37492
rect 3052 36540 3108 36596
rect 2156 36428 2212 36484
rect 2828 36428 2884 36484
rect 1708 35980 1764 36036
rect 2380 36258 2436 36260
rect 2380 36206 2382 36258
rect 2382 36206 2434 36258
rect 2434 36206 2436 36258
rect 2380 36204 2436 36206
rect 2604 36258 2660 36260
rect 2604 36206 2606 36258
rect 2606 36206 2658 36258
rect 2658 36206 2660 36258
rect 2604 36204 2660 36206
rect 1372 33852 1428 33908
rect 1932 34412 1988 34468
rect 2156 34972 2212 35028
rect 2156 34524 2212 34580
rect 2044 33964 2100 34020
rect 1932 33570 1988 33572
rect 1932 33518 1934 33570
rect 1934 33518 1986 33570
rect 1986 33518 1988 33570
rect 1932 33516 1988 33518
rect 3052 35420 3108 35476
rect 3612 36988 3668 37044
rect 4396 39340 4452 39396
rect 4732 39394 4788 39396
rect 4732 39342 4734 39394
rect 4734 39342 4786 39394
rect 4786 39342 4788 39394
rect 4732 39340 4788 39342
rect 4732 38946 4788 38948
rect 4732 38894 4734 38946
rect 4734 38894 4786 38946
rect 4786 38894 4788 38946
rect 4732 38892 4788 38894
rect 4396 38780 4452 38836
rect 3948 36204 4004 36260
rect 2492 34860 2548 34916
rect 2380 34300 2436 34356
rect 2604 34748 2660 34804
rect 2156 33516 2212 33572
rect 1820 32620 1876 32676
rect 1820 32396 1876 32452
rect 2156 33068 2212 33124
rect 2380 33068 2436 33124
rect 2492 33964 2548 34020
rect 2268 32620 2324 32676
rect 2492 32620 2548 32676
rect 2380 32396 2436 32452
rect 2156 31778 2212 31780
rect 2156 31726 2158 31778
rect 2158 31726 2210 31778
rect 2210 31726 2212 31778
rect 2156 31724 2212 31726
rect 2156 31106 2212 31108
rect 2156 31054 2158 31106
rect 2158 31054 2210 31106
rect 2210 31054 2212 31106
rect 2156 31052 2212 31054
rect 1260 28028 1316 28084
rect 1596 30940 1652 30996
rect 1148 16156 1204 16212
rect 1260 27580 1316 27636
rect 2044 29596 2100 29652
rect 1708 28812 1764 28868
rect 1932 28700 1988 28756
rect 1820 28642 1876 28644
rect 1820 28590 1822 28642
rect 1822 28590 1874 28642
rect 1874 28590 1876 28642
rect 1820 28588 1876 28590
rect 1932 27916 1988 27972
rect 1932 27132 1988 27188
rect 2268 28812 2324 28868
rect 2380 28700 2436 28756
rect 2268 28364 2324 28420
rect 3612 34748 3668 34804
rect 2940 34300 2996 34356
rect 3388 34242 3444 34244
rect 3388 34190 3390 34242
rect 3390 34190 3442 34242
rect 3442 34190 3444 34242
rect 3388 34188 3444 34190
rect 2716 33516 2772 33572
rect 2828 31948 2884 32004
rect 2940 31836 2996 31892
rect 2604 28364 2660 28420
rect 2716 30940 2772 30996
rect 2268 27804 2324 27860
rect 2828 31724 2884 31780
rect 3164 32060 3220 32116
rect 2716 27132 2772 27188
rect 1708 24892 1764 24948
rect 1372 24556 1428 24612
rect 1484 23772 1540 23828
rect 2156 26348 2212 26404
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 2044 23378 2100 23380
rect 2044 23326 2046 23378
rect 2046 23326 2098 23378
rect 2098 23326 2100 23378
rect 2044 23324 2100 23326
rect 1708 22764 1764 22820
rect 1708 22540 1764 22596
rect 1708 21868 1764 21924
rect 1820 21756 1876 21812
rect 1932 20076 1988 20132
rect 2156 21868 2212 21924
rect 2156 20300 2212 20356
rect 2380 25394 2436 25396
rect 2380 25342 2382 25394
rect 2382 25342 2434 25394
rect 2434 25342 2436 25394
rect 2380 25340 2436 25342
rect 2604 25004 2660 25060
rect 2492 24892 2548 24948
rect 3612 34188 3668 34244
rect 3612 32620 3668 32676
rect 3500 32060 3556 32116
rect 3276 31666 3332 31668
rect 3276 31614 3278 31666
rect 3278 31614 3330 31666
rect 3330 31614 3332 31666
rect 3276 31612 3332 31614
rect 3052 29932 3108 29988
rect 2940 28028 2996 28084
rect 3164 29260 3220 29316
rect 3724 30994 3780 30996
rect 3724 30942 3726 30994
rect 3726 30942 3778 30994
rect 3778 30942 3780 30994
rect 3724 30940 3780 30942
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 5292 46898 5348 46900
rect 5292 46846 5294 46898
rect 5294 46846 5346 46898
rect 5346 46846 5348 46898
rect 5292 46844 5348 46846
rect 5628 47180 5684 47236
rect 5516 44492 5572 44548
rect 5068 41916 5124 41972
rect 7420 52162 7476 52164
rect 7420 52110 7422 52162
rect 7422 52110 7474 52162
rect 7474 52110 7476 52162
rect 7420 52108 7476 52110
rect 7196 51884 7252 51940
rect 6860 51548 6916 51604
rect 6860 51266 6916 51268
rect 6860 51214 6862 51266
rect 6862 51214 6914 51266
rect 6914 51214 6916 51266
rect 6860 51212 6916 51214
rect 6748 50316 6804 50372
rect 6636 49980 6692 50036
rect 6860 50540 6916 50596
rect 7084 50594 7140 50596
rect 7084 50542 7086 50594
rect 7086 50542 7138 50594
rect 7138 50542 7140 50594
rect 7084 50540 7140 50542
rect 7084 49980 7140 50036
rect 7308 50034 7364 50036
rect 7308 49982 7310 50034
rect 7310 49982 7362 50034
rect 7362 49982 7364 50034
rect 7308 49980 7364 49982
rect 6188 46732 6244 46788
rect 5740 46002 5796 46004
rect 5740 45950 5742 46002
rect 5742 45950 5794 46002
rect 5794 45950 5796 46002
rect 5740 45948 5796 45950
rect 6300 45836 6356 45892
rect 5964 45052 6020 45108
rect 5740 44828 5796 44884
rect 5740 44434 5796 44436
rect 5740 44382 5742 44434
rect 5742 44382 5794 44434
rect 5794 44382 5796 44434
rect 5740 44380 5796 44382
rect 6076 44492 6132 44548
rect 6300 44380 6356 44436
rect 6524 47346 6580 47348
rect 6524 47294 6526 47346
rect 6526 47294 6578 47346
rect 6578 47294 6580 47346
rect 6524 47292 6580 47294
rect 6860 46786 6916 46788
rect 6860 46734 6862 46786
rect 6862 46734 6914 46786
rect 6914 46734 6916 46786
rect 6860 46732 6916 46734
rect 6748 45948 6804 46004
rect 6748 45778 6804 45780
rect 6748 45726 6750 45778
rect 6750 45726 6802 45778
rect 6802 45726 6804 45778
rect 6748 45724 6804 45726
rect 6636 45218 6692 45220
rect 6636 45166 6638 45218
rect 6638 45166 6690 45218
rect 6690 45166 6692 45218
rect 6636 45164 6692 45166
rect 6524 45052 6580 45108
rect 7532 48300 7588 48356
rect 7084 48076 7140 48132
rect 7420 47404 7476 47460
rect 7308 46844 7364 46900
rect 7868 50706 7924 50708
rect 7868 50654 7870 50706
rect 7870 50654 7922 50706
rect 7922 50654 7924 50706
rect 7868 50652 7924 50654
rect 8316 52668 8372 52724
rect 9100 53170 9156 53172
rect 9100 53118 9102 53170
rect 9102 53118 9154 53170
rect 9154 53118 9156 53170
rect 9100 53116 9156 53118
rect 8092 50652 8148 50708
rect 7756 49698 7812 49700
rect 7756 49646 7758 49698
rect 7758 49646 7810 49698
rect 7810 49646 7812 49698
rect 7756 49644 7812 49646
rect 7308 45330 7364 45332
rect 7308 45278 7310 45330
rect 7310 45278 7362 45330
rect 7362 45278 7364 45330
rect 7308 45276 7364 45278
rect 7420 45218 7476 45220
rect 7420 45166 7422 45218
rect 7422 45166 7474 45218
rect 7474 45166 7476 45218
rect 7420 45164 7476 45166
rect 7084 44828 7140 44884
rect 7196 44322 7252 44324
rect 7196 44270 7198 44322
rect 7198 44270 7250 44322
rect 7250 44270 7252 44322
rect 7196 44268 7252 44270
rect 6412 43596 6468 43652
rect 6300 43260 6356 43316
rect 5740 42812 5796 42868
rect 5964 42754 6020 42756
rect 5964 42702 5966 42754
rect 5966 42702 6018 42754
rect 6018 42702 6020 42754
rect 5964 42700 6020 42702
rect 6188 42476 6244 42532
rect 5740 42364 5796 42420
rect 5516 41804 5572 41860
rect 5292 39340 5348 39396
rect 5068 38946 5124 38948
rect 5068 38894 5070 38946
rect 5070 38894 5122 38946
rect 5122 38894 5124 38946
rect 5068 38892 5124 38894
rect 4956 38162 5012 38164
rect 4956 38110 4958 38162
rect 4958 38110 5010 38162
rect 5010 38110 5012 38162
rect 4956 38108 5012 38110
rect 4844 37772 4900 37828
rect 5068 37548 5124 37604
rect 4732 37324 4788 37380
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 5068 36876 5124 36932
rect 4396 36316 4452 36372
rect 4284 35756 4340 35812
rect 5404 38834 5460 38836
rect 5404 38782 5406 38834
rect 5406 38782 5458 38834
rect 5458 38782 5460 38834
rect 5404 38780 5460 38782
rect 6300 42364 6356 42420
rect 6300 41970 6356 41972
rect 6300 41918 6302 41970
rect 6302 41918 6354 41970
rect 6354 41918 6356 41970
rect 6300 41916 6356 41918
rect 7084 43596 7140 43652
rect 6636 43484 6692 43540
rect 7084 43372 7140 43428
rect 7196 43148 7252 43204
rect 6860 42140 6916 42196
rect 6636 42082 6692 42084
rect 6636 42030 6638 42082
rect 6638 42030 6690 42082
rect 6690 42030 6692 42082
rect 6636 42028 6692 42030
rect 6972 42082 7028 42084
rect 6972 42030 6974 42082
rect 6974 42030 7026 42082
rect 7026 42030 7028 42082
rect 6972 42028 7028 42030
rect 6972 41692 7028 41748
rect 6860 41244 6916 41300
rect 6076 40908 6132 40964
rect 6076 39900 6132 39956
rect 6188 40572 6244 40628
rect 5628 39676 5684 39732
rect 6076 39730 6132 39732
rect 6076 39678 6078 39730
rect 6078 39678 6130 39730
rect 6130 39678 6132 39730
rect 6076 39676 6132 39678
rect 5964 38834 6020 38836
rect 5964 38782 5966 38834
rect 5966 38782 6018 38834
rect 6018 38782 6020 38834
rect 5964 38780 6020 38782
rect 6076 37436 6132 37492
rect 5740 37154 5796 37156
rect 5740 37102 5742 37154
rect 5742 37102 5794 37154
rect 5794 37102 5796 37154
rect 5740 37100 5796 37102
rect 5516 36876 5572 36932
rect 5628 36370 5684 36372
rect 5628 36318 5630 36370
rect 5630 36318 5682 36370
rect 5682 36318 5684 36370
rect 5628 36316 5684 36318
rect 5852 36204 5908 36260
rect 5404 35980 5460 36036
rect 4060 34018 4116 34020
rect 4060 33966 4062 34018
rect 4062 33966 4114 34018
rect 4114 33966 4116 34018
rect 4060 33964 4116 33966
rect 4172 34972 4228 35028
rect 4060 33404 4116 33460
rect 4060 33068 4116 33124
rect 4060 32562 4116 32564
rect 4060 32510 4062 32562
rect 4062 32510 4114 32562
rect 4114 32510 4116 32562
rect 4060 32508 4116 32510
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4844 34524 4900 34580
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4284 33516 4340 33572
rect 4844 32674 4900 32676
rect 4844 32622 4846 32674
rect 4846 32622 4898 32674
rect 4898 32622 4900 32674
rect 4844 32620 4900 32622
rect 4956 33292 5012 33348
rect 4172 32396 4228 32452
rect 4508 32450 4564 32452
rect 4508 32398 4510 32450
rect 4510 32398 4562 32450
rect 4562 32398 4564 32450
rect 4508 32396 4564 32398
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 5180 32060 5236 32116
rect 6412 39618 6468 39620
rect 6412 39566 6414 39618
rect 6414 39566 6466 39618
rect 6466 39566 6468 39618
rect 6412 39564 6468 39566
rect 6300 39506 6356 39508
rect 6300 39454 6302 39506
rect 6302 39454 6354 39506
rect 6354 39454 6356 39506
rect 6300 39452 6356 39454
rect 6412 37772 6468 37828
rect 6636 36988 6692 37044
rect 6524 36706 6580 36708
rect 6524 36654 6526 36706
rect 6526 36654 6578 36706
rect 6578 36654 6580 36706
rect 6524 36652 6580 36654
rect 8204 51100 8260 51156
rect 8316 50316 8372 50372
rect 9996 54572 10052 54628
rect 9660 54402 9716 54404
rect 9660 54350 9662 54402
rect 9662 54350 9714 54402
rect 9714 54350 9716 54402
rect 9660 54348 9716 54350
rect 10556 55074 10612 55076
rect 10556 55022 10558 55074
rect 10558 55022 10610 55074
rect 10610 55022 10612 55074
rect 10556 55020 10612 55022
rect 11004 55074 11060 55076
rect 11004 55022 11006 55074
rect 11006 55022 11058 55074
rect 11058 55022 11060 55074
rect 11004 55020 11060 55022
rect 11228 54796 11284 54852
rect 9660 53618 9716 53620
rect 9660 53566 9662 53618
rect 9662 53566 9714 53618
rect 9714 53566 9716 53618
rect 9660 53564 9716 53566
rect 10892 54348 10948 54404
rect 11004 54236 11060 54292
rect 10892 54124 10948 54180
rect 25340 60508 25396 60564
rect 16156 60172 16212 60228
rect 17948 60226 18004 60228
rect 17948 60174 17950 60226
rect 17950 60174 18002 60226
rect 18002 60174 18004 60226
rect 17948 60172 18004 60174
rect 13580 59890 13636 59892
rect 13580 59838 13582 59890
rect 13582 59838 13634 59890
rect 13634 59838 13636 59890
rect 13580 59836 13636 59838
rect 12908 58940 12964 58996
rect 12124 57372 12180 57428
rect 12684 57372 12740 57428
rect 12572 56140 12628 56196
rect 12572 55970 12628 55972
rect 12572 55918 12574 55970
rect 12574 55918 12626 55970
rect 12626 55918 12628 55970
rect 12572 55916 12628 55918
rect 11676 55468 11732 55524
rect 12684 55132 12740 55188
rect 11788 55020 11844 55076
rect 11676 54572 11732 54628
rect 11788 54236 11844 54292
rect 11452 53788 11508 53844
rect 11564 53676 11620 53732
rect 10220 53452 10276 53508
rect 9884 53228 9940 53284
rect 9100 52274 9156 52276
rect 9100 52222 9102 52274
rect 9102 52222 9154 52274
rect 9154 52222 9156 52274
rect 9100 52220 9156 52222
rect 10556 53506 10612 53508
rect 10556 53454 10558 53506
rect 10558 53454 10610 53506
rect 10610 53454 10612 53506
rect 10556 53452 10612 53454
rect 11228 53452 11284 53508
rect 10220 52220 10276 52276
rect 8764 51938 8820 51940
rect 8764 51886 8766 51938
rect 8766 51886 8818 51938
rect 8818 51886 8820 51938
rect 8764 51884 8820 51886
rect 10220 51884 10276 51940
rect 10108 51772 10164 51828
rect 8652 51602 8708 51604
rect 8652 51550 8654 51602
rect 8654 51550 8706 51602
rect 8706 51550 8708 51602
rect 8652 51548 8708 51550
rect 9100 50988 9156 51044
rect 8652 50092 8708 50148
rect 8540 49868 8596 49924
rect 8316 49308 8372 49364
rect 8316 48242 8372 48244
rect 8316 48190 8318 48242
rect 8318 48190 8370 48242
rect 8370 48190 8372 48242
rect 8316 48188 8372 48190
rect 8316 47628 8372 47684
rect 8316 47180 8372 47236
rect 8988 50482 9044 50484
rect 8988 50430 8990 50482
rect 8990 50430 9042 50482
rect 9042 50430 9044 50482
rect 8988 50428 9044 50430
rect 9548 50764 9604 50820
rect 9324 50652 9380 50708
rect 9436 50540 9492 50596
rect 9100 49980 9156 50036
rect 8876 49698 8932 49700
rect 8876 49646 8878 49698
rect 8878 49646 8930 49698
rect 8930 49646 8932 49698
rect 8876 49644 8932 49646
rect 8764 48636 8820 48692
rect 8428 47516 8484 47572
rect 8652 47292 8708 47348
rect 9212 47740 9268 47796
rect 8988 47068 9044 47124
rect 9212 47346 9268 47348
rect 9212 47294 9214 47346
rect 9214 47294 9266 47346
rect 9266 47294 9268 47346
rect 9212 47292 9268 47294
rect 8876 46732 8932 46788
rect 8764 45948 8820 46004
rect 7420 42252 7476 42308
rect 7532 43148 7588 43204
rect 7308 42140 7364 42196
rect 7532 42028 7588 42084
rect 7196 41804 7252 41860
rect 7084 41186 7140 41188
rect 7084 41134 7086 41186
rect 7086 41134 7138 41186
rect 7138 41134 7140 41186
rect 7084 41132 7140 41134
rect 7420 41356 7476 41412
rect 7084 40236 7140 40292
rect 7196 40684 7252 40740
rect 6972 39676 7028 39732
rect 6860 39618 6916 39620
rect 6860 39566 6862 39618
rect 6862 39566 6914 39618
rect 6914 39566 6916 39618
rect 6860 39564 6916 39566
rect 6748 35196 6804 35252
rect 6188 34914 6244 34916
rect 6188 34862 6190 34914
rect 6190 34862 6242 34914
rect 6242 34862 6244 34914
rect 6188 34860 6244 34862
rect 5964 34748 6020 34804
rect 6300 34748 6356 34804
rect 5628 34524 5684 34580
rect 5964 33516 6020 33572
rect 5404 32844 5460 32900
rect 4732 31948 4788 32004
rect 5068 31948 5124 32004
rect 3948 31724 4004 31780
rect 4284 31724 4340 31780
rect 3836 30156 3892 30212
rect 3948 31500 4004 31556
rect 3500 29986 3556 29988
rect 3500 29934 3502 29986
rect 3502 29934 3554 29986
rect 3554 29934 3556 29986
rect 3500 29932 3556 29934
rect 3388 28140 3444 28196
rect 3500 29148 3556 29204
rect 4844 31276 4900 31332
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4732 30044 4788 30100
rect 4732 29596 4788 29652
rect 4620 29260 4676 29316
rect 4508 29148 4564 29204
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4396 28812 4452 28868
rect 5852 32620 5908 32676
rect 5516 31724 5572 31780
rect 5964 32508 6020 32564
rect 6748 34972 6804 35028
rect 6860 34748 6916 34804
rect 6412 33964 6468 34020
rect 6524 32620 6580 32676
rect 6188 32002 6244 32004
rect 6188 31950 6190 32002
rect 6190 31950 6242 32002
rect 6242 31950 6244 32002
rect 6188 31948 6244 31950
rect 6188 31612 6244 31668
rect 6412 31724 6468 31780
rect 6188 31388 6244 31444
rect 5852 30940 5908 30996
rect 5628 30268 5684 30324
rect 5516 28812 5572 28868
rect 5740 30210 5796 30212
rect 5740 30158 5742 30210
rect 5742 30158 5794 30210
rect 5794 30158 5796 30210
rect 5740 30156 5796 30158
rect 5628 28588 5684 28644
rect 6076 30210 6132 30212
rect 6076 30158 6078 30210
rect 6078 30158 6130 30210
rect 6130 30158 6132 30210
rect 6076 30156 6132 30158
rect 6860 33516 6916 33572
rect 8204 45276 8260 45332
rect 7868 44380 7924 44436
rect 8316 44380 8372 44436
rect 8988 45612 9044 45668
rect 8764 45106 8820 45108
rect 8764 45054 8766 45106
rect 8766 45054 8818 45106
rect 8818 45054 8820 45106
rect 8764 45052 8820 45054
rect 8540 44268 8596 44324
rect 7980 42812 8036 42868
rect 8092 42476 8148 42532
rect 8316 42812 8372 42868
rect 8092 42082 8148 42084
rect 8092 42030 8094 42082
rect 8094 42030 8146 42082
rect 8146 42030 8148 42082
rect 8092 42028 8148 42030
rect 7868 41580 7924 41636
rect 7644 41244 7700 41300
rect 7532 41186 7588 41188
rect 7532 41134 7534 41186
rect 7534 41134 7586 41186
rect 7586 41134 7588 41186
rect 7532 41132 7588 41134
rect 7644 40908 7700 40964
rect 7532 40514 7588 40516
rect 7532 40462 7534 40514
rect 7534 40462 7586 40514
rect 7586 40462 7588 40514
rect 7532 40460 7588 40462
rect 7308 39676 7364 39732
rect 7756 40626 7812 40628
rect 7756 40574 7758 40626
rect 7758 40574 7810 40626
rect 7810 40574 7812 40626
rect 7756 40572 7812 40574
rect 8092 41020 8148 41076
rect 8316 42252 8372 42308
rect 8876 43650 8932 43652
rect 8876 43598 8878 43650
rect 8878 43598 8930 43650
rect 8930 43598 8932 43650
rect 8876 43596 8932 43598
rect 9996 50652 10052 50708
rect 9660 49868 9716 49924
rect 9548 47292 9604 47348
rect 10220 50764 10276 50820
rect 10108 50594 10164 50596
rect 10108 50542 10110 50594
rect 10110 50542 10162 50594
rect 10162 50542 10164 50594
rect 10108 50540 10164 50542
rect 9884 49084 9940 49140
rect 9660 47180 9716 47236
rect 9660 46956 9716 47012
rect 9548 46674 9604 46676
rect 9548 46622 9550 46674
rect 9550 46622 9602 46674
rect 9602 46622 9604 46674
rect 9548 46620 9604 46622
rect 9884 47740 9940 47796
rect 9772 46844 9828 46900
rect 9884 47068 9940 47124
rect 10668 50540 10724 50596
rect 10444 50370 10500 50372
rect 10444 50318 10446 50370
rect 10446 50318 10498 50370
rect 10498 50318 10500 50370
rect 10444 50316 10500 50318
rect 10444 49138 10500 49140
rect 10444 49086 10446 49138
rect 10446 49086 10498 49138
rect 10498 49086 10500 49138
rect 10444 49084 10500 49086
rect 10556 48188 10612 48244
rect 10556 47516 10612 47572
rect 10108 46956 10164 47012
rect 10332 47180 10388 47236
rect 10220 46844 10276 46900
rect 9660 45666 9716 45668
rect 9660 45614 9662 45666
rect 9662 45614 9714 45666
rect 9714 45614 9716 45666
rect 9660 45612 9716 45614
rect 10108 45836 10164 45892
rect 9772 45500 9828 45556
rect 9548 45106 9604 45108
rect 9548 45054 9550 45106
rect 9550 45054 9602 45106
rect 9602 45054 9604 45106
rect 9548 45052 9604 45054
rect 9324 44492 9380 44548
rect 9100 43596 9156 43652
rect 9660 43650 9716 43652
rect 9660 43598 9662 43650
rect 9662 43598 9714 43650
rect 9714 43598 9716 43650
rect 9660 43596 9716 43598
rect 9884 43596 9940 43652
rect 8988 43538 9044 43540
rect 8988 43486 8990 43538
rect 8990 43486 9042 43538
rect 9042 43486 9044 43538
rect 8988 43484 9044 43486
rect 9548 43538 9604 43540
rect 9548 43486 9550 43538
rect 9550 43486 9602 43538
rect 9602 43486 9604 43538
rect 9548 43484 9604 43486
rect 8876 43314 8932 43316
rect 8876 43262 8878 43314
rect 8878 43262 8930 43314
rect 8930 43262 8932 43314
rect 8876 43260 8932 43262
rect 8652 42364 8708 42420
rect 10668 47180 10724 47236
rect 10444 46786 10500 46788
rect 10444 46734 10446 46786
rect 10446 46734 10498 46786
rect 10498 46734 10500 46786
rect 10444 46732 10500 46734
rect 12348 55074 12404 55076
rect 12348 55022 12350 55074
rect 12350 55022 12402 55074
rect 12402 55022 12404 55074
rect 12348 55020 12404 55022
rect 12124 54402 12180 54404
rect 12124 54350 12126 54402
rect 12126 54350 12178 54402
rect 12178 54350 12180 54402
rect 12124 54348 12180 54350
rect 12236 54290 12292 54292
rect 12236 54238 12238 54290
rect 12238 54238 12290 54290
rect 12290 54238 12292 54290
rect 12236 54236 12292 54238
rect 12460 53900 12516 53956
rect 11900 53564 11956 53620
rect 12348 53618 12404 53620
rect 12348 53566 12350 53618
rect 12350 53566 12402 53618
rect 12402 53566 12404 53618
rect 12348 53564 12404 53566
rect 12796 54514 12852 54516
rect 12796 54462 12798 54514
rect 12798 54462 12850 54514
rect 12850 54462 12852 54514
rect 12796 54460 12852 54462
rect 11228 50876 11284 50932
rect 11004 49250 11060 49252
rect 11004 49198 11006 49250
rect 11006 49198 11058 49250
rect 11058 49198 11060 49250
rect 11004 49196 11060 49198
rect 11340 48860 11396 48916
rect 10892 47516 10948 47572
rect 11228 47628 11284 47684
rect 11116 46844 11172 46900
rect 10892 46732 10948 46788
rect 10220 44380 10276 44436
rect 10332 44492 10388 44548
rect 10220 44044 10276 44100
rect 9996 43484 10052 43540
rect 10108 43372 10164 43428
rect 9884 42588 9940 42644
rect 8652 41970 8708 41972
rect 8652 41918 8654 41970
rect 8654 41918 8706 41970
rect 8706 41918 8708 41970
rect 8652 41916 8708 41918
rect 8876 41804 8932 41860
rect 8764 41580 8820 41636
rect 8316 41186 8372 41188
rect 8316 41134 8318 41186
rect 8318 41134 8370 41186
rect 8370 41134 8372 41186
rect 8316 41132 8372 41134
rect 9772 41858 9828 41860
rect 9772 41806 9774 41858
rect 9774 41806 9826 41858
rect 9826 41806 9828 41858
rect 9772 41804 9828 41806
rect 8092 40460 8148 40516
rect 7868 39788 7924 39844
rect 7308 38668 7364 38724
rect 9548 41074 9604 41076
rect 9548 41022 9550 41074
rect 9550 41022 9602 41074
rect 9602 41022 9604 41074
rect 9548 41020 9604 41022
rect 8540 39676 8596 39732
rect 8876 40236 8932 40292
rect 7868 39618 7924 39620
rect 7868 39566 7870 39618
rect 7870 39566 7922 39618
rect 7922 39566 7924 39618
rect 7868 39564 7924 39566
rect 10332 42642 10388 42644
rect 10332 42590 10334 42642
rect 10334 42590 10386 42642
rect 10386 42590 10388 42642
rect 10332 42588 10388 42590
rect 10108 41692 10164 41748
rect 9884 41356 9940 41412
rect 9772 40962 9828 40964
rect 9772 40910 9774 40962
rect 9774 40910 9826 40962
rect 9826 40910 9828 40962
rect 9772 40908 9828 40910
rect 10332 40626 10388 40628
rect 10332 40574 10334 40626
rect 10334 40574 10386 40626
rect 10386 40574 10388 40626
rect 10332 40572 10388 40574
rect 9884 40348 9940 40404
rect 9772 39788 9828 39844
rect 8540 39452 8596 39508
rect 7196 36652 7252 36708
rect 7084 35756 7140 35812
rect 7868 37660 7924 37716
rect 7980 37324 8036 37380
rect 7196 35868 7252 35924
rect 7084 33906 7140 33908
rect 7084 33854 7086 33906
rect 7086 33854 7138 33906
rect 7138 33854 7140 33906
rect 7084 33852 7140 33854
rect 8652 39116 8708 39172
rect 7420 35644 7476 35700
rect 7756 35756 7812 35812
rect 7980 35810 8036 35812
rect 7980 35758 7982 35810
rect 7982 35758 8034 35810
rect 8034 35758 8036 35810
rect 7980 35756 8036 35758
rect 8652 38050 8708 38052
rect 8652 37998 8654 38050
rect 8654 37998 8706 38050
rect 8706 37998 8708 38050
rect 8652 37996 8708 37998
rect 8316 37660 8372 37716
rect 8652 37490 8708 37492
rect 8652 37438 8654 37490
rect 8654 37438 8706 37490
rect 8706 37438 8708 37490
rect 8652 37436 8708 37438
rect 7644 35308 7700 35364
rect 7308 34860 7364 34916
rect 7420 35196 7476 35252
rect 7084 33458 7140 33460
rect 7084 33406 7086 33458
rect 7086 33406 7138 33458
rect 7138 33406 7140 33458
rect 7084 33404 7140 33406
rect 7196 33346 7252 33348
rect 7196 33294 7198 33346
rect 7198 33294 7250 33346
rect 7250 33294 7252 33346
rect 7196 33292 7252 33294
rect 6636 31164 6692 31220
rect 6300 29260 6356 29316
rect 6188 29148 6244 29204
rect 4508 28140 4564 28196
rect 2940 25676 2996 25732
rect 2940 24444 2996 24500
rect 2604 23884 2660 23940
rect 2604 22540 2660 22596
rect 2492 21532 2548 21588
rect 1484 18396 1540 18452
rect 1596 18620 1652 18676
rect 1372 16716 1428 16772
rect 1260 15484 1316 15540
rect 2044 18508 2100 18564
rect 2044 17778 2100 17780
rect 2044 17726 2046 17778
rect 2046 17726 2098 17778
rect 2098 17726 2100 17778
rect 2044 17724 2100 17726
rect 2268 18172 2324 18228
rect 2268 16716 2324 16772
rect 2268 15932 2324 15988
rect 2604 20748 2660 20804
rect 2716 20972 2772 21028
rect 2604 20578 2660 20580
rect 2604 20526 2606 20578
rect 2606 20526 2658 20578
rect 2658 20526 2660 20578
rect 2604 20524 2660 20526
rect 2492 20300 2548 20356
rect 4060 27916 4116 27972
rect 3724 27858 3780 27860
rect 3724 27806 3726 27858
rect 3726 27806 3778 27858
rect 3778 27806 3780 27858
rect 3724 27804 3780 27806
rect 3948 27804 4004 27860
rect 3500 26348 3556 26404
rect 3500 25452 3556 25508
rect 4508 27970 4564 27972
rect 4508 27918 4510 27970
rect 4510 27918 4562 27970
rect 4562 27918 4564 27970
rect 4508 27916 4564 27918
rect 5516 28028 5572 28084
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4060 27020 4116 27076
rect 4620 27074 4676 27076
rect 4620 27022 4622 27074
rect 4622 27022 4674 27074
rect 4674 27022 4676 27074
rect 4620 27020 4676 27022
rect 4732 26962 4788 26964
rect 4732 26910 4734 26962
rect 4734 26910 4786 26962
rect 4786 26910 4788 26962
rect 4732 26908 4788 26910
rect 5628 27858 5684 27860
rect 5628 27806 5630 27858
rect 5630 27806 5682 27858
rect 5682 27806 5684 27858
rect 5628 27804 5684 27806
rect 4844 26236 4900 26292
rect 4284 26124 4340 26180
rect 3836 25004 3892 25060
rect 3500 24668 3556 24724
rect 3836 24220 3892 24276
rect 3724 23548 3780 23604
rect 3164 23100 3220 23156
rect 3052 21532 3108 21588
rect 3164 22764 3220 22820
rect 3052 20802 3108 20804
rect 3052 20750 3054 20802
rect 3054 20750 3106 20802
rect 3106 20750 3108 20802
rect 3052 20748 3108 20750
rect 2940 19740 2996 19796
rect 2716 18450 2772 18452
rect 2716 18398 2718 18450
rect 2718 18398 2770 18450
rect 2770 18398 2772 18450
rect 2716 18396 2772 18398
rect 3052 17836 3108 17892
rect 2828 17276 2884 17332
rect 2604 17106 2660 17108
rect 2604 17054 2606 17106
rect 2606 17054 2658 17106
rect 2658 17054 2660 17106
rect 2604 17052 2660 17054
rect 2716 15596 2772 15652
rect 2716 15372 2772 15428
rect 2492 14642 2548 14644
rect 2492 14590 2494 14642
rect 2494 14590 2546 14642
rect 2546 14590 2548 14642
rect 2492 14588 2548 14590
rect 3500 23154 3556 23156
rect 3500 23102 3502 23154
rect 3502 23102 3554 23154
rect 3554 23102 3556 23154
rect 3500 23100 3556 23102
rect 3500 22876 3556 22932
rect 3388 21868 3444 21924
rect 3276 21026 3332 21028
rect 3276 20974 3278 21026
rect 3278 20974 3330 21026
rect 3330 20974 3332 21026
rect 3276 20972 3332 20974
rect 3276 19404 3332 19460
rect 2380 13804 2436 13860
rect 1932 13132 1988 13188
rect 2940 14306 2996 14308
rect 2940 14254 2942 14306
rect 2942 14254 2994 14306
rect 2994 14254 2996 14306
rect 2940 14252 2996 14254
rect 3164 15932 3220 15988
rect 3500 21698 3556 21700
rect 3500 21646 3502 21698
rect 3502 21646 3554 21698
rect 3554 21646 3556 21698
rect 3500 21644 3556 21646
rect 3612 18732 3668 18788
rect 3612 18450 3668 18452
rect 3612 18398 3614 18450
rect 3614 18398 3666 18450
rect 3666 18398 3668 18450
rect 3612 18396 3668 18398
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25394 4340 25396
rect 4284 25342 4286 25394
rect 4286 25342 4338 25394
rect 4338 25342 4340 25394
rect 4284 25340 4340 25342
rect 4396 25564 4452 25620
rect 4956 25564 5012 25620
rect 4060 24780 4116 24836
rect 4732 24780 4788 24836
rect 5628 26402 5684 26404
rect 5628 26350 5630 26402
rect 5630 26350 5682 26402
rect 5682 26350 5684 26402
rect 5628 26348 5684 26350
rect 5964 26236 6020 26292
rect 5516 26124 5572 26180
rect 5852 26178 5908 26180
rect 5852 26126 5854 26178
rect 5854 26126 5906 26178
rect 5906 26126 5908 26178
rect 5852 26124 5908 26126
rect 5740 25676 5796 25732
rect 5292 25228 5348 25284
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4060 23938 4116 23940
rect 4060 23886 4062 23938
rect 4062 23886 4114 23938
rect 4114 23886 4116 23938
rect 4060 23884 4116 23886
rect 3948 21756 4004 21812
rect 4060 23212 4116 23268
rect 3948 20802 4004 20804
rect 3948 20750 3950 20802
rect 3950 20750 4002 20802
rect 4002 20750 4004 20802
rect 3948 20748 4004 20750
rect 4620 22988 4676 23044
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4284 21756 4340 21812
rect 4620 22316 4676 22372
rect 5068 24050 5124 24052
rect 5068 23998 5070 24050
rect 5070 23998 5122 24050
rect 5122 23998 5124 24050
rect 5068 23996 5124 23998
rect 5068 22146 5124 22148
rect 5068 22094 5070 22146
rect 5070 22094 5122 22146
rect 5122 22094 5124 22146
rect 5068 22092 5124 22094
rect 5180 21756 5236 21812
rect 4172 21644 4228 21700
rect 4172 21026 4228 21028
rect 4172 20974 4174 21026
rect 4174 20974 4226 21026
rect 4226 20974 4228 21026
rect 4172 20972 4228 20974
rect 4396 21532 4452 21588
rect 4732 21474 4788 21476
rect 4732 21422 4734 21474
rect 4734 21422 4786 21474
rect 4786 21422 4788 21474
rect 4732 21420 4788 21422
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3948 20524 4004 20580
rect 3724 17724 3780 17780
rect 3836 19740 3892 19796
rect 3948 18508 4004 18564
rect 3948 18172 4004 18228
rect 3948 17106 4004 17108
rect 3948 17054 3950 17106
rect 3950 17054 4002 17106
rect 4002 17054 4004 17106
rect 3948 17052 4004 17054
rect 3388 15372 3444 15428
rect 3388 15202 3444 15204
rect 3388 15150 3390 15202
rect 3390 15150 3442 15202
rect 3442 15150 3444 15202
rect 3388 15148 3444 15150
rect 3612 16210 3668 16212
rect 3612 16158 3614 16210
rect 3614 16158 3666 16210
rect 3666 16158 3668 16210
rect 3612 16156 3668 16158
rect 5180 20578 5236 20580
rect 5180 20526 5182 20578
rect 5182 20526 5234 20578
rect 5234 20526 5236 20578
rect 5180 20524 5236 20526
rect 5852 25282 5908 25284
rect 5852 25230 5854 25282
rect 5854 25230 5906 25282
rect 5906 25230 5908 25282
rect 5852 25228 5908 25230
rect 5964 25116 6020 25172
rect 5628 24834 5684 24836
rect 5628 24782 5630 24834
rect 5630 24782 5682 24834
rect 5682 24782 5684 24834
rect 5628 24780 5684 24782
rect 5852 25004 5908 25060
rect 5852 24722 5908 24724
rect 5852 24670 5854 24722
rect 5854 24670 5906 24722
rect 5906 24670 5908 24722
rect 5852 24668 5908 24670
rect 5852 23548 5908 23604
rect 5628 22988 5684 23044
rect 5404 22092 5460 22148
rect 5740 20972 5796 21028
rect 5516 20860 5572 20916
rect 5180 20130 5236 20132
rect 5180 20078 5182 20130
rect 5182 20078 5234 20130
rect 5234 20078 5236 20130
rect 5180 20076 5236 20078
rect 5292 19964 5348 20020
rect 4620 19740 4676 19796
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4732 19068 4788 19124
rect 4956 19740 5012 19796
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4396 17612 4452 17668
rect 4396 17106 4452 17108
rect 4396 17054 4398 17106
rect 4398 17054 4450 17106
rect 4450 17054 4452 17106
rect 4396 17052 4452 17054
rect 4956 19516 5012 19572
rect 4956 17612 5012 17668
rect 4956 17442 5012 17444
rect 4956 17390 4958 17442
rect 4958 17390 5010 17442
rect 5010 17390 5012 17442
rect 4956 17388 5012 17390
rect 4284 16828 4340 16884
rect 4060 16156 4116 16212
rect 4172 16268 4228 16324
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 5180 16380 5236 16436
rect 4732 16268 4788 16324
rect 5628 19122 5684 19124
rect 5628 19070 5630 19122
rect 5630 19070 5682 19122
rect 5682 19070 5684 19122
rect 5628 19068 5684 19070
rect 5516 18284 5572 18340
rect 5628 17724 5684 17780
rect 6300 28082 6356 28084
rect 6300 28030 6302 28082
rect 6302 28030 6354 28082
rect 6354 28030 6356 28082
rect 6300 28028 6356 28030
rect 6188 27468 6244 27524
rect 6188 27186 6244 27188
rect 6188 27134 6190 27186
rect 6190 27134 6242 27186
rect 6242 27134 6244 27186
rect 6188 27132 6244 27134
rect 6860 31666 6916 31668
rect 6860 31614 6862 31666
rect 6862 31614 6914 31666
rect 6914 31614 6916 31666
rect 6860 31612 6916 31614
rect 6972 31554 7028 31556
rect 6972 31502 6974 31554
rect 6974 31502 7026 31554
rect 7026 31502 7028 31554
rect 6972 31500 7028 31502
rect 6860 31388 6916 31444
rect 7084 30828 7140 30884
rect 6860 29932 6916 29988
rect 7084 30492 7140 30548
rect 6972 29314 7028 29316
rect 6972 29262 6974 29314
rect 6974 29262 7026 29314
rect 7026 29262 7028 29314
rect 6972 29260 7028 29262
rect 7532 34972 7588 35028
rect 7868 34748 7924 34804
rect 7756 34524 7812 34580
rect 7644 33516 7700 33572
rect 7532 33292 7588 33348
rect 8540 35698 8596 35700
rect 8540 35646 8542 35698
rect 8542 35646 8594 35698
rect 8594 35646 8596 35698
rect 8540 35644 8596 35646
rect 9996 39618 10052 39620
rect 9996 39566 9998 39618
rect 9998 39566 10050 39618
rect 10050 39566 10052 39618
rect 9996 39564 10052 39566
rect 9772 38892 9828 38948
rect 9548 38050 9604 38052
rect 9548 37998 9550 38050
rect 9550 37998 9602 38050
rect 9602 37998 9604 38050
rect 9548 37996 9604 37998
rect 9100 37938 9156 37940
rect 9100 37886 9102 37938
rect 9102 37886 9154 37938
rect 9154 37886 9156 37938
rect 9100 37884 9156 37886
rect 9324 37826 9380 37828
rect 9324 37774 9326 37826
rect 9326 37774 9378 37826
rect 9378 37774 9380 37826
rect 9324 37772 9380 37774
rect 8988 37378 9044 37380
rect 8988 37326 8990 37378
rect 8990 37326 9042 37378
rect 9042 37326 9044 37378
rect 8988 37324 9044 37326
rect 9996 38668 10052 38724
rect 10108 38780 10164 38836
rect 11004 46060 11060 46116
rect 10780 45724 10836 45780
rect 10556 45218 10612 45220
rect 10556 45166 10558 45218
rect 10558 45166 10610 45218
rect 10610 45166 10612 45218
rect 10556 45164 10612 45166
rect 10780 45052 10836 45108
rect 10892 44322 10948 44324
rect 10892 44270 10894 44322
rect 10894 44270 10946 44322
rect 10946 44270 10948 44322
rect 10892 44268 10948 44270
rect 11676 52668 11732 52724
rect 11676 51884 11732 51940
rect 12572 51772 12628 51828
rect 11788 51548 11844 51604
rect 11564 51212 11620 51268
rect 12684 51266 12740 51268
rect 12684 51214 12686 51266
rect 12686 51214 12738 51266
rect 12738 51214 12740 51266
rect 12684 51212 12740 51214
rect 14028 59836 14084 59892
rect 14140 59276 14196 59332
rect 13804 58940 13860 58996
rect 13804 58716 13860 58772
rect 13468 58658 13524 58660
rect 13468 58606 13470 58658
rect 13470 58606 13522 58658
rect 13522 58606 13524 58658
rect 13468 58604 13524 58606
rect 14812 59388 14868 59444
rect 14924 59330 14980 59332
rect 14924 59278 14926 59330
rect 14926 59278 14978 59330
rect 14978 59278 14980 59330
rect 14924 59276 14980 59278
rect 14476 58492 14532 58548
rect 15260 58828 15316 58884
rect 14140 58380 14196 58436
rect 13580 57820 13636 57876
rect 13132 56924 13188 56980
rect 14812 58156 14868 58212
rect 14588 57874 14644 57876
rect 14588 57822 14590 57874
rect 14590 57822 14642 57874
rect 14642 57822 14644 57874
rect 14588 57820 14644 57822
rect 13916 56924 13972 56980
rect 14028 57484 14084 57540
rect 14028 57036 14084 57092
rect 13020 56866 13076 56868
rect 13020 56814 13022 56866
rect 13022 56814 13074 56866
rect 13074 56814 13076 56866
rect 13020 56812 13076 56814
rect 13580 56866 13636 56868
rect 13580 56814 13582 56866
rect 13582 56814 13634 56866
rect 13634 56814 13636 56866
rect 13580 56812 13636 56814
rect 14140 56476 14196 56532
rect 13356 55916 13412 55972
rect 13244 54738 13300 54740
rect 13244 54686 13246 54738
rect 13246 54686 13298 54738
rect 13298 54686 13300 54738
rect 13244 54684 13300 54686
rect 12908 53730 12964 53732
rect 12908 53678 12910 53730
rect 12910 53678 12962 53730
rect 12962 53678 12964 53730
rect 12908 53676 12964 53678
rect 13020 54572 13076 54628
rect 13132 54514 13188 54516
rect 13132 54462 13134 54514
rect 13134 54462 13186 54514
rect 13186 54462 13188 54514
rect 13132 54460 13188 54462
rect 13244 53004 13300 53060
rect 11788 50764 11844 50820
rect 12348 50876 12404 50932
rect 11564 50540 11620 50596
rect 12012 50316 12068 50372
rect 11452 46396 11508 46452
rect 11452 46060 11508 46116
rect 11340 46002 11396 46004
rect 11340 45950 11342 46002
rect 11342 45950 11394 46002
rect 11394 45950 11396 46002
rect 11340 45948 11396 45950
rect 11228 45724 11284 45780
rect 11452 45612 11508 45668
rect 11900 48300 11956 48356
rect 11900 47404 11956 47460
rect 12348 50316 12404 50372
rect 12460 50764 12516 50820
rect 12796 51100 12852 51156
rect 12572 50652 12628 50708
rect 12124 49644 12180 49700
rect 12236 49084 12292 49140
rect 12684 50540 12740 50596
rect 13020 50594 13076 50596
rect 13020 50542 13022 50594
rect 13022 50542 13074 50594
rect 13074 50542 13076 50594
rect 13020 50540 13076 50542
rect 12572 48802 12628 48804
rect 12572 48750 12574 48802
rect 12574 48750 12626 48802
rect 12626 48750 12628 48802
rect 12572 48748 12628 48750
rect 13916 55020 13972 55076
rect 13916 54796 13972 54852
rect 13804 54626 13860 54628
rect 13804 54574 13806 54626
rect 13806 54574 13858 54626
rect 13858 54574 13860 54626
rect 13804 54572 13860 54574
rect 13916 54460 13972 54516
rect 13692 54124 13748 54180
rect 13580 54012 13636 54068
rect 13804 54012 13860 54068
rect 13692 53900 13748 53956
rect 13580 53506 13636 53508
rect 13580 53454 13582 53506
rect 13582 53454 13634 53506
rect 13634 53454 13636 53506
rect 13580 53452 13636 53454
rect 13804 53340 13860 53396
rect 13692 52834 13748 52836
rect 13692 52782 13694 52834
rect 13694 52782 13746 52834
rect 13746 52782 13748 52834
rect 13692 52780 13748 52782
rect 13468 52332 13524 52388
rect 13804 52556 13860 52612
rect 13692 52162 13748 52164
rect 13692 52110 13694 52162
rect 13694 52110 13746 52162
rect 13746 52110 13748 52162
rect 13692 52108 13748 52110
rect 13916 51996 13972 52052
rect 14364 56252 14420 56308
rect 14140 55186 14196 55188
rect 14140 55134 14142 55186
rect 14142 55134 14194 55186
rect 14194 55134 14196 55186
rect 14140 55132 14196 55134
rect 14252 55468 14308 55524
rect 14252 54514 14308 54516
rect 14252 54462 14254 54514
rect 14254 54462 14306 54514
rect 14306 54462 14308 54514
rect 14252 54460 14308 54462
rect 14700 56754 14756 56756
rect 14700 56702 14702 56754
rect 14702 56702 14754 56754
rect 14754 56702 14756 56754
rect 14700 56700 14756 56702
rect 14700 55970 14756 55972
rect 14700 55918 14702 55970
rect 14702 55918 14754 55970
rect 14754 55918 14756 55970
rect 14700 55916 14756 55918
rect 14588 55468 14644 55524
rect 15036 57650 15092 57652
rect 15036 57598 15038 57650
rect 15038 57598 15090 57650
rect 15090 57598 15092 57650
rect 15036 57596 15092 57598
rect 15932 58604 15988 58660
rect 15372 58380 15428 58436
rect 15820 58492 15876 58548
rect 15484 58156 15540 58212
rect 15484 57820 15540 57876
rect 15036 56978 15092 56980
rect 15036 56926 15038 56978
rect 15038 56926 15090 56978
rect 15090 56926 15092 56978
rect 15036 56924 15092 56926
rect 15372 56588 15428 56644
rect 15260 55356 15316 55412
rect 14364 53564 14420 53620
rect 14028 53116 14084 53172
rect 13356 51772 13412 51828
rect 13580 51884 13636 51940
rect 13468 51660 13524 51716
rect 13356 51212 13412 51268
rect 13356 50764 13412 50820
rect 14476 53116 14532 53172
rect 14140 52892 14196 52948
rect 13692 50876 13748 50932
rect 15596 57090 15652 57092
rect 15596 57038 15598 57090
rect 15598 57038 15650 57090
rect 15650 57038 15652 57090
rect 15596 57036 15652 57038
rect 15708 56476 15764 56532
rect 16044 58380 16100 58436
rect 16156 59442 16212 59444
rect 16156 59390 16158 59442
rect 16158 59390 16210 59442
rect 16210 59390 16212 59442
rect 16156 59388 16212 59390
rect 16268 59052 16324 59108
rect 16380 57932 16436 57988
rect 15932 57596 15988 57652
rect 16940 58156 16996 58212
rect 16940 57708 16996 57764
rect 16156 57148 16212 57204
rect 15596 56306 15652 56308
rect 15596 56254 15598 56306
rect 15598 56254 15650 56306
rect 15650 56254 15652 56306
rect 15596 56252 15652 56254
rect 15484 55410 15540 55412
rect 15484 55358 15486 55410
rect 15486 55358 15538 55410
rect 15538 55358 15540 55410
rect 15484 55356 15540 55358
rect 15484 55132 15540 55188
rect 14812 54348 14868 54404
rect 14700 53228 14756 53284
rect 14252 52220 14308 52276
rect 14476 52332 14532 52388
rect 14700 52108 14756 52164
rect 14812 52892 14868 52948
rect 14812 52668 14868 52724
rect 14476 51884 14532 51940
rect 14252 51548 14308 51604
rect 13804 50652 13860 50708
rect 14364 50594 14420 50596
rect 14364 50542 14366 50594
rect 14366 50542 14418 50594
rect 14418 50542 14420 50594
rect 14364 50540 14420 50542
rect 14700 51266 14756 51268
rect 14700 51214 14702 51266
rect 14702 51214 14754 51266
rect 14754 51214 14756 51266
rect 14700 51212 14756 51214
rect 13804 49868 13860 49924
rect 13916 49532 13972 49588
rect 13916 49196 13972 49252
rect 12908 48914 12964 48916
rect 12908 48862 12910 48914
rect 12910 48862 12962 48914
rect 12962 48862 12964 48914
rect 12908 48860 12964 48862
rect 12348 47964 12404 48020
rect 11676 46956 11732 47012
rect 11788 46620 11844 46676
rect 11676 45948 11732 46004
rect 11788 45612 11844 45668
rect 11564 45106 11620 45108
rect 11564 45054 11566 45106
rect 11566 45054 11618 45106
rect 11618 45054 11620 45106
rect 11564 45052 11620 45054
rect 11564 44828 11620 44884
rect 11004 43538 11060 43540
rect 11004 43486 11006 43538
rect 11006 43486 11058 43538
rect 11058 43486 11060 43538
rect 11004 43484 11060 43486
rect 10556 42754 10612 42756
rect 10556 42702 10558 42754
rect 10558 42702 10610 42754
rect 10610 42702 10612 42754
rect 10556 42700 10612 42702
rect 10780 41804 10836 41860
rect 11340 44380 11396 44436
rect 11676 43538 11732 43540
rect 11676 43486 11678 43538
rect 11678 43486 11730 43538
rect 11730 43486 11732 43538
rect 11676 43484 11732 43486
rect 12012 45612 12068 45668
rect 12348 45164 12404 45220
rect 12236 44434 12292 44436
rect 12236 44382 12238 44434
rect 12238 44382 12290 44434
rect 12290 44382 12292 44434
rect 12236 44380 12292 44382
rect 12796 48188 12852 48244
rect 12684 47458 12740 47460
rect 12684 47406 12686 47458
rect 12686 47406 12738 47458
rect 12738 47406 12740 47458
rect 12684 47404 12740 47406
rect 13132 48354 13188 48356
rect 13132 48302 13134 48354
rect 13134 48302 13186 48354
rect 13186 48302 13188 48354
rect 13132 48300 13188 48302
rect 13580 48524 13636 48580
rect 13132 46956 13188 47012
rect 13020 46898 13076 46900
rect 13020 46846 13022 46898
rect 13022 46846 13074 46898
rect 13074 46846 13076 46898
rect 13020 46844 13076 46846
rect 13468 47404 13524 47460
rect 13468 47234 13524 47236
rect 13468 47182 13470 47234
rect 13470 47182 13522 47234
rect 13522 47182 13524 47234
rect 13468 47180 13524 47182
rect 13804 47292 13860 47348
rect 12572 45948 12628 46004
rect 14140 49868 14196 49924
rect 14140 47852 14196 47908
rect 14476 49698 14532 49700
rect 14476 49646 14478 49698
rect 14478 49646 14530 49698
rect 14530 49646 14532 49698
rect 14476 49644 14532 49646
rect 14252 48300 14308 48356
rect 14028 46844 14084 46900
rect 14364 48860 14420 48916
rect 14812 49644 14868 49700
rect 14588 48524 14644 48580
rect 14700 48242 14756 48244
rect 14700 48190 14702 48242
rect 14702 48190 14754 48242
rect 14754 48190 14756 48242
rect 14700 48188 14756 48190
rect 14364 47292 14420 47348
rect 14700 47068 14756 47124
rect 14476 46844 14532 46900
rect 14700 46674 14756 46676
rect 14700 46622 14702 46674
rect 14702 46622 14754 46674
rect 14754 46622 14756 46674
rect 14700 46620 14756 46622
rect 14252 46508 14308 46564
rect 13020 45948 13076 46004
rect 13916 46060 13972 46116
rect 13468 45890 13524 45892
rect 13468 45838 13470 45890
rect 13470 45838 13522 45890
rect 13522 45838 13524 45890
rect 13468 45836 13524 45838
rect 12908 45778 12964 45780
rect 12908 45726 12910 45778
rect 12910 45726 12962 45778
rect 12962 45726 12964 45778
rect 12908 45724 12964 45726
rect 12796 45612 12852 45668
rect 13020 45500 13076 45556
rect 12460 43708 12516 43764
rect 12796 43596 12852 43652
rect 14252 46060 14308 46116
rect 14028 45388 14084 45444
rect 13804 45276 13860 45332
rect 12012 42588 12068 42644
rect 12012 41916 12068 41972
rect 11228 41692 11284 41748
rect 11900 41692 11956 41748
rect 11788 41132 11844 41188
rect 11340 41020 11396 41076
rect 11340 40402 11396 40404
rect 11340 40350 11342 40402
rect 11342 40350 11394 40402
rect 11394 40350 11396 40402
rect 11340 40348 11396 40350
rect 10556 38780 10612 38836
rect 10780 38780 10836 38836
rect 10220 37660 10276 37716
rect 9884 36988 9940 37044
rect 10108 36428 10164 36484
rect 8876 36204 8932 36260
rect 8876 35922 8932 35924
rect 8876 35870 8878 35922
rect 8878 35870 8930 35922
rect 8930 35870 8932 35922
rect 8876 35868 8932 35870
rect 9772 35698 9828 35700
rect 9772 35646 9774 35698
rect 9774 35646 9826 35698
rect 9826 35646 9828 35698
rect 9772 35644 9828 35646
rect 8092 34914 8148 34916
rect 8092 34862 8094 34914
rect 8094 34862 8146 34914
rect 8146 34862 8148 34914
rect 8092 34860 8148 34862
rect 8316 34690 8372 34692
rect 8316 34638 8318 34690
rect 8318 34638 8370 34690
rect 8370 34638 8372 34690
rect 8316 34636 8372 34638
rect 8652 34914 8708 34916
rect 8652 34862 8654 34914
rect 8654 34862 8706 34914
rect 8706 34862 8708 34914
rect 8652 34860 8708 34862
rect 8204 33740 8260 33796
rect 8092 33404 8148 33460
rect 8540 34748 8596 34804
rect 7868 33068 7924 33124
rect 7420 31500 7476 31556
rect 7532 30940 7588 30996
rect 7756 31666 7812 31668
rect 7756 31614 7758 31666
rect 7758 31614 7810 31666
rect 7810 31614 7812 31666
rect 7756 31612 7812 31614
rect 8428 33964 8484 34020
rect 8540 33180 8596 33236
rect 8652 34636 8708 34692
rect 9660 34914 9716 34916
rect 9660 34862 9662 34914
rect 9662 34862 9714 34914
rect 9714 34862 9716 34914
rect 9660 34860 9716 34862
rect 9100 34524 9156 34580
rect 8988 33852 9044 33908
rect 8764 33292 8820 33348
rect 9996 34914 10052 34916
rect 9996 34862 9998 34914
rect 9998 34862 10050 34914
rect 10050 34862 10052 34914
rect 9996 34860 10052 34862
rect 9996 33740 10052 33796
rect 10444 34524 10500 34580
rect 10780 35756 10836 35812
rect 10668 35698 10724 35700
rect 10668 35646 10670 35698
rect 10670 35646 10722 35698
rect 10722 35646 10724 35698
rect 10668 35644 10724 35646
rect 10556 35084 10612 35140
rect 10220 34300 10276 34356
rect 10556 34076 10612 34132
rect 11004 39618 11060 39620
rect 11004 39566 11006 39618
rect 11006 39566 11058 39618
rect 11058 39566 11060 39618
rect 11004 39564 11060 39566
rect 11788 39676 11844 39732
rect 11452 39618 11508 39620
rect 11452 39566 11454 39618
rect 11454 39566 11506 39618
rect 11506 39566 11508 39618
rect 11452 39564 11508 39566
rect 11004 38668 11060 38724
rect 11228 38834 11284 38836
rect 11228 38782 11230 38834
rect 11230 38782 11282 38834
rect 11282 38782 11284 38834
rect 11228 38780 11284 38782
rect 11788 38780 11844 38836
rect 11676 38722 11732 38724
rect 11676 38670 11678 38722
rect 11678 38670 11730 38722
rect 11730 38670 11732 38722
rect 11676 38668 11732 38670
rect 11116 37660 11172 37716
rect 11452 37660 11508 37716
rect 11340 37042 11396 37044
rect 11340 36990 11342 37042
rect 11342 36990 11394 37042
rect 11394 36990 11396 37042
rect 11340 36988 11396 36990
rect 11004 36482 11060 36484
rect 11004 36430 11006 36482
rect 11006 36430 11058 36482
rect 11058 36430 11060 36482
rect 11004 36428 11060 36430
rect 11004 35756 11060 35812
rect 11228 35868 11284 35924
rect 11564 36428 11620 36484
rect 11004 34972 11060 35028
rect 10220 33346 10276 33348
rect 10220 33294 10222 33346
rect 10222 33294 10274 33346
rect 10274 33294 10276 33346
rect 10220 33292 10276 33294
rect 10220 33122 10276 33124
rect 10220 33070 10222 33122
rect 10222 33070 10274 33122
rect 10274 33070 10276 33122
rect 10220 33068 10276 33070
rect 10108 32620 10164 32676
rect 10332 32956 10388 33012
rect 7980 31164 8036 31220
rect 7868 30994 7924 30996
rect 7868 30942 7870 30994
rect 7870 30942 7922 30994
rect 7922 30942 7924 30994
rect 7868 30940 7924 30942
rect 7644 30716 7700 30772
rect 7756 30492 7812 30548
rect 7868 30268 7924 30324
rect 7308 30210 7364 30212
rect 7308 30158 7310 30210
rect 7310 30158 7362 30210
rect 7362 30158 7364 30210
rect 7308 30156 7364 30158
rect 7420 30098 7476 30100
rect 7420 30046 7422 30098
rect 7422 30046 7474 30098
rect 7474 30046 7476 30098
rect 7420 30044 7476 30046
rect 7196 29708 7252 29764
rect 7756 29708 7812 29764
rect 8316 31164 8372 31220
rect 8092 30716 8148 30772
rect 7644 28588 7700 28644
rect 6748 27132 6804 27188
rect 7756 27186 7812 27188
rect 7756 27134 7758 27186
rect 7758 27134 7810 27186
rect 7810 27134 7812 27186
rect 7756 27132 7812 27134
rect 6972 26908 7028 26964
rect 6748 26796 6804 26852
rect 6748 26290 6804 26292
rect 6748 26238 6750 26290
rect 6750 26238 6802 26290
rect 6802 26238 6804 26290
rect 6748 26236 6804 26238
rect 6412 26124 6468 26180
rect 8540 31948 8596 32004
rect 9660 32060 9716 32116
rect 9212 31890 9268 31892
rect 9212 31838 9214 31890
rect 9214 31838 9266 31890
rect 9266 31838 9268 31890
rect 9212 31836 9268 31838
rect 8988 31778 9044 31780
rect 8988 31726 8990 31778
rect 8990 31726 9042 31778
rect 9042 31726 9044 31778
rect 8988 31724 9044 31726
rect 9100 31554 9156 31556
rect 9100 31502 9102 31554
rect 9102 31502 9154 31554
rect 9154 31502 9156 31554
rect 9100 31500 9156 31502
rect 9436 31500 9492 31556
rect 8764 31388 8820 31444
rect 8540 31276 8596 31332
rect 9772 31948 9828 32004
rect 9660 31276 9716 31332
rect 9772 31724 9828 31780
rect 10108 31164 10164 31220
rect 8876 30994 8932 30996
rect 8876 30942 8878 30994
rect 8878 30942 8930 30994
rect 8930 30942 8932 30994
rect 8876 30940 8932 30942
rect 8540 30098 8596 30100
rect 8540 30046 8542 30098
rect 8542 30046 8594 30098
rect 8594 30046 8596 30098
rect 8540 30044 8596 30046
rect 8428 28028 8484 28084
rect 8092 27580 8148 27636
rect 8092 27132 8148 27188
rect 7868 27074 7924 27076
rect 7868 27022 7870 27074
rect 7870 27022 7922 27074
rect 7922 27022 7924 27074
rect 7868 27020 7924 27022
rect 8204 26962 8260 26964
rect 8204 26910 8206 26962
rect 8206 26910 8258 26962
rect 8258 26910 8260 26962
rect 8204 26908 8260 26910
rect 9548 29148 9604 29204
rect 9436 28588 9492 28644
rect 9324 27244 9380 27300
rect 8988 26908 9044 26964
rect 7756 26290 7812 26292
rect 7756 26238 7758 26290
rect 7758 26238 7810 26290
rect 7810 26238 7812 26290
rect 7756 26236 7812 26238
rect 6748 25506 6804 25508
rect 6748 25454 6750 25506
rect 6750 25454 6802 25506
rect 6802 25454 6804 25506
rect 6748 25452 6804 25454
rect 6972 25228 7028 25284
rect 6748 24780 6804 24836
rect 6748 24498 6804 24500
rect 6748 24446 6750 24498
rect 6750 24446 6802 24498
rect 6802 24446 6804 24498
rect 6748 24444 6804 24446
rect 6636 24220 6692 24276
rect 6748 23938 6804 23940
rect 6748 23886 6750 23938
rect 6750 23886 6802 23938
rect 6802 23886 6804 23938
rect 6748 23884 6804 23886
rect 6076 22092 6132 22148
rect 6412 22876 6468 22932
rect 6636 23436 6692 23492
rect 6412 22092 6468 22148
rect 6188 21586 6244 21588
rect 6188 21534 6190 21586
rect 6190 21534 6242 21586
rect 6242 21534 6244 21586
rect 6188 21532 6244 21534
rect 5964 20748 6020 20804
rect 6076 20636 6132 20692
rect 6300 21420 6356 21476
rect 6524 20972 6580 21028
rect 6636 23100 6692 23156
rect 5964 19964 6020 20020
rect 5964 18396 6020 18452
rect 5516 16380 5572 16436
rect 5404 16268 5460 16324
rect 5180 16098 5236 16100
rect 5180 16046 5182 16098
rect 5182 16046 5234 16098
rect 5234 16046 5236 16098
rect 5180 16044 5236 16046
rect 4620 15932 4676 15988
rect 4956 15874 5012 15876
rect 4956 15822 4958 15874
rect 4958 15822 5010 15874
rect 5010 15822 5012 15874
rect 4956 15820 5012 15822
rect 3948 15708 4004 15764
rect 3836 15596 3892 15652
rect 3948 15148 4004 15204
rect 3500 14476 3556 14532
rect 3612 14700 3668 14756
rect 3500 14252 3556 14308
rect 2828 13132 2884 13188
rect 2044 13074 2100 13076
rect 2044 13022 2046 13074
rect 2046 13022 2098 13074
rect 2098 13022 2100 13074
rect 2044 13020 2100 13022
rect 3388 13020 3444 13076
rect 1708 11452 1764 11508
rect 2828 12066 2884 12068
rect 2828 12014 2830 12066
rect 2830 12014 2882 12066
rect 2882 12014 2884 12066
rect 2828 12012 2884 12014
rect 4284 15538 4340 15540
rect 4284 15486 4286 15538
rect 4286 15486 4338 15538
rect 4338 15486 4340 15538
rect 4284 15484 4340 15486
rect 5964 17164 6020 17220
rect 5852 17106 5908 17108
rect 5852 17054 5854 17106
rect 5854 17054 5906 17106
rect 5906 17054 5908 17106
rect 5852 17052 5908 17054
rect 6524 19964 6580 20020
rect 6636 20076 6692 20132
rect 6300 19740 6356 19796
rect 6412 19852 6468 19908
rect 6524 19628 6580 19684
rect 7756 25228 7812 25284
rect 7420 24780 7476 24836
rect 7532 24668 7588 24724
rect 7196 24220 7252 24276
rect 6972 24108 7028 24164
rect 7084 23938 7140 23940
rect 7084 23886 7086 23938
rect 7086 23886 7138 23938
rect 7138 23886 7140 23938
rect 7084 23884 7140 23886
rect 7980 24668 8036 24724
rect 7644 24108 7700 24164
rect 8204 24556 8260 24612
rect 8092 24162 8148 24164
rect 8092 24110 8094 24162
rect 8094 24110 8146 24162
rect 8146 24110 8148 24162
rect 8092 24108 8148 24110
rect 7420 23324 7476 23380
rect 6972 22370 7028 22372
rect 6972 22318 6974 22370
rect 6974 22318 7026 22370
rect 7026 22318 7028 22370
rect 6972 22316 7028 22318
rect 6972 20188 7028 20244
rect 7196 20018 7252 20020
rect 7196 19966 7198 20018
rect 7198 19966 7250 20018
rect 7250 19966 7252 20018
rect 7196 19964 7252 19966
rect 6972 19234 7028 19236
rect 6972 19182 6974 19234
rect 6974 19182 7026 19234
rect 7026 19182 7028 19234
rect 6972 19180 7028 19182
rect 6636 19068 6692 19124
rect 6748 19010 6804 19012
rect 6748 18958 6750 19010
rect 6750 18958 6802 19010
rect 6802 18958 6804 19010
rect 6748 18956 6804 18958
rect 6524 18450 6580 18452
rect 6524 18398 6526 18450
rect 6526 18398 6578 18450
rect 6578 18398 6580 18450
rect 6524 18396 6580 18398
rect 6748 18396 6804 18452
rect 6300 17442 6356 17444
rect 6300 17390 6302 17442
rect 6302 17390 6354 17442
rect 6354 17390 6356 17442
rect 6300 17388 6356 17390
rect 6860 17778 6916 17780
rect 6860 17726 6862 17778
rect 6862 17726 6914 17778
rect 6914 17726 6916 17778
rect 6860 17724 6916 17726
rect 6748 16940 6804 16996
rect 6972 16994 7028 16996
rect 6972 16942 6974 16994
rect 6974 16942 7026 16994
rect 7026 16942 7028 16994
rect 6972 16940 7028 16942
rect 6860 16882 6916 16884
rect 6860 16830 6862 16882
rect 6862 16830 6914 16882
rect 6914 16830 6916 16882
rect 6860 16828 6916 16830
rect 6300 16268 6356 16324
rect 6076 16098 6132 16100
rect 6076 16046 6078 16098
rect 6078 16046 6130 16098
rect 6130 16046 6132 16098
rect 6076 16044 6132 16046
rect 6188 16156 6244 16212
rect 5852 15820 5908 15876
rect 4732 15372 4788 15428
rect 4844 15314 4900 15316
rect 4844 15262 4846 15314
rect 4846 15262 4898 15314
rect 4898 15262 4900 15314
rect 4844 15260 4900 15262
rect 5516 15426 5572 15428
rect 5516 15374 5518 15426
rect 5518 15374 5570 15426
rect 5570 15374 5572 15426
rect 5516 15372 5572 15374
rect 5292 15260 5348 15316
rect 4172 14588 4228 14644
rect 4284 15036 4340 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5740 15148 5796 15204
rect 4732 14252 4788 14308
rect 4620 13916 4676 13972
rect 4060 13804 4116 13860
rect 3836 12908 3892 12964
rect 4844 13804 4900 13860
rect 4732 13468 4788 13524
rect 5068 14306 5124 14308
rect 5068 14254 5070 14306
rect 5070 14254 5122 14306
rect 5122 14254 5124 14306
rect 5068 14252 5124 14254
rect 5404 14140 5460 14196
rect 5180 13580 5236 13636
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4060 13020 4116 13076
rect 4060 12684 4116 12740
rect 5068 13020 5124 13076
rect 3500 12012 3556 12068
rect 2492 11506 2548 11508
rect 2492 11454 2494 11506
rect 2494 11454 2546 11506
rect 2546 11454 2548 11506
rect 2492 11452 2548 11454
rect 3724 12066 3780 12068
rect 3724 12014 3726 12066
rect 3726 12014 3778 12066
rect 3778 12014 3780 12066
rect 3724 12012 3780 12014
rect 4172 11954 4228 11956
rect 4172 11902 4174 11954
rect 4174 11902 4226 11954
rect 4226 11902 4228 11954
rect 4172 11900 4228 11902
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4956 11282 5012 11284
rect 4956 11230 4958 11282
rect 4958 11230 5010 11282
rect 5010 11230 5012 11282
rect 4956 11228 5012 11230
rect 5068 11116 5124 11172
rect 2044 10556 2100 10612
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 5516 14028 5572 14084
rect 5516 13692 5572 13748
rect 5628 13580 5684 13636
rect 6076 15314 6132 15316
rect 6076 15262 6078 15314
rect 6078 15262 6130 15314
rect 6130 15262 6132 15314
rect 6076 15260 6132 15262
rect 6412 15260 6468 15316
rect 5852 14812 5908 14868
rect 5852 14364 5908 14420
rect 5964 14140 6020 14196
rect 5852 13916 5908 13972
rect 6300 14642 6356 14644
rect 6300 14590 6302 14642
rect 6302 14590 6354 14642
rect 6354 14590 6356 14642
rect 6300 14588 6356 14590
rect 7532 21756 7588 21812
rect 8540 26460 8596 26516
rect 8540 26290 8596 26292
rect 8540 26238 8542 26290
rect 8542 26238 8594 26290
rect 8594 26238 8596 26290
rect 8540 26236 8596 26238
rect 8428 26178 8484 26180
rect 8428 26126 8430 26178
rect 8430 26126 8482 26178
rect 8482 26126 8484 26178
rect 8428 26124 8484 26126
rect 8428 25228 8484 25284
rect 9436 25116 9492 25172
rect 9548 27468 9604 27524
rect 8876 25004 8932 25060
rect 9884 29650 9940 29652
rect 9884 29598 9886 29650
rect 9886 29598 9938 29650
rect 9938 29598 9940 29650
rect 9884 29596 9940 29598
rect 10108 29372 10164 29428
rect 9996 27692 10052 27748
rect 9660 25618 9716 25620
rect 9660 25566 9662 25618
rect 9662 25566 9714 25618
rect 9714 25566 9716 25618
rect 9660 25564 9716 25566
rect 9548 24444 9604 24500
rect 8764 24108 8820 24164
rect 8876 24332 8932 24388
rect 9212 23714 9268 23716
rect 9212 23662 9214 23714
rect 9214 23662 9266 23714
rect 9266 23662 9268 23714
rect 9212 23660 9268 23662
rect 8764 23212 8820 23268
rect 8428 23154 8484 23156
rect 8428 23102 8430 23154
rect 8430 23102 8482 23154
rect 8482 23102 8484 23154
rect 8428 23100 8484 23102
rect 8092 23042 8148 23044
rect 8092 22990 8094 23042
rect 8094 22990 8146 23042
rect 8146 22990 8148 23042
rect 8092 22988 8148 22990
rect 8652 22370 8708 22372
rect 8652 22318 8654 22370
rect 8654 22318 8706 22370
rect 8706 22318 8708 22370
rect 8652 22316 8708 22318
rect 7532 20412 7588 20468
rect 7756 20914 7812 20916
rect 7756 20862 7758 20914
rect 7758 20862 7810 20914
rect 7810 20862 7812 20914
rect 7756 20860 7812 20862
rect 7756 20188 7812 20244
rect 8092 20636 8148 20692
rect 8316 20748 8372 20804
rect 7868 19964 7924 20020
rect 7756 19740 7812 19796
rect 7756 18844 7812 18900
rect 7420 17612 7476 17668
rect 8092 19180 8148 19236
rect 8316 20300 8372 20356
rect 8876 22204 8932 22260
rect 8540 20188 8596 20244
rect 9100 21532 9156 21588
rect 8988 20412 9044 20468
rect 8988 20130 9044 20132
rect 8988 20078 8990 20130
rect 8990 20078 9042 20130
rect 9042 20078 9044 20130
rect 8988 20076 9044 20078
rect 8652 19852 8708 19908
rect 9996 26402 10052 26404
rect 9996 26350 9998 26402
rect 9998 26350 10050 26402
rect 10050 26350 10052 26402
rect 9996 26348 10052 26350
rect 10556 33458 10612 33460
rect 10556 33406 10558 33458
rect 10558 33406 10610 33458
rect 10610 33406 10612 33458
rect 10556 33404 10612 33406
rect 12796 42588 12852 42644
rect 12684 42082 12740 42084
rect 12684 42030 12686 42082
rect 12686 42030 12738 42082
rect 12738 42030 12740 42082
rect 12684 42028 12740 42030
rect 12572 41244 12628 41300
rect 12124 41132 12180 41188
rect 12460 41074 12516 41076
rect 12460 41022 12462 41074
rect 12462 41022 12514 41074
rect 12514 41022 12516 41074
rect 12460 41020 12516 41022
rect 12012 40572 12068 40628
rect 12684 40962 12740 40964
rect 12684 40910 12686 40962
rect 12686 40910 12738 40962
rect 12738 40910 12740 40962
rect 12684 40908 12740 40910
rect 13244 41804 13300 41860
rect 12908 41244 12964 41300
rect 13244 40908 13300 40964
rect 12684 38892 12740 38948
rect 13132 40236 13188 40292
rect 12460 37212 12516 37268
rect 12684 37884 12740 37940
rect 12236 36988 12292 37044
rect 11900 36764 11956 36820
rect 11788 34354 11844 34356
rect 11788 34302 11790 34354
rect 11790 34302 11842 34354
rect 11842 34302 11844 34354
rect 11788 34300 11844 34302
rect 12012 35756 12068 35812
rect 12124 36204 12180 36260
rect 12348 35980 12404 36036
rect 10780 33234 10836 33236
rect 10780 33182 10782 33234
rect 10782 33182 10834 33234
rect 10834 33182 10836 33234
rect 10780 33180 10836 33182
rect 10892 32172 10948 32228
rect 10668 32060 10724 32116
rect 11228 32060 11284 32116
rect 12012 32732 12068 32788
rect 11564 32284 11620 32340
rect 11004 31554 11060 31556
rect 11004 31502 11006 31554
rect 11006 31502 11058 31554
rect 11058 31502 11060 31554
rect 11004 31500 11060 31502
rect 13356 40124 13412 40180
rect 13356 38892 13412 38948
rect 13244 38668 13300 38724
rect 13692 42642 13748 42644
rect 13692 42590 13694 42642
rect 13694 42590 13746 42642
rect 13746 42590 13748 42642
rect 13692 42588 13748 42590
rect 13916 41970 13972 41972
rect 13916 41918 13918 41970
rect 13918 41918 13970 41970
rect 13970 41918 13972 41970
rect 13916 41916 13972 41918
rect 14140 45052 14196 45108
rect 14140 43708 14196 43764
rect 14700 45164 14756 45220
rect 15148 53340 15204 53396
rect 15036 53058 15092 53060
rect 15036 53006 15038 53058
rect 15038 53006 15090 53058
rect 15090 53006 15092 53058
rect 15036 53004 15092 53006
rect 15148 52946 15204 52948
rect 15148 52894 15150 52946
rect 15150 52894 15202 52946
rect 15202 52894 15204 52946
rect 15148 52892 15204 52894
rect 15372 53116 15428 53172
rect 16492 56924 16548 56980
rect 15932 56082 15988 56084
rect 15932 56030 15934 56082
rect 15934 56030 15986 56082
rect 15986 56030 15988 56082
rect 15932 56028 15988 56030
rect 16156 55804 16212 55860
rect 15820 54348 15876 54404
rect 15932 54908 15988 54964
rect 19964 59890 20020 59892
rect 19964 59838 19966 59890
rect 19966 59838 20018 59890
rect 20018 59838 20020 59890
rect 19964 59836 20020 59838
rect 20860 59890 20916 59892
rect 20860 59838 20862 59890
rect 20862 59838 20914 59890
rect 20914 59838 20916 59890
rect 20860 59836 20916 59838
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 20300 59778 20356 59780
rect 20300 59726 20302 59778
rect 20302 59726 20354 59778
rect 20354 59726 20356 59778
rect 20300 59724 20356 59726
rect 17948 59330 18004 59332
rect 17948 59278 17950 59330
rect 17950 59278 18002 59330
rect 18002 59278 18004 59330
rect 17948 59276 18004 59278
rect 19516 58828 19572 58884
rect 17164 57932 17220 57988
rect 17052 56700 17108 56756
rect 16828 56476 16884 56532
rect 16716 56028 16772 56084
rect 17948 57708 18004 57764
rect 17836 57148 17892 57204
rect 18844 58044 18900 58100
rect 19180 57932 19236 57988
rect 18844 57820 18900 57876
rect 19404 57762 19460 57764
rect 19404 57710 19406 57762
rect 19406 57710 19458 57762
rect 19458 57710 19460 57762
rect 19404 57708 19460 57710
rect 18508 57036 18564 57092
rect 18172 56924 18228 56980
rect 17276 55580 17332 55636
rect 16268 55132 16324 55188
rect 16156 54572 16212 54628
rect 15596 53676 15652 53732
rect 15932 53788 15988 53844
rect 15484 53564 15540 53620
rect 15148 52722 15204 52724
rect 15148 52670 15150 52722
rect 15150 52670 15202 52722
rect 15202 52670 15204 52722
rect 15148 52668 15204 52670
rect 15372 52668 15428 52724
rect 15260 52274 15316 52276
rect 15260 52222 15262 52274
rect 15262 52222 15314 52274
rect 15314 52222 15316 52274
rect 15260 52220 15316 52222
rect 15036 52108 15092 52164
rect 16268 54348 16324 54404
rect 16156 54236 16212 54292
rect 16380 53900 16436 53956
rect 16268 53730 16324 53732
rect 16268 53678 16270 53730
rect 16270 53678 16322 53730
rect 16322 53678 16324 53730
rect 16268 53676 16324 53678
rect 15932 53004 15988 53060
rect 15820 52556 15876 52612
rect 15148 51548 15204 51604
rect 15484 51324 15540 51380
rect 15260 50652 15316 50708
rect 15484 49868 15540 49924
rect 15260 49420 15316 49476
rect 15372 49532 15428 49588
rect 15260 48748 15316 48804
rect 15484 49420 15540 49476
rect 15820 51212 15876 51268
rect 16044 52668 16100 52724
rect 16268 52108 16324 52164
rect 16156 51996 16212 52052
rect 16044 50764 16100 50820
rect 15708 50482 15764 50484
rect 15708 50430 15710 50482
rect 15710 50430 15762 50482
rect 15762 50430 15764 50482
rect 15708 50428 15764 50430
rect 15708 49810 15764 49812
rect 15708 49758 15710 49810
rect 15710 49758 15762 49810
rect 15762 49758 15764 49810
rect 15708 49756 15764 49758
rect 16380 51100 16436 51156
rect 16268 50652 16324 50708
rect 17388 54908 17444 54964
rect 17612 54626 17668 54628
rect 17612 54574 17614 54626
rect 17614 54574 17666 54626
rect 17666 54574 17668 54626
rect 17612 54572 17668 54574
rect 16604 53058 16660 53060
rect 16604 53006 16606 53058
rect 16606 53006 16658 53058
rect 16658 53006 16660 53058
rect 16604 53004 16660 53006
rect 16604 52556 16660 52612
rect 16828 53618 16884 53620
rect 16828 53566 16830 53618
rect 16830 53566 16882 53618
rect 16882 53566 16884 53618
rect 16828 53564 16884 53566
rect 16940 53506 16996 53508
rect 16940 53454 16942 53506
rect 16942 53454 16994 53506
rect 16994 53454 16996 53506
rect 16940 53452 16996 53454
rect 17500 54012 17556 54068
rect 17612 53788 17668 53844
rect 17276 53730 17332 53732
rect 17276 53678 17278 53730
rect 17278 53678 17330 53730
rect 17330 53678 17332 53730
rect 17276 53676 17332 53678
rect 17164 53618 17220 53620
rect 17164 53566 17166 53618
rect 17166 53566 17218 53618
rect 17218 53566 17220 53618
rect 17164 53564 17220 53566
rect 17052 53228 17108 53284
rect 17500 52892 17556 52948
rect 17388 52108 17444 52164
rect 16828 51436 16884 51492
rect 16044 49644 16100 49700
rect 16044 49420 16100 49476
rect 15484 47852 15540 47908
rect 15372 47346 15428 47348
rect 15372 47294 15374 47346
rect 15374 47294 15426 47346
rect 15426 47294 15428 47346
rect 15372 47292 15428 47294
rect 15484 47068 15540 47124
rect 15372 46844 15428 46900
rect 14924 45388 14980 45444
rect 15036 46508 15092 46564
rect 15372 46396 15428 46452
rect 15148 45890 15204 45892
rect 15148 45838 15150 45890
rect 15150 45838 15202 45890
rect 15202 45838 15204 45890
rect 15148 45836 15204 45838
rect 15372 45106 15428 45108
rect 15372 45054 15374 45106
rect 15374 45054 15426 45106
rect 15426 45054 15428 45106
rect 15372 45052 15428 45054
rect 15484 44940 15540 44996
rect 15596 45052 15652 45108
rect 15036 44716 15092 44772
rect 14700 43650 14756 43652
rect 14700 43598 14702 43650
rect 14702 43598 14754 43650
rect 14754 43598 14756 43650
rect 14700 43596 14756 43598
rect 15148 42924 15204 42980
rect 15372 42924 15428 42980
rect 14252 42754 14308 42756
rect 14252 42702 14254 42754
rect 14254 42702 14306 42754
rect 14306 42702 14308 42754
rect 14252 42700 14308 42702
rect 14140 41804 14196 41860
rect 13580 40908 13636 40964
rect 13692 39900 13748 39956
rect 13804 39564 13860 39620
rect 13468 37996 13524 38052
rect 13692 37884 13748 37940
rect 13356 37548 13412 37604
rect 14140 41074 14196 41076
rect 14140 41022 14142 41074
rect 14142 41022 14194 41074
rect 14194 41022 14196 41074
rect 14140 41020 14196 41022
rect 14028 39788 14084 39844
rect 14028 39618 14084 39620
rect 14028 39566 14030 39618
rect 14030 39566 14082 39618
rect 14082 39566 14084 39618
rect 14028 39564 14084 39566
rect 14476 41244 14532 41300
rect 15036 42082 15092 42084
rect 15036 42030 15038 42082
rect 15038 42030 15090 42082
rect 15090 42030 15092 42082
rect 15036 42028 15092 42030
rect 15148 41916 15204 41972
rect 15260 42588 15316 42644
rect 15260 41356 15316 41412
rect 14252 40124 14308 40180
rect 14588 40402 14644 40404
rect 14588 40350 14590 40402
rect 14590 40350 14642 40402
rect 14642 40350 14644 40402
rect 14588 40348 14644 40350
rect 14476 39564 14532 39620
rect 14364 38834 14420 38836
rect 14364 38782 14366 38834
rect 14366 38782 14418 38834
rect 14418 38782 14420 38834
rect 14364 38780 14420 38782
rect 13916 37548 13972 37604
rect 13356 37324 13412 37380
rect 13916 37212 13972 37268
rect 14700 40124 14756 40180
rect 15036 41074 15092 41076
rect 15036 41022 15038 41074
rect 15038 41022 15090 41074
rect 15090 41022 15092 41074
rect 15036 41020 15092 41022
rect 15372 41244 15428 41300
rect 14924 40572 14980 40628
rect 14812 39506 14868 39508
rect 14812 39454 14814 39506
rect 14814 39454 14866 39506
rect 14866 39454 14868 39506
rect 14812 39452 14868 39454
rect 14700 39340 14756 39396
rect 14700 38722 14756 38724
rect 14700 38670 14702 38722
rect 14702 38670 14754 38722
rect 14754 38670 14756 38722
rect 14700 38668 14756 38670
rect 14588 37996 14644 38052
rect 14364 37212 14420 37268
rect 13580 36428 13636 36484
rect 12684 33628 12740 33684
rect 12796 33458 12852 33460
rect 12796 33406 12798 33458
rect 12798 33406 12850 33458
rect 12850 33406 12852 33458
rect 12796 33404 12852 33406
rect 12236 32172 12292 32228
rect 12348 33346 12404 33348
rect 12348 33294 12350 33346
rect 12350 33294 12402 33346
rect 12402 33294 12404 33346
rect 12348 33292 12404 33294
rect 12236 31836 12292 31892
rect 11676 31218 11732 31220
rect 11676 31166 11678 31218
rect 11678 31166 11730 31218
rect 11730 31166 11732 31218
rect 11676 31164 11732 31166
rect 10892 30828 10948 30884
rect 11228 30828 11284 30884
rect 10556 28754 10612 28756
rect 10556 28702 10558 28754
rect 10558 28702 10610 28754
rect 10610 28702 10612 28754
rect 10556 28700 10612 28702
rect 10332 28588 10388 28644
rect 10220 27356 10276 27412
rect 10220 27186 10276 27188
rect 10220 27134 10222 27186
rect 10222 27134 10274 27186
rect 10274 27134 10276 27186
rect 10220 27132 10276 27134
rect 10556 28082 10612 28084
rect 10556 28030 10558 28082
rect 10558 28030 10610 28082
rect 10610 28030 10612 28082
rect 10556 28028 10612 28030
rect 10892 27916 10948 27972
rect 11004 27020 11060 27076
rect 11564 30210 11620 30212
rect 11564 30158 11566 30210
rect 11566 30158 11618 30210
rect 11618 30158 11620 30210
rect 11564 30156 11620 30158
rect 11340 28028 11396 28084
rect 11564 28028 11620 28084
rect 11340 27804 11396 27860
rect 11676 27970 11732 27972
rect 11676 27918 11678 27970
rect 11678 27918 11730 27970
rect 11730 27918 11732 27970
rect 11676 27916 11732 27918
rect 10108 23996 10164 24052
rect 10444 26908 10500 26964
rect 9324 21756 9380 21812
rect 8316 18844 8372 18900
rect 8316 18338 8372 18340
rect 8316 18286 8318 18338
rect 8318 18286 8370 18338
rect 8370 18286 8372 18338
rect 8316 18284 8372 18286
rect 8204 18172 8260 18228
rect 7980 17724 8036 17780
rect 8316 17164 8372 17220
rect 8652 19404 8708 19460
rect 8428 16940 8484 16996
rect 7980 16044 8036 16100
rect 7420 15932 7476 15988
rect 7308 15372 7364 15428
rect 7084 15202 7140 15204
rect 7084 15150 7086 15202
rect 7086 15150 7138 15202
rect 7138 15150 7140 15202
rect 7084 15148 7140 15150
rect 6860 14530 6916 14532
rect 6860 14478 6862 14530
rect 6862 14478 6914 14530
rect 6914 14478 6916 14530
rect 6860 14476 6916 14478
rect 6188 13916 6244 13972
rect 6300 13356 6356 13412
rect 5740 12738 5796 12740
rect 5740 12686 5742 12738
rect 5742 12686 5794 12738
rect 5794 12686 5796 12738
rect 5740 12684 5796 12686
rect 5964 12124 6020 12180
rect 5628 11900 5684 11956
rect 5740 11228 5796 11284
rect 5852 10668 5908 10724
rect 5964 10892 6020 10948
rect 6076 11116 6132 11172
rect 6636 12796 6692 12852
rect 6860 13244 6916 13300
rect 6524 12012 6580 12068
rect 6524 11394 6580 11396
rect 6524 11342 6526 11394
rect 6526 11342 6578 11394
rect 6578 11342 6580 11394
rect 6524 11340 6580 11342
rect 7196 13970 7252 13972
rect 7196 13918 7198 13970
rect 7198 13918 7250 13970
rect 7250 13918 7252 13970
rect 7196 13916 7252 13918
rect 9772 23378 9828 23380
rect 9772 23326 9774 23378
rect 9774 23326 9826 23378
rect 9826 23326 9828 23378
rect 9772 23324 9828 23326
rect 9772 22988 9828 23044
rect 9660 22204 9716 22260
rect 9548 20802 9604 20804
rect 9548 20750 9550 20802
rect 9550 20750 9602 20802
rect 9602 20750 9604 20802
rect 9548 20748 9604 20750
rect 9436 20690 9492 20692
rect 9436 20638 9438 20690
rect 9438 20638 9490 20690
rect 9490 20638 9492 20690
rect 9436 20636 9492 20638
rect 9884 21474 9940 21476
rect 9884 21422 9886 21474
rect 9886 21422 9938 21474
rect 9938 21422 9940 21474
rect 9884 21420 9940 21422
rect 10332 25788 10388 25844
rect 10332 24610 10388 24612
rect 10332 24558 10334 24610
rect 10334 24558 10386 24610
rect 10386 24558 10388 24610
rect 10332 24556 10388 24558
rect 10220 23436 10276 23492
rect 10108 20636 10164 20692
rect 9436 19180 9492 19236
rect 9772 20018 9828 20020
rect 9772 19966 9774 20018
rect 9774 19966 9826 20018
rect 9826 19966 9828 20018
rect 9772 19964 9828 19966
rect 9884 19516 9940 19572
rect 9996 19964 10052 20020
rect 9548 18172 9604 18228
rect 9884 19234 9940 19236
rect 9884 19182 9886 19234
rect 9886 19182 9938 19234
rect 9938 19182 9940 19234
rect 9884 19180 9940 19182
rect 10668 26908 10724 26964
rect 10780 25394 10836 25396
rect 10780 25342 10782 25394
rect 10782 25342 10834 25394
rect 10834 25342 10836 25394
rect 10780 25340 10836 25342
rect 11004 25282 11060 25284
rect 11004 25230 11006 25282
rect 11006 25230 11058 25282
rect 11058 25230 11060 25282
rect 11004 25228 11060 25230
rect 10892 24220 10948 24276
rect 11452 26796 11508 26852
rect 12124 31164 12180 31220
rect 12572 32450 12628 32452
rect 12572 32398 12574 32450
rect 12574 32398 12626 32450
rect 12626 32398 12628 32450
rect 12572 32396 12628 32398
rect 14028 36988 14084 37044
rect 13916 36204 13972 36260
rect 14140 36540 14196 36596
rect 13804 34636 13860 34692
rect 13132 33516 13188 33572
rect 13244 33906 13300 33908
rect 13244 33854 13246 33906
rect 13246 33854 13298 33906
rect 13298 33854 13300 33906
rect 13244 33852 13300 33854
rect 13132 32284 13188 32340
rect 13020 31948 13076 32004
rect 12684 31836 12740 31892
rect 12684 31388 12740 31444
rect 12796 31218 12852 31220
rect 12796 31166 12798 31218
rect 12798 31166 12850 31218
rect 12850 31166 12852 31218
rect 12796 31164 12852 31166
rect 13356 32396 13412 32452
rect 13468 31164 13524 31220
rect 12460 30994 12516 30996
rect 12460 30942 12462 30994
rect 12462 30942 12514 30994
rect 12514 30942 12516 30994
rect 12460 30940 12516 30942
rect 12908 30156 12964 30212
rect 13132 30940 13188 30996
rect 12236 27916 12292 27972
rect 13020 29036 13076 29092
rect 13132 28700 13188 28756
rect 12796 28642 12852 28644
rect 12796 28590 12798 28642
rect 12798 28590 12850 28642
rect 12850 28590 12852 28642
rect 12796 28588 12852 28590
rect 12460 28028 12516 28084
rect 12348 27804 12404 27860
rect 11900 26962 11956 26964
rect 11900 26910 11902 26962
rect 11902 26910 11954 26962
rect 11954 26910 11956 26962
rect 11900 26908 11956 26910
rect 11788 26796 11844 26852
rect 11788 26572 11844 26628
rect 12460 26572 12516 26628
rect 12572 26796 12628 26852
rect 12236 26514 12292 26516
rect 12236 26462 12238 26514
rect 12238 26462 12290 26514
rect 12290 26462 12292 26514
rect 12236 26460 12292 26462
rect 13468 28588 13524 28644
rect 13356 27970 13412 27972
rect 13356 27918 13358 27970
rect 13358 27918 13410 27970
rect 13410 27918 13412 27970
rect 13356 27916 13412 27918
rect 13244 26796 13300 26852
rect 12908 26684 12964 26740
rect 12684 26236 12740 26292
rect 12012 25676 12068 25732
rect 12012 25228 12068 25284
rect 11788 24556 11844 24612
rect 11900 24444 11956 24500
rect 10780 22540 10836 22596
rect 10892 22258 10948 22260
rect 10892 22206 10894 22258
rect 10894 22206 10946 22258
rect 10946 22206 10948 22258
rect 10892 22204 10948 22206
rect 11004 22988 11060 23044
rect 11004 21868 11060 21924
rect 11228 22428 11284 22484
rect 11788 23548 11844 23604
rect 11900 23436 11956 23492
rect 11788 22540 11844 22596
rect 12572 25452 12628 25508
rect 12460 25282 12516 25284
rect 12460 25230 12462 25282
rect 12462 25230 12514 25282
rect 12514 25230 12516 25282
rect 12460 25228 12516 25230
rect 12348 24780 12404 24836
rect 12236 24162 12292 24164
rect 12236 24110 12238 24162
rect 12238 24110 12290 24162
rect 12290 24110 12292 24162
rect 12236 24108 12292 24110
rect 12796 26178 12852 26180
rect 12796 26126 12798 26178
rect 12798 26126 12850 26178
rect 12850 26126 12852 26178
rect 12796 26124 12852 26126
rect 13020 25452 13076 25508
rect 13132 25340 13188 25396
rect 12908 25004 12964 25060
rect 12684 24892 12740 24948
rect 13132 24892 13188 24948
rect 13468 26012 13524 26068
rect 14028 34300 14084 34356
rect 14700 37772 14756 37828
rect 14700 36652 14756 36708
rect 13804 32956 13860 33012
rect 14252 33122 14308 33124
rect 14252 33070 14254 33122
rect 14254 33070 14306 33122
rect 14306 33070 14308 33122
rect 14252 33068 14308 33070
rect 15036 39564 15092 39620
rect 15260 39618 15316 39620
rect 15260 39566 15262 39618
rect 15262 39566 15314 39618
rect 15314 39566 15316 39618
rect 15260 39564 15316 39566
rect 15260 38220 15316 38276
rect 15148 37884 15204 37940
rect 15148 36988 15204 37044
rect 14924 36204 14980 36260
rect 15148 36652 15204 36708
rect 15932 48188 15988 48244
rect 15820 48076 15876 48132
rect 16156 48524 16212 48580
rect 16604 50316 16660 50372
rect 16380 49922 16436 49924
rect 16380 49870 16382 49922
rect 16382 49870 16434 49922
rect 16434 49870 16436 49922
rect 16380 49868 16436 49870
rect 16268 47740 16324 47796
rect 16380 49644 16436 49700
rect 16268 47346 16324 47348
rect 16268 47294 16270 47346
rect 16270 47294 16322 47346
rect 16322 47294 16324 47346
rect 16268 47292 16324 47294
rect 16716 50034 16772 50036
rect 16716 49982 16718 50034
rect 16718 49982 16770 50034
rect 16770 49982 16772 50034
rect 16716 49980 16772 49982
rect 16828 49308 16884 49364
rect 17164 51660 17220 51716
rect 17276 51548 17332 51604
rect 17388 51884 17444 51940
rect 17612 52332 17668 52388
rect 17612 51996 17668 52052
rect 17948 55468 18004 55524
rect 17948 54514 18004 54516
rect 17948 54462 17950 54514
rect 17950 54462 18002 54514
rect 18002 54462 18004 54514
rect 17948 54460 18004 54462
rect 17836 54402 17892 54404
rect 17836 54350 17838 54402
rect 17838 54350 17890 54402
rect 17890 54350 17892 54402
rect 17836 54348 17892 54350
rect 17836 54124 17892 54180
rect 18284 56642 18340 56644
rect 18284 56590 18286 56642
rect 18286 56590 18338 56642
rect 18338 56590 18340 56642
rect 18284 56588 18340 56590
rect 18284 55468 18340 55524
rect 18508 56866 18564 56868
rect 18508 56814 18510 56866
rect 18510 56814 18562 56866
rect 18562 56814 18564 56866
rect 18508 56812 18564 56814
rect 19292 57538 19348 57540
rect 19292 57486 19294 57538
rect 19294 57486 19346 57538
rect 19346 57486 19348 57538
rect 19292 57484 19348 57486
rect 19404 57260 19460 57316
rect 19180 56700 19236 56756
rect 18956 56252 19012 56308
rect 18508 56082 18564 56084
rect 18508 56030 18510 56082
rect 18510 56030 18562 56082
rect 18562 56030 18564 56082
rect 18508 56028 18564 56030
rect 18060 53452 18116 53508
rect 18172 55020 18228 55076
rect 18732 55244 18788 55300
rect 18284 54796 18340 54852
rect 18620 55132 18676 55188
rect 18060 53228 18116 53284
rect 17836 53058 17892 53060
rect 17836 53006 17838 53058
rect 17838 53006 17890 53058
rect 17890 53006 17892 53058
rect 17836 53004 17892 53006
rect 17612 49868 17668 49924
rect 17388 49308 17444 49364
rect 16604 48972 16660 49028
rect 16492 48300 16548 48356
rect 16604 48748 16660 48804
rect 16604 47740 16660 47796
rect 16156 46956 16212 47012
rect 15932 46786 15988 46788
rect 15932 46734 15934 46786
rect 15934 46734 15986 46786
rect 15986 46734 15988 46786
rect 15932 46732 15988 46734
rect 16156 46674 16212 46676
rect 16156 46622 16158 46674
rect 16158 46622 16210 46674
rect 16210 46622 16212 46674
rect 16156 46620 16212 46622
rect 16268 46562 16324 46564
rect 16268 46510 16270 46562
rect 16270 46510 16322 46562
rect 16322 46510 16324 46562
rect 16268 46508 16324 46510
rect 16268 44492 16324 44548
rect 17276 46732 17332 46788
rect 16716 46284 16772 46340
rect 16828 46060 16884 46116
rect 16380 44268 16436 44324
rect 17612 49026 17668 49028
rect 17612 48974 17614 49026
rect 17614 48974 17666 49026
rect 17666 48974 17668 49026
rect 17612 48972 17668 48974
rect 18508 54684 18564 54740
rect 18620 54514 18676 54516
rect 18620 54462 18622 54514
rect 18622 54462 18674 54514
rect 18674 54462 18676 54514
rect 18620 54460 18676 54462
rect 18508 54124 18564 54180
rect 18508 53340 18564 53396
rect 19180 54684 19236 54740
rect 18844 53676 18900 53732
rect 20076 58492 20132 58548
rect 19628 58434 19684 58436
rect 19628 58382 19630 58434
rect 19630 58382 19682 58434
rect 19682 58382 19684 58434
rect 19628 58380 19684 58382
rect 19628 58044 19684 58100
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19740 57708 19796 57764
rect 19964 57820 20020 57876
rect 19628 57484 19684 57540
rect 20188 56812 20244 56868
rect 19740 56754 19796 56756
rect 19740 56702 19742 56754
rect 19742 56702 19794 56754
rect 19794 56702 19796 56754
rect 19740 56700 19796 56702
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 20188 56364 20244 56420
rect 20188 56140 20244 56196
rect 19516 55356 19572 55412
rect 19740 55132 19796 55188
rect 20188 55468 20244 55524
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19516 54572 19572 54628
rect 19852 54402 19908 54404
rect 19852 54350 19854 54402
rect 19854 54350 19906 54402
rect 19906 54350 19908 54402
rect 19852 54348 19908 54350
rect 19404 53564 19460 53620
rect 19516 54236 19572 54292
rect 19068 52668 19124 52724
rect 19180 53452 19236 53508
rect 18172 52332 18228 52388
rect 18844 51772 18900 51828
rect 18396 51660 18452 51716
rect 18060 49644 18116 49700
rect 18284 49308 18340 49364
rect 18844 51436 18900 51492
rect 18956 49868 19012 49924
rect 18396 49084 18452 49140
rect 18508 49532 18564 49588
rect 18284 48972 18340 49028
rect 18060 48242 18116 48244
rect 18060 48190 18062 48242
rect 18062 48190 18114 48242
rect 18114 48190 18116 48242
rect 18060 48188 18116 48190
rect 18060 47516 18116 47572
rect 18508 48748 18564 48804
rect 18508 48300 18564 48356
rect 18172 47404 18228 47460
rect 18284 47964 18340 48020
rect 17948 46956 18004 47012
rect 17724 46786 17780 46788
rect 17724 46734 17726 46786
rect 17726 46734 17778 46786
rect 17778 46734 17780 46786
rect 17724 46732 17780 46734
rect 17388 46620 17444 46676
rect 17724 46508 17780 46564
rect 17276 45724 17332 45780
rect 17612 45948 17668 46004
rect 17388 45500 17444 45556
rect 16716 44882 16772 44884
rect 16716 44830 16718 44882
rect 16718 44830 16770 44882
rect 16770 44830 16772 44882
rect 16716 44828 16772 44830
rect 16156 43650 16212 43652
rect 16156 43598 16158 43650
rect 16158 43598 16210 43650
rect 16210 43598 16212 43650
rect 16156 43596 16212 43598
rect 17388 44268 17444 44324
rect 17724 45836 17780 45892
rect 17612 45724 17668 45780
rect 16268 42140 16324 42196
rect 16044 41804 16100 41860
rect 15708 41244 15764 41300
rect 15484 40908 15540 40964
rect 15484 40236 15540 40292
rect 15820 39564 15876 39620
rect 15932 39452 15988 39508
rect 16044 40908 16100 40964
rect 16268 40962 16324 40964
rect 16268 40910 16270 40962
rect 16270 40910 16322 40962
rect 16322 40910 16324 40962
rect 16268 40908 16324 40910
rect 16604 40908 16660 40964
rect 17164 41804 17220 41860
rect 16940 41692 16996 41748
rect 16940 41186 16996 41188
rect 16940 41134 16942 41186
rect 16942 41134 16994 41186
rect 16994 41134 16996 41186
rect 16940 41132 16996 41134
rect 17500 41970 17556 41972
rect 17500 41918 17502 41970
rect 17502 41918 17554 41970
rect 17554 41918 17556 41970
rect 17500 41916 17556 41918
rect 17612 41132 17668 41188
rect 16828 40124 16884 40180
rect 16828 39842 16884 39844
rect 16828 39790 16830 39842
rect 16830 39790 16882 39842
rect 16882 39790 16884 39842
rect 16828 39788 16884 39790
rect 16604 39506 16660 39508
rect 16604 39454 16606 39506
rect 16606 39454 16658 39506
rect 16658 39454 16660 39506
rect 16604 39452 16660 39454
rect 16492 39116 16548 39172
rect 16156 38780 16212 38836
rect 15596 38220 15652 38276
rect 15596 38050 15652 38052
rect 15596 37998 15598 38050
rect 15598 37998 15650 38050
rect 15650 37998 15652 38050
rect 15596 37996 15652 37998
rect 15708 37884 15764 37940
rect 15932 37996 15988 38052
rect 16940 39564 16996 39620
rect 16268 38220 16324 38276
rect 16044 37212 16100 37268
rect 15372 36540 15428 36596
rect 15260 35532 15316 35588
rect 15372 35196 15428 35252
rect 14812 34636 14868 34692
rect 15372 34412 15428 34468
rect 16044 36370 16100 36372
rect 16044 36318 16046 36370
rect 16046 36318 16098 36370
rect 16098 36318 16100 36370
rect 16044 36316 16100 36318
rect 17164 38892 17220 38948
rect 17276 39116 17332 39172
rect 17612 39506 17668 39508
rect 17612 39454 17614 39506
rect 17614 39454 17666 39506
rect 17666 39454 17668 39506
rect 17612 39452 17668 39454
rect 17612 39228 17668 39284
rect 17164 36540 17220 36596
rect 16268 36204 16324 36260
rect 16828 35868 16884 35924
rect 17500 37266 17556 37268
rect 17500 37214 17502 37266
rect 17502 37214 17554 37266
rect 17554 37214 17556 37266
rect 17500 37212 17556 37214
rect 17500 36594 17556 36596
rect 17500 36542 17502 36594
rect 17502 36542 17554 36594
rect 17554 36542 17556 36594
rect 17500 36540 17556 36542
rect 17724 38946 17780 38948
rect 17724 38894 17726 38946
rect 17726 38894 17778 38946
rect 17778 38894 17780 38946
rect 17724 38892 17780 38894
rect 19292 53116 19348 53172
rect 19852 54124 19908 54180
rect 20076 53564 20132 53620
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 22540 59836 22596 59892
rect 20860 59164 20916 59220
rect 20972 58828 21028 58884
rect 22092 59612 22148 59668
rect 21756 59052 21812 59108
rect 21420 58940 21476 58996
rect 20524 57260 20580 57316
rect 20748 57484 20804 57540
rect 20524 56140 20580 56196
rect 20636 57036 20692 57092
rect 20972 57036 21028 57092
rect 21196 57708 21252 57764
rect 21980 58546 22036 58548
rect 21980 58494 21982 58546
rect 21982 58494 22034 58546
rect 22034 58494 22036 58546
rect 21980 58492 22036 58494
rect 23212 59890 23268 59892
rect 23212 59838 23214 59890
rect 23214 59838 23266 59890
rect 23266 59838 23268 59890
rect 23212 59836 23268 59838
rect 23436 58994 23492 58996
rect 23436 58942 23438 58994
rect 23438 58942 23490 58994
rect 23490 58942 23492 58994
rect 23436 58940 23492 58942
rect 21532 58044 21588 58100
rect 21868 57650 21924 57652
rect 21868 57598 21870 57650
rect 21870 57598 21922 57650
rect 21922 57598 21924 57650
rect 21868 57596 21924 57598
rect 21644 56812 21700 56868
rect 22092 57650 22148 57652
rect 22092 57598 22094 57650
rect 22094 57598 22146 57650
rect 22146 57598 22148 57650
rect 22092 57596 22148 57598
rect 22092 57148 22148 57204
rect 23212 57426 23268 57428
rect 23212 57374 23214 57426
rect 23214 57374 23266 57426
rect 23266 57374 23268 57426
rect 23212 57372 23268 57374
rect 23660 59164 23716 59220
rect 24556 59218 24612 59220
rect 24556 59166 24558 59218
rect 24558 59166 24610 59218
rect 24610 59166 24612 59218
rect 24556 59164 24612 59166
rect 23884 58828 23940 58884
rect 23884 58492 23940 58548
rect 23548 56924 23604 56980
rect 22764 56588 22820 56644
rect 21196 56306 21252 56308
rect 21196 56254 21198 56306
rect 21198 56254 21250 56306
rect 21250 56254 21252 56306
rect 21196 56252 21252 56254
rect 21868 55244 21924 55300
rect 20860 55132 20916 55188
rect 21980 55074 22036 55076
rect 21980 55022 21982 55074
rect 21982 55022 22034 55074
rect 22034 55022 22036 55074
rect 21980 55020 22036 55022
rect 22092 54908 22148 54964
rect 22652 55580 22708 55636
rect 22204 54684 22260 54740
rect 20972 54626 21028 54628
rect 20972 54574 20974 54626
rect 20974 54574 21026 54626
rect 21026 54574 21028 54626
rect 20972 54572 21028 54574
rect 20636 54124 20692 54180
rect 20748 54460 20804 54516
rect 21532 54460 21588 54516
rect 21308 53788 21364 53844
rect 21532 53730 21588 53732
rect 21532 53678 21534 53730
rect 21534 53678 21586 53730
rect 21586 53678 21588 53730
rect 21532 53676 21588 53678
rect 20300 53452 20356 53508
rect 19964 53004 20020 53060
rect 19740 52780 19796 52836
rect 20524 52834 20580 52836
rect 20524 52782 20526 52834
rect 20526 52782 20578 52834
rect 20578 52782 20580 52834
rect 20524 52780 20580 52782
rect 20636 52556 20692 52612
rect 20524 52220 20580 52276
rect 20412 51996 20468 52052
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 20076 51602 20132 51604
rect 20076 51550 20078 51602
rect 20078 51550 20130 51602
rect 20130 51550 20132 51602
rect 20076 51548 20132 51550
rect 19516 51212 19572 51268
rect 20524 50594 20580 50596
rect 20524 50542 20526 50594
rect 20526 50542 20578 50594
rect 20578 50542 20580 50594
rect 20524 50540 20580 50542
rect 20636 50482 20692 50484
rect 20636 50430 20638 50482
rect 20638 50430 20690 50482
rect 20690 50430 20692 50482
rect 20636 50428 20692 50430
rect 19516 49810 19572 49812
rect 19516 49758 19518 49810
rect 19518 49758 19570 49810
rect 19570 49758 19572 49810
rect 19516 49756 19572 49758
rect 20300 50370 20356 50372
rect 20300 50318 20302 50370
rect 20302 50318 20354 50370
rect 20354 50318 20356 50370
rect 20300 50316 20356 50318
rect 20748 50316 20804 50372
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 20300 50092 20356 50148
rect 20076 49756 20132 49812
rect 19180 48188 19236 48244
rect 19964 49586 20020 49588
rect 19964 49534 19966 49586
rect 19966 49534 20018 49586
rect 20018 49534 20020 49586
rect 19964 49532 20020 49534
rect 19292 47740 19348 47796
rect 18508 46844 18564 46900
rect 18620 47628 18676 47684
rect 18284 46562 18340 46564
rect 18284 46510 18286 46562
rect 18286 46510 18338 46562
rect 18338 46510 18340 46562
rect 18284 46508 18340 46510
rect 18172 46114 18228 46116
rect 18172 46062 18174 46114
rect 18174 46062 18226 46114
rect 18226 46062 18228 46114
rect 18172 46060 18228 46062
rect 18844 46060 18900 46116
rect 18956 46002 19012 46004
rect 18956 45950 18958 46002
rect 18958 45950 19010 46002
rect 19010 45950 19012 46002
rect 18956 45948 19012 45950
rect 18620 45890 18676 45892
rect 18620 45838 18622 45890
rect 18622 45838 18674 45890
rect 18674 45838 18676 45890
rect 18620 45836 18676 45838
rect 18060 45612 18116 45668
rect 17948 43426 18004 43428
rect 17948 43374 17950 43426
rect 17950 43374 18002 43426
rect 18002 43374 18004 43426
rect 17948 43372 18004 43374
rect 18060 45106 18116 45108
rect 18060 45054 18062 45106
rect 18062 45054 18114 45106
rect 18114 45054 18116 45106
rect 18060 45052 18116 45054
rect 18620 44604 18676 44660
rect 18508 43484 18564 43540
rect 17948 42700 18004 42756
rect 18396 43260 18452 43316
rect 18732 43484 18788 43540
rect 18508 43036 18564 43092
rect 17948 42140 18004 42196
rect 17948 41804 18004 41860
rect 17948 40460 18004 40516
rect 18172 42028 18228 42084
rect 18396 42194 18452 42196
rect 18396 42142 18398 42194
rect 18398 42142 18450 42194
rect 18450 42142 18452 42194
rect 18396 42140 18452 42142
rect 19740 49420 19796 49476
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 20524 48242 20580 48244
rect 20524 48190 20526 48242
rect 20526 48190 20578 48242
rect 20578 48190 20580 48242
rect 20524 48188 20580 48190
rect 19852 47628 19908 47684
rect 19964 47740 20020 47796
rect 20524 47740 20580 47796
rect 20300 47458 20356 47460
rect 20300 47406 20302 47458
rect 20302 47406 20354 47458
rect 20354 47406 20356 47458
rect 20300 47404 20356 47406
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19740 46844 19796 46900
rect 20188 46844 20244 46900
rect 20076 46002 20132 46004
rect 20076 45950 20078 46002
rect 20078 45950 20130 46002
rect 20130 45950 20132 46002
rect 20076 45948 20132 45950
rect 19740 45724 19796 45780
rect 20076 45612 20132 45668
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 20188 45106 20244 45108
rect 20188 45054 20190 45106
rect 20190 45054 20242 45106
rect 20242 45054 20244 45106
rect 20188 45052 20244 45054
rect 21756 53228 21812 53284
rect 21756 53004 21812 53060
rect 21308 52892 21364 52948
rect 21420 52722 21476 52724
rect 21420 52670 21422 52722
rect 21422 52670 21474 52722
rect 21474 52670 21476 52722
rect 21420 52668 21476 52670
rect 21532 52556 21588 52612
rect 21756 52780 21812 52836
rect 21420 51772 21476 51828
rect 21532 51490 21588 51492
rect 21532 51438 21534 51490
rect 21534 51438 21586 51490
rect 21586 51438 21588 51490
rect 21532 51436 21588 51438
rect 21196 51212 21252 51268
rect 21084 47852 21140 47908
rect 20860 45836 20916 45892
rect 20860 45666 20916 45668
rect 20860 45614 20862 45666
rect 20862 45614 20914 45666
rect 20914 45614 20916 45666
rect 20860 45612 20916 45614
rect 20524 45276 20580 45332
rect 20524 44322 20580 44324
rect 20524 44270 20526 44322
rect 20526 44270 20578 44322
rect 20578 44270 20580 44322
rect 20524 44268 20580 44270
rect 20636 45106 20692 45108
rect 20636 45054 20638 45106
rect 20638 45054 20690 45106
rect 20690 45054 20692 45106
rect 20636 45052 20692 45054
rect 19516 44044 19572 44100
rect 20524 44044 20580 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20300 43820 20356 43876
rect 19068 43596 19124 43652
rect 19852 43596 19908 43652
rect 19516 43538 19572 43540
rect 19516 43486 19518 43538
rect 19518 43486 19570 43538
rect 19570 43486 19572 43538
rect 19516 43484 19572 43486
rect 19292 43260 19348 43316
rect 20300 43484 20356 43540
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 18396 40962 18452 40964
rect 18396 40910 18398 40962
rect 18398 40910 18450 40962
rect 18450 40910 18452 40962
rect 18396 40908 18452 40910
rect 18172 40348 18228 40404
rect 18060 40124 18116 40180
rect 18396 39618 18452 39620
rect 18396 39566 18398 39618
rect 18398 39566 18450 39618
rect 18450 39566 18452 39618
rect 18396 39564 18452 39566
rect 18844 40962 18900 40964
rect 18844 40910 18846 40962
rect 18846 40910 18898 40962
rect 18898 40910 18900 40962
rect 18844 40908 18900 40910
rect 17948 39506 18004 39508
rect 17948 39454 17950 39506
rect 17950 39454 18002 39506
rect 18002 39454 18004 39506
rect 17948 39452 18004 39454
rect 18508 39394 18564 39396
rect 18508 39342 18510 39394
rect 18510 39342 18562 39394
rect 18562 39342 18564 39394
rect 18508 39340 18564 39342
rect 17948 39116 18004 39172
rect 18508 37938 18564 37940
rect 18508 37886 18510 37938
rect 18510 37886 18562 37938
rect 18562 37886 18564 37938
rect 18508 37884 18564 37886
rect 17948 37266 18004 37268
rect 17948 37214 17950 37266
rect 17950 37214 18002 37266
rect 18002 37214 18004 37266
rect 17948 37212 18004 37214
rect 18620 36764 18676 36820
rect 17612 36092 17668 36148
rect 15596 35644 15652 35700
rect 17052 35420 17108 35476
rect 15036 34076 15092 34132
rect 14700 33068 14756 33124
rect 14588 32956 14644 33012
rect 14924 32844 14980 32900
rect 14028 32060 14084 32116
rect 13804 31164 13860 31220
rect 13692 31052 13748 31108
rect 13692 30380 13748 30436
rect 14028 30940 14084 30996
rect 13804 29372 13860 29428
rect 14028 30604 14084 30660
rect 14140 30380 14196 30436
rect 14924 32508 14980 32564
rect 14364 31778 14420 31780
rect 14364 31726 14366 31778
rect 14366 31726 14418 31778
rect 14418 31726 14420 31778
rect 14364 31724 14420 31726
rect 14476 31052 14532 31108
rect 15260 31836 15316 31892
rect 14588 31724 14644 31780
rect 14700 31612 14756 31668
rect 15148 31612 15204 31668
rect 15036 31388 15092 31444
rect 14812 31106 14868 31108
rect 14812 31054 14814 31106
rect 14814 31054 14866 31106
rect 14866 31054 14868 31106
rect 14812 31052 14868 31054
rect 14252 29372 14308 29428
rect 14140 28924 14196 28980
rect 13804 27858 13860 27860
rect 13804 27806 13806 27858
rect 13806 27806 13858 27858
rect 13858 27806 13860 27858
rect 13804 27804 13860 27806
rect 14476 29202 14532 29204
rect 14476 29150 14478 29202
rect 14478 29150 14530 29202
rect 14530 29150 14532 29202
rect 14476 29148 14532 29150
rect 14364 29036 14420 29092
rect 14700 28754 14756 28756
rect 14700 28702 14702 28754
rect 14702 28702 14754 28754
rect 14754 28702 14756 28754
rect 14700 28700 14756 28702
rect 14364 28642 14420 28644
rect 14364 28590 14366 28642
rect 14366 28590 14418 28642
rect 14418 28590 14420 28642
rect 14364 28588 14420 28590
rect 14028 27020 14084 27076
rect 15820 34130 15876 34132
rect 15820 34078 15822 34130
rect 15822 34078 15874 34130
rect 15874 34078 15876 34130
rect 15820 34076 15876 34078
rect 15708 33292 15764 33348
rect 16044 34914 16100 34916
rect 16044 34862 16046 34914
rect 16046 34862 16098 34914
rect 16098 34862 16100 34914
rect 16044 34860 16100 34862
rect 16828 34690 16884 34692
rect 16828 34638 16830 34690
rect 16830 34638 16882 34690
rect 16882 34638 16884 34690
rect 16828 34636 16884 34638
rect 16044 33852 16100 33908
rect 16044 33346 16100 33348
rect 16044 33294 16046 33346
rect 16046 33294 16098 33346
rect 16098 33294 16100 33346
rect 16044 33292 16100 33294
rect 15932 33068 15988 33124
rect 16828 33740 16884 33796
rect 16940 33404 16996 33460
rect 16380 33292 16436 33348
rect 15484 32396 15540 32452
rect 15596 31836 15652 31892
rect 16044 32562 16100 32564
rect 16044 32510 16046 32562
rect 16046 32510 16098 32562
rect 16098 32510 16100 32562
rect 16044 32508 16100 32510
rect 16268 32508 16324 32564
rect 15372 31164 15428 31220
rect 15708 31106 15764 31108
rect 15708 31054 15710 31106
rect 15710 31054 15762 31106
rect 15762 31054 15764 31106
rect 15708 31052 15764 31054
rect 16044 30940 16100 30996
rect 14588 27804 14644 27860
rect 15260 29426 15316 29428
rect 15260 29374 15262 29426
rect 15262 29374 15314 29426
rect 15314 29374 15316 29426
rect 15260 29372 15316 29374
rect 14700 27692 14756 27748
rect 15260 28924 15316 28980
rect 13580 25228 13636 25284
rect 14588 26514 14644 26516
rect 14588 26462 14590 26514
rect 14590 26462 14642 26514
rect 14642 26462 14644 26514
rect 14588 26460 14644 26462
rect 13804 26236 13860 26292
rect 13356 24892 13412 24948
rect 13580 25004 13636 25060
rect 13468 24780 13524 24836
rect 13356 24722 13412 24724
rect 13356 24670 13358 24722
rect 13358 24670 13410 24722
rect 13410 24670 13412 24722
rect 13356 24668 13412 24670
rect 13692 24892 13748 24948
rect 14924 27858 14980 27860
rect 14924 27806 14926 27858
rect 14926 27806 14978 27858
rect 14978 27806 14980 27858
rect 14924 27804 14980 27806
rect 15148 27244 15204 27300
rect 15036 26908 15092 26964
rect 14812 26290 14868 26292
rect 14812 26238 14814 26290
rect 14814 26238 14866 26290
rect 14866 26238 14868 26290
rect 14812 26236 14868 26238
rect 14476 25228 14532 25284
rect 14252 24780 14308 24836
rect 13692 24162 13748 24164
rect 13692 24110 13694 24162
rect 13694 24110 13746 24162
rect 13746 24110 13748 24162
rect 13692 24108 13748 24110
rect 13580 23436 13636 23492
rect 13468 22930 13524 22932
rect 13468 22878 13470 22930
rect 13470 22878 13522 22930
rect 13522 22878 13524 22930
rect 13468 22876 13524 22878
rect 12012 22540 12068 22596
rect 11564 22316 11620 22372
rect 11676 22204 11732 22260
rect 11116 21756 11172 21812
rect 10556 21362 10612 21364
rect 10556 21310 10558 21362
rect 10558 21310 10610 21362
rect 10610 21310 10612 21362
rect 10556 21308 10612 21310
rect 10220 19180 10276 19236
rect 10332 20524 10388 20580
rect 11116 21586 11172 21588
rect 11116 21534 11118 21586
rect 11118 21534 11170 21586
rect 11170 21534 11172 21586
rect 11116 21532 11172 21534
rect 10780 21474 10836 21476
rect 10780 21422 10782 21474
rect 10782 21422 10834 21474
rect 10834 21422 10836 21474
rect 10780 21420 10836 21422
rect 10556 19068 10612 19124
rect 9772 18338 9828 18340
rect 9772 18286 9774 18338
rect 9774 18286 9826 18338
rect 9826 18286 9828 18338
rect 9772 18284 9828 18286
rect 9884 17666 9940 17668
rect 9884 17614 9886 17666
rect 9886 17614 9938 17666
rect 9938 17614 9940 17666
rect 9884 17612 9940 17614
rect 9436 17388 9492 17444
rect 8988 17164 9044 17220
rect 8652 15708 8708 15764
rect 8764 16044 8820 16100
rect 7532 14476 7588 14532
rect 7084 13580 7140 13636
rect 7644 12796 7700 12852
rect 7084 12684 7140 12740
rect 7980 12684 8036 12740
rect 7308 11788 7364 11844
rect 6412 10780 6468 10836
rect 6636 11228 6692 11284
rect 6860 10610 6916 10612
rect 6860 10558 6862 10610
rect 6862 10558 6914 10610
rect 6914 10558 6916 10610
rect 6860 10556 6916 10558
rect 6636 10444 6692 10500
rect 7084 10444 7140 10500
rect 7756 11788 7812 11844
rect 7756 11116 7812 11172
rect 7756 10834 7812 10836
rect 7756 10782 7758 10834
rect 7758 10782 7810 10834
rect 7810 10782 7812 10834
rect 7756 10780 7812 10782
rect 7308 10108 7364 10164
rect 6748 9266 6804 9268
rect 6748 9214 6750 9266
rect 6750 9214 6802 9266
rect 6802 9214 6804 9266
rect 6748 9212 6804 9214
rect 7084 8930 7140 8932
rect 7084 8878 7086 8930
rect 7086 8878 7138 8930
rect 7138 8878 7140 8930
rect 7084 8876 7140 8878
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 9100 14364 9156 14420
rect 9324 15484 9380 15540
rect 9212 14306 9268 14308
rect 9212 14254 9214 14306
rect 9214 14254 9266 14306
rect 9266 14254 9268 14306
rect 9212 14252 9268 14254
rect 8988 13746 9044 13748
rect 8988 13694 8990 13746
rect 8990 13694 9042 13746
rect 9042 13694 9044 13746
rect 8988 13692 9044 13694
rect 8764 13468 8820 13524
rect 8540 13356 8596 13412
rect 8428 13244 8484 13300
rect 8652 13020 8708 13076
rect 8540 12796 8596 12852
rect 8988 12236 9044 12292
rect 8988 11900 9044 11956
rect 8204 11788 8260 11844
rect 8428 11676 8484 11732
rect 8204 11452 8260 11508
rect 7980 8540 8036 8596
rect 8316 10780 8372 10836
rect 8876 11340 8932 11396
rect 8540 10722 8596 10724
rect 8540 10670 8542 10722
rect 8542 10670 8594 10722
rect 8594 10670 8596 10722
rect 8540 10668 8596 10670
rect 8988 10610 9044 10612
rect 8988 10558 8990 10610
rect 8990 10558 9042 10610
rect 9042 10558 9044 10610
rect 8988 10556 9044 10558
rect 9884 17164 9940 17220
rect 9548 16940 9604 16996
rect 10332 18674 10388 18676
rect 10332 18622 10334 18674
rect 10334 18622 10386 18674
rect 10386 18622 10388 18674
rect 10332 18620 10388 18622
rect 10220 18172 10276 18228
rect 10108 17052 10164 17108
rect 10108 16716 10164 16772
rect 10332 16716 10388 16772
rect 10668 17164 10724 17220
rect 11228 19404 11284 19460
rect 10780 17276 10836 17332
rect 12348 22258 12404 22260
rect 12348 22206 12350 22258
rect 12350 22206 12402 22258
rect 12402 22206 12404 22258
rect 12348 22204 12404 22206
rect 12012 22146 12068 22148
rect 12012 22094 12014 22146
rect 12014 22094 12066 22146
rect 12066 22094 12068 22146
rect 12012 22092 12068 22094
rect 12572 22146 12628 22148
rect 12572 22094 12574 22146
rect 12574 22094 12626 22146
rect 12626 22094 12628 22146
rect 12572 22092 12628 22094
rect 12012 21756 12068 21812
rect 12684 21644 12740 21700
rect 12572 21474 12628 21476
rect 12572 21422 12574 21474
rect 12574 21422 12626 21474
rect 12626 21422 12628 21474
rect 12572 21420 12628 21422
rect 12012 21308 12068 21364
rect 12460 21308 12516 21364
rect 11900 20860 11956 20916
rect 12572 20860 12628 20916
rect 11900 20188 11956 20244
rect 11788 20130 11844 20132
rect 11788 20078 11790 20130
rect 11790 20078 11842 20130
rect 11842 20078 11844 20130
rect 11788 20076 11844 20078
rect 11788 19234 11844 19236
rect 11788 19182 11790 19234
rect 11790 19182 11842 19234
rect 11842 19182 11844 19234
rect 11788 19180 11844 19182
rect 11004 17836 11060 17892
rect 10444 16268 10500 16324
rect 11340 18396 11396 18452
rect 11340 17948 11396 18004
rect 11004 16828 11060 16884
rect 9996 16044 10052 16100
rect 9324 11676 9380 11732
rect 9436 13580 9492 13636
rect 9884 14418 9940 14420
rect 9884 14366 9886 14418
rect 9886 14366 9938 14418
rect 9938 14366 9940 14418
rect 9884 14364 9940 14366
rect 9660 14252 9716 14308
rect 9548 13356 9604 13412
rect 9884 12796 9940 12852
rect 9996 13020 10052 13076
rect 8316 9548 8372 9604
rect 8540 8540 8596 8596
rect 8876 9154 8932 9156
rect 8876 9102 8878 9154
rect 8878 9102 8930 9154
rect 8930 9102 8932 9154
rect 8876 9100 8932 9102
rect 8764 9042 8820 9044
rect 8764 8990 8766 9042
rect 8766 8990 8818 9042
rect 8818 8990 8820 9042
rect 8764 8988 8820 8990
rect 9324 9660 9380 9716
rect 9436 10780 9492 10836
rect 9660 10556 9716 10612
rect 10220 13916 10276 13972
rect 10668 13692 10724 13748
rect 10444 13468 10500 13524
rect 10108 12066 10164 12068
rect 10108 12014 10110 12066
rect 10110 12014 10162 12066
rect 10162 12014 10164 12066
rect 10108 12012 10164 12014
rect 10108 11564 10164 11620
rect 9884 11506 9940 11508
rect 9884 11454 9886 11506
rect 9886 11454 9938 11506
rect 9938 11454 9940 11506
rect 9884 11452 9940 11454
rect 10220 10780 10276 10836
rect 10556 12236 10612 12292
rect 9772 10332 9828 10388
rect 10220 10332 10276 10388
rect 9996 9884 10052 9940
rect 9884 9660 9940 9716
rect 9548 9548 9604 9604
rect 9548 8092 9604 8148
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 10220 8988 10276 9044
rect 11452 15314 11508 15316
rect 11452 15262 11454 15314
rect 11454 15262 11506 15314
rect 11506 15262 11508 15314
rect 11452 15260 11508 15262
rect 12572 20076 12628 20132
rect 12012 20018 12068 20020
rect 12012 19966 12014 20018
rect 12014 19966 12066 20018
rect 12066 19966 12068 20018
rect 12012 19964 12068 19966
rect 12124 19068 12180 19124
rect 11900 18508 11956 18564
rect 11676 17442 11732 17444
rect 11676 17390 11678 17442
rect 11678 17390 11730 17442
rect 11730 17390 11732 17442
rect 11676 17388 11732 17390
rect 12012 17890 12068 17892
rect 12012 17838 12014 17890
rect 12014 17838 12066 17890
rect 12066 17838 12068 17890
rect 12012 17836 12068 17838
rect 11900 15596 11956 15652
rect 12012 16492 12068 16548
rect 11788 15484 11844 15540
rect 12348 19906 12404 19908
rect 12348 19854 12350 19906
rect 12350 19854 12402 19906
rect 12402 19854 12404 19906
rect 12348 19852 12404 19854
rect 12348 19234 12404 19236
rect 12348 19182 12350 19234
rect 12350 19182 12402 19234
rect 12402 19182 12404 19234
rect 12348 19180 12404 19182
rect 12236 18620 12292 18676
rect 13020 21420 13076 21476
rect 13580 22652 13636 22708
rect 13916 23436 13972 23492
rect 14140 23714 14196 23716
rect 14140 23662 14142 23714
rect 14142 23662 14194 23714
rect 14194 23662 14196 23714
rect 14140 23660 14196 23662
rect 14028 23212 14084 23268
rect 13916 23100 13972 23156
rect 14140 22876 14196 22932
rect 13692 20802 13748 20804
rect 13692 20750 13694 20802
rect 13694 20750 13746 20802
rect 13746 20750 13748 20802
rect 13692 20748 13748 20750
rect 14700 24892 14756 24948
rect 14588 23212 14644 23268
rect 14700 24108 14756 24164
rect 14812 23436 14868 23492
rect 14476 22540 14532 22596
rect 15148 25452 15204 25508
rect 16492 32620 16548 32676
rect 16380 32396 16436 32452
rect 16268 31836 16324 31892
rect 16268 31218 16324 31220
rect 16268 31166 16270 31218
rect 16270 31166 16322 31218
rect 16322 31166 16324 31218
rect 16268 31164 16324 31166
rect 16492 31388 16548 31444
rect 16604 31500 16660 31556
rect 16492 30994 16548 30996
rect 16492 30942 16494 30994
rect 16494 30942 16546 30994
rect 16546 30942 16548 30994
rect 16492 30940 16548 30942
rect 16828 31778 16884 31780
rect 16828 31726 16830 31778
rect 16830 31726 16882 31778
rect 16882 31726 16884 31778
rect 16828 31724 16884 31726
rect 16716 31052 16772 31108
rect 16940 31388 16996 31444
rect 16380 30044 16436 30100
rect 16492 29538 16548 29540
rect 16492 29486 16494 29538
rect 16494 29486 16546 29538
rect 16546 29486 16548 29538
rect 16492 29484 16548 29486
rect 16604 29372 16660 29428
rect 16940 29596 16996 29652
rect 16716 29148 16772 29204
rect 16156 29036 16212 29092
rect 15484 26796 15540 26852
rect 15484 26572 15540 26628
rect 15036 25004 15092 25060
rect 14924 22764 14980 22820
rect 15148 23154 15204 23156
rect 15148 23102 15150 23154
rect 15150 23102 15202 23154
rect 15202 23102 15204 23154
rect 15148 23100 15204 23102
rect 15036 22540 15092 22596
rect 13132 19964 13188 20020
rect 13468 19740 13524 19796
rect 13692 19516 13748 19572
rect 13804 19404 13860 19460
rect 13916 22092 13972 22148
rect 13020 18956 13076 19012
rect 13020 18620 13076 18676
rect 12684 18508 12740 18564
rect 13132 17724 13188 17780
rect 13132 17052 13188 17108
rect 12908 16882 12964 16884
rect 12908 16830 12910 16882
rect 12910 16830 12962 16882
rect 12962 16830 12964 16882
rect 12908 16828 12964 16830
rect 12908 16604 12964 16660
rect 12684 16098 12740 16100
rect 12684 16046 12686 16098
rect 12686 16046 12738 16098
rect 12738 16046 12740 16098
rect 12684 16044 12740 16046
rect 11564 14476 11620 14532
rect 11228 14364 11284 14420
rect 11564 14028 11620 14084
rect 10892 13580 10948 13636
rect 11004 13804 11060 13860
rect 11676 13692 11732 13748
rect 11116 13580 11172 13636
rect 10780 13522 10836 13524
rect 10780 13470 10782 13522
rect 10782 13470 10834 13522
rect 10834 13470 10836 13522
rect 10780 13468 10836 13470
rect 11228 13356 11284 13412
rect 10892 12012 10948 12068
rect 10780 10668 10836 10724
rect 11788 12236 11844 12292
rect 11900 12124 11956 12180
rect 11004 10780 11060 10836
rect 10444 8930 10500 8932
rect 10444 8878 10446 8930
rect 10446 8878 10498 8930
rect 10498 8878 10500 8930
rect 10444 8876 10500 8878
rect 11228 10498 11284 10500
rect 11228 10446 11230 10498
rect 11230 10446 11282 10498
rect 11282 10446 11284 10498
rect 11228 10444 11284 10446
rect 12572 14418 12628 14420
rect 12572 14366 12574 14418
rect 12574 14366 12626 14418
rect 12626 14366 12628 14418
rect 12572 14364 12628 14366
rect 12236 13916 12292 13972
rect 12572 14028 12628 14084
rect 12460 13804 12516 13860
rect 12684 13692 12740 13748
rect 12460 12178 12516 12180
rect 12460 12126 12462 12178
rect 12462 12126 12514 12178
rect 12514 12126 12516 12178
rect 12460 12124 12516 12126
rect 11676 11004 11732 11060
rect 11676 10610 11732 10612
rect 11676 10558 11678 10610
rect 11678 10558 11730 10610
rect 11730 10558 11732 10610
rect 11676 10556 11732 10558
rect 11900 10332 11956 10388
rect 11788 10108 11844 10164
rect 11564 9996 11620 10052
rect 12124 11618 12180 11620
rect 12124 11566 12126 11618
rect 12126 11566 12178 11618
rect 12178 11566 12180 11618
rect 12124 11564 12180 11566
rect 12348 11564 12404 11620
rect 12348 11394 12404 11396
rect 12348 11342 12350 11394
rect 12350 11342 12402 11394
rect 12402 11342 12404 11394
rect 12348 11340 12404 11342
rect 13132 16380 13188 16436
rect 14028 21308 14084 21364
rect 14700 21308 14756 21364
rect 13356 18674 13412 18676
rect 13356 18622 13358 18674
rect 13358 18622 13410 18674
rect 13410 18622 13412 18674
rect 13356 18620 13412 18622
rect 14252 19122 14308 19124
rect 14252 19070 14254 19122
rect 14254 19070 14306 19122
rect 14306 19070 14308 19122
rect 14252 19068 14308 19070
rect 13468 18450 13524 18452
rect 13468 18398 13470 18450
rect 13470 18398 13522 18450
rect 13522 18398 13524 18450
rect 13468 18396 13524 18398
rect 13804 18450 13860 18452
rect 13804 18398 13806 18450
rect 13806 18398 13858 18450
rect 13858 18398 13860 18450
rect 13804 18396 13860 18398
rect 13580 17836 13636 17892
rect 14924 22092 14980 22148
rect 15820 26460 15876 26516
rect 15932 26796 15988 26852
rect 15820 26290 15876 26292
rect 15820 26238 15822 26290
rect 15822 26238 15874 26290
rect 15874 26238 15876 26290
rect 15820 26236 15876 26238
rect 15484 25788 15540 25844
rect 15596 26124 15652 26180
rect 16268 28588 16324 28644
rect 17052 28812 17108 28868
rect 17164 35308 17220 35364
rect 16604 28364 16660 28420
rect 16044 25564 16100 25620
rect 16492 26066 16548 26068
rect 16492 26014 16494 26066
rect 16494 26014 16546 26066
rect 16546 26014 16548 26066
rect 16492 26012 16548 26014
rect 16716 27746 16772 27748
rect 16716 27694 16718 27746
rect 16718 27694 16770 27746
rect 16770 27694 16772 27746
rect 16716 27692 16772 27694
rect 17612 35308 17668 35364
rect 18284 36204 18340 36260
rect 18396 36092 18452 36148
rect 18508 36316 18564 36372
rect 17276 34354 17332 34356
rect 17276 34302 17278 34354
rect 17278 34302 17330 34354
rect 17330 34302 17332 34354
rect 17276 34300 17332 34302
rect 17836 34412 17892 34468
rect 17500 34242 17556 34244
rect 17500 34190 17502 34242
rect 17502 34190 17554 34242
rect 17554 34190 17556 34242
rect 17500 34188 17556 34190
rect 17612 34130 17668 34132
rect 17612 34078 17614 34130
rect 17614 34078 17666 34130
rect 17666 34078 17668 34130
rect 17612 34076 17668 34078
rect 17388 33740 17444 33796
rect 17276 33628 17332 33684
rect 17836 33852 17892 33908
rect 17388 32620 17444 32676
rect 17612 32396 17668 32452
rect 18844 35698 18900 35700
rect 18844 35646 18846 35698
rect 18846 35646 18898 35698
rect 18898 35646 18900 35698
rect 18844 35644 18900 35646
rect 19292 41970 19348 41972
rect 19292 41918 19294 41970
rect 19294 41918 19346 41970
rect 19346 41918 19348 41970
rect 19292 41916 19348 41918
rect 20636 43820 20692 43876
rect 20636 43372 20692 43428
rect 21644 51212 21700 51268
rect 21868 52668 21924 52724
rect 21868 51324 21924 51380
rect 21756 50482 21812 50484
rect 21756 50430 21758 50482
rect 21758 50430 21810 50482
rect 21810 50430 21812 50482
rect 21756 50428 21812 50430
rect 21308 50204 21364 50260
rect 21644 50092 21700 50148
rect 21308 49644 21364 49700
rect 21532 49308 21588 49364
rect 21420 49138 21476 49140
rect 21420 49086 21422 49138
rect 21422 49086 21474 49138
rect 21474 49086 21476 49138
rect 21420 49084 21476 49086
rect 21308 47516 21364 47572
rect 21756 48860 21812 48916
rect 22204 53564 22260 53620
rect 22316 53452 22372 53508
rect 22540 54460 22596 54516
rect 22540 53788 22596 53844
rect 22764 55244 22820 55300
rect 23100 56028 23156 56084
rect 23660 56700 23716 56756
rect 24108 57596 24164 57652
rect 23996 56812 24052 56868
rect 24108 57372 24164 57428
rect 23548 56194 23604 56196
rect 23548 56142 23550 56194
rect 23550 56142 23602 56194
rect 23602 56142 23604 56194
rect 23548 56140 23604 56142
rect 23772 55410 23828 55412
rect 23772 55358 23774 55410
rect 23774 55358 23826 55410
rect 23826 55358 23828 55410
rect 23772 55356 23828 55358
rect 23884 55244 23940 55300
rect 22988 55132 23044 55188
rect 23100 55074 23156 55076
rect 23100 55022 23102 55074
rect 23102 55022 23154 55074
rect 23154 55022 23156 55074
rect 23100 55020 23156 55022
rect 23212 54684 23268 54740
rect 22764 53900 22820 53956
rect 22652 53564 22708 53620
rect 22204 53058 22260 53060
rect 22204 53006 22206 53058
rect 22206 53006 22258 53058
rect 22258 53006 22260 53058
rect 22204 53004 22260 53006
rect 22316 51100 22372 51156
rect 23212 53116 23268 53172
rect 24556 58828 24612 58884
rect 25228 59612 25284 59668
rect 25004 59164 25060 59220
rect 24668 58156 24724 58212
rect 24332 57762 24388 57764
rect 24332 57710 24334 57762
rect 24334 57710 24386 57762
rect 24386 57710 24388 57762
rect 24332 57708 24388 57710
rect 24780 57372 24836 57428
rect 24668 57260 24724 57316
rect 24444 57148 24500 57204
rect 24556 56754 24612 56756
rect 24556 56702 24558 56754
rect 24558 56702 24610 56754
rect 24610 56702 24612 56754
rect 24556 56700 24612 56702
rect 24444 56642 24500 56644
rect 24444 56590 24446 56642
rect 24446 56590 24498 56642
rect 24498 56590 24500 56642
rect 24444 56588 24500 56590
rect 24332 56364 24388 56420
rect 24220 56140 24276 56196
rect 24444 55916 24500 55972
rect 25004 58492 25060 58548
rect 25004 57596 25060 57652
rect 25116 57932 25172 57988
rect 25116 56700 25172 56756
rect 25228 57036 25284 57092
rect 24892 55916 24948 55972
rect 24332 55804 24388 55860
rect 24220 55132 24276 55188
rect 24780 55298 24836 55300
rect 24780 55246 24782 55298
rect 24782 55246 24834 55298
rect 24834 55246 24836 55298
rect 24780 55244 24836 55246
rect 25340 55410 25396 55412
rect 25340 55358 25342 55410
rect 25342 55358 25394 55410
rect 25394 55358 25396 55410
rect 25340 55356 25396 55358
rect 25228 54908 25284 54964
rect 25116 54348 25172 54404
rect 23548 54012 23604 54068
rect 23548 52780 23604 52836
rect 23548 52556 23604 52612
rect 23996 53954 24052 53956
rect 23996 53902 23998 53954
rect 23998 53902 24050 53954
rect 24050 53902 24052 53954
rect 23996 53900 24052 53902
rect 27356 59890 27412 59892
rect 27356 59838 27358 59890
rect 27358 59838 27410 59890
rect 27410 59838 27412 59890
rect 27356 59836 27412 59838
rect 26348 59612 26404 59668
rect 26236 59388 26292 59444
rect 27468 59442 27524 59444
rect 27468 59390 27470 59442
rect 27470 59390 27522 59442
rect 27522 59390 27524 59442
rect 27468 59388 27524 59390
rect 25564 59218 25620 59220
rect 25564 59166 25566 59218
rect 25566 59166 25618 59218
rect 25618 59166 25620 59218
rect 25564 59164 25620 59166
rect 26124 58994 26180 58996
rect 26124 58942 26126 58994
rect 26126 58942 26178 58994
rect 26178 58942 26180 58994
rect 26124 58940 26180 58942
rect 26796 58940 26852 58996
rect 26460 58044 26516 58100
rect 27020 58434 27076 58436
rect 27020 58382 27022 58434
rect 27022 58382 27074 58434
rect 27074 58382 27076 58434
rect 27020 58380 27076 58382
rect 26012 57650 26068 57652
rect 26012 57598 26014 57650
rect 26014 57598 26066 57650
rect 26066 57598 26068 57650
rect 26012 57596 26068 57598
rect 25676 56924 25732 56980
rect 25676 56252 25732 56308
rect 25564 56194 25620 56196
rect 25564 56142 25566 56194
rect 25566 56142 25618 56194
rect 25618 56142 25620 56194
rect 25564 56140 25620 56142
rect 26460 57260 26516 57316
rect 27020 56812 27076 56868
rect 28140 59724 28196 59780
rect 27804 59164 27860 59220
rect 27916 59052 27972 59108
rect 27804 58940 27860 58996
rect 27804 58434 27860 58436
rect 27804 58382 27806 58434
rect 27806 58382 27858 58434
rect 27858 58382 27860 58434
rect 27804 58380 27860 58382
rect 28028 58604 28084 58660
rect 27580 56866 27636 56868
rect 27580 56814 27582 56866
rect 27582 56814 27634 56866
rect 27634 56814 27636 56866
rect 27580 56812 27636 56814
rect 27692 56924 27748 56980
rect 25900 56082 25956 56084
rect 25900 56030 25902 56082
rect 25902 56030 25954 56082
rect 25954 56030 25956 56082
rect 25900 56028 25956 56030
rect 28028 57708 28084 57764
rect 28364 58716 28420 58772
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 29596 59948 29652 60004
rect 33964 60002 34020 60004
rect 33964 59950 33966 60002
rect 33966 59950 34018 60002
rect 34018 59950 34020 60002
rect 33964 59948 34020 59950
rect 34972 60002 35028 60004
rect 34972 59950 34974 60002
rect 34974 59950 35026 60002
rect 35026 59950 35028 60002
rect 34972 59948 35028 59950
rect 29708 59836 29764 59892
rect 28588 58380 28644 58436
rect 29148 59612 29204 59668
rect 27468 55858 27524 55860
rect 27468 55806 27470 55858
rect 27470 55806 27522 55858
rect 27522 55806 27524 55858
rect 27468 55804 27524 55806
rect 24220 52892 24276 52948
rect 23996 51884 24052 51940
rect 22764 50540 22820 50596
rect 22092 48412 22148 48468
rect 22316 48300 22372 48356
rect 22204 47628 22260 47684
rect 21308 46562 21364 46564
rect 21308 46510 21310 46562
rect 21310 46510 21362 46562
rect 21362 46510 21364 46562
rect 21308 46508 21364 46510
rect 21420 46450 21476 46452
rect 21420 46398 21422 46450
rect 21422 46398 21474 46450
rect 21474 46398 21476 46450
rect 21420 46396 21476 46398
rect 21756 46620 21812 46676
rect 21420 45388 21476 45444
rect 22092 46172 22148 46228
rect 21980 45164 22036 45220
rect 23324 48466 23380 48468
rect 23324 48414 23326 48466
rect 23326 48414 23378 48466
rect 23378 48414 23380 48466
rect 23324 48412 23380 48414
rect 23996 51324 24052 51380
rect 24220 52556 24276 52612
rect 24332 52162 24388 52164
rect 24332 52110 24334 52162
rect 24334 52110 24386 52162
rect 24386 52110 24388 52162
rect 24332 52108 24388 52110
rect 25228 53564 25284 53620
rect 25676 55020 25732 55076
rect 26572 55356 26628 55412
rect 25452 53900 25508 53956
rect 26236 54460 26292 54516
rect 25900 53788 25956 53844
rect 25340 53340 25396 53396
rect 25340 52780 25396 52836
rect 25788 53170 25844 53172
rect 25788 53118 25790 53170
rect 25790 53118 25842 53170
rect 25842 53118 25844 53170
rect 25788 53116 25844 53118
rect 25452 52108 25508 52164
rect 24444 51548 24500 51604
rect 22540 47570 22596 47572
rect 22540 47518 22542 47570
rect 22542 47518 22594 47570
rect 22594 47518 22596 47570
rect 22540 47516 22596 47518
rect 24108 50204 24164 50260
rect 23884 48748 23940 48804
rect 23772 48300 23828 48356
rect 23548 47740 23604 47796
rect 23660 47964 23716 48020
rect 22988 46844 23044 46900
rect 23324 46844 23380 46900
rect 22876 46786 22932 46788
rect 22876 46734 22878 46786
rect 22878 46734 22930 46786
rect 22930 46734 22932 46786
rect 22876 46732 22932 46734
rect 23324 46674 23380 46676
rect 23324 46622 23326 46674
rect 23326 46622 23378 46674
rect 23378 46622 23380 46674
rect 23324 46620 23380 46622
rect 23212 45612 23268 45668
rect 21756 44380 21812 44436
rect 21196 42700 21252 42756
rect 20524 42364 20580 42420
rect 20860 42476 20916 42532
rect 20300 41916 20356 41972
rect 19068 40908 19124 40964
rect 19404 41804 19460 41860
rect 20748 41970 20804 41972
rect 20748 41918 20750 41970
rect 20750 41918 20802 41970
rect 20802 41918 20804 41970
rect 20748 41916 20804 41918
rect 20524 41804 20580 41860
rect 19740 41746 19796 41748
rect 19740 41694 19742 41746
rect 19742 41694 19794 41746
rect 19794 41694 19796 41746
rect 19740 41692 19796 41694
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19068 40236 19124 40292
rect 19404 39228 19460 39284
rect 19180 38834 19236 38836
rect 19180 38782 19182 38834
rect 19182 38782 19234 38834
rect 19234 38782 19236 38834
rect 19180 38780 19236 38782
rect 20188 40236 20244 40292
rect 20412 40348 20468 40404
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20636 41020 20692 41076
rect 20636 40796 20692 40852
rect 21756 43596 21812 43652
rect 22652 44994 22708 44996
rect 22652 44942 22654 44994
rect 22654 44942 22706 44994
rect 22706 44942 22708 44994
rect 22652 44940 22708 44942
rect 22876 44716 22932 44772
rect 21868 43484 21924 43540
rect 21532 43036 21588 43092
rect 22316 44322 22372 44324
rect 22316 44270 22318 44322
rect 22318 44270 22370 44322
rect 22370 44270 22372 44322
rect 22316 44268 22372 44270
rect 22092 43484 22148 43540
rect 21980 42924 22036 42980
rect 21420 42082 21476 42084
rect 21420 42030 21422 42082
rect 21422 42030 21474 42082
rect 21474 42030 21476 42082
rect 21420 42028 21476 42030
rect 21980 42530 22036 42532
rect 21980 42478 21982 42530
rect 21982 42478 22034 42530
rect 22034 42478 22036 42530
rect 21980 42476 22036 42478
rect 21756 42140 21812 42196
rect 21644 41804 21700 41860
rect 22428 41970 22484 41972
rect 22428 41918 22430 41970
rect 22430 41918 22482 41970
rect 22482 41918 22484 41970
rect 22428 41916 22484 41918
rect 21868 41804 21924 41860
rect 21644 40908 21700 40964
rect 21756 41074 21812 41076
rect 21756 41022 21758 41074
rect 21758 41022 21810 41074
rect 21810 41022 21812 41074
rect 21756 41020 21812 41022
rect 22652 42924 22708 42980
rect 22540 41804 22596 41860
rect 22092 41746 22148 41748
rect 22092 41694 22094 41746
rect 22094 41694 22146 41746
rect 22146 41694 22148 41746
rect 22092 41692 22148 41694
rect 23100 45052 23156 45108
rect 23324 45276 23380 45332
rect 23436 45106 23492 45108
rect 23436 45054 23438 45106
rect 23438 45054 23490 45106
rect 23490 45054 23492 45106
rect 23436 45052 23492 45054
rect 23996 48412 24052 48468
rect 23996 47740 24052 47796
rect 23884 46172 23940 46228
rect 23548 44604 23604 44660
rect 23772 46060 23828 46116
rect 23996 45836 24052 45892
rect 23884 45500 23940 45556
rect 25452 51660 25508 51716
rect 25228 51602 25284 51604
rect 25228 51550 25230 51602
rect 25230 51550 25282 51602
rect 25282 51550 25284 51602
rect 25228 51548 25284 51550
rect 24780 51324 24836 51380
rect 26012 52444 26068 52500
rect 27580 55580 27636 55636
rect 26684 55186 26740 55188
rect 26684 55134 26686 55186
rect 26686 55134 26738 55186
rect 26738 55134 26740 55186
rect 26684 55132 26740 55134
rect 26908 55074 26964 55076
rect 26908 55022 26910 55074
rect 26910 55022 26962 55074
rect 26962 55022 26964 55074
rect 26908 55020 26964 55022
rect 26572 53900 26628 53956
rect 26684 53730 26740 53732
rect 26684 53678 26686 53730
rect 26686 53678 26738 53730
rect 26738 53678 26740 53730
rect 26684 53676 26740 53678
rect 27132 55298 27188 55300
rect 27132 55246 27134 55298
rect 27134 55246 27186 55298
rect 27186 55246 27188 55298
rect 27132 55244 27188 55246
rect 27468 55356 27524 55412
rect 27244 54236 27300 54292
rect 27356 53788 27412 53844
rect 27804 55692 27860 55748
rect 27916 55468 27972 55524
rect 28140 55692 28196 55748
rect 27804 54572 27860 54628
rect 27692 54124 27748 54180
rect 26460 53452 26516 53508
rect 27692 53954 27748 53956
rect 27692 53902 27694 53954
rect 27694 53902 27746 53954
rect 27746 53902 27748 53954
rect 27692 53900 27748 53902
rect 27020 53170 27076 53172
rect 27020 53118 27022 53170
rect 27022 53118 27074 53170
rect 27074 53118 27076 53170
rect 27020 53116 27076 53118
rect 26572 52444 26628 52500
rect 25564 51548 25620 51604
rect 24556 49980 24612 50036
rect 24444 47458 24500 47460
rect 24444 47406 24446 47458
rect 24446 47406 24498 47458
rect 24498 47406 24500 47458
rect 24444 47404 24500 47406
rect 24780 48748 24836 48804
rect 25004 47628 25060 47684
rect 24668 46956 24724 47012
rect 24332 46674 24388 46676
rect 24332 46622 24334 46674
rect 24334 46622 24386 46674
rect 24386 46622 24388 46674
rect 24332 46620 24388 46622
rect 24556 46786 24612 46788
rect 24556 46734 24558 46786
rect 24558 46734 24610 46786
rect 24610 46734 24612 46786
rect 24556 46732 24612 46734
rect 24108 45276 24164 45332
rect 24556 45890 24612 45892
rect 24556 45838 24558 45890
rect 24558 45838 24610 45890
rect 24610 45838 24612 45890
rect 24556 45836 24612 45838
rect 26348 51602 26404 51604
rect 26348 51550 26350 51602
rect 26350 51550 26402 51602
rect 26402 51550 26404 51602
rect 26348 51548 26404 51550
rect 26796 51772 26852 51828
rect 27020 52556 27076 52612
rect 26796 51378 26852 51380
rect 26796 51326 26798 51378
rect 26798 51326 26850 51378
rect 26850 51326 26852 51378
rect 26796 51324 26852 51326
rect 25788 50988 25844 51044
rect 25676 50034 25732 50036
rect 25676 49982 25678 50034
rect 25678 49982 25730 50034
rect 25730 49982 25732 50034
rect 25676 49980 25732 49982
rect 25340 49084 25396 49140
rect 25452 48802 25508 48804
rect 25452 48750 25454 48802
rect 25454 48750 25506 48802
rect 25506 48750 25508 48802
rect 25452 48748 25508 48750
rect 24780 46114 24836 46116
rect 24780 46062 24782 46114
rect 24782 46062 24834 46114
rect 24834 46062 24836 46114
rect 24780 46060 24836 46062
rect 24780 45276 24836 45332
rect 23996 45106 24052 45108
rect 23996 45054 23998 45106
rect 23998 45054 24050 45106
rect 24050 45054 24052 45106
rect 23996 45052 24052 45054
rect 23212 44268 23268 44324
rect 23100 42754 23156 42756
rect 23100 42702 23102 42754
rect 23102 42702 23154 42754
rect 23154 42702 23156 42754
rect 23100 42700 23156 42702
rect 23212 43596 23268 43652
rect 22652 41356 22708 41412
rect 22540 41132 22596 41188
rect 22204 40572 22260 40628
rect 22092 40460 22148 40516
rect 21420 40402 21476 40404
rect 21420 40350 21422 40402
rect 21422 40350 21474 40402
rect 21474 40350 21476 40402
rect 21420 40348 21476 40350
rect 20076 38892 20132 38948
rect 19404 37884 19460 37940
rect 19516 38332 19572 38388
rect 19292 35980 19348 36036
rect 20412 38556 20468 38612
rect 19852 38050 19908 38052
rect 19852 37998 19854 38050
rect 19854 37998 19906 38050
rect 19906 37998 19908 38050
rect 19852 37996 19908 37998
rect 20748 37996 20804 38052
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20188 36988 20244 37044
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19628 35698 19684 35700
rect 19628 35646 19630 35698
rect 19630 35646 19682 35698
rect 19682 35646 19684 35698
rect 19628 35644 19684 35646
rect 20300 36652 20356 36708
rect 20300 36428 20356 36484
rect 20412 37772 20468 37828
rect 18620 34860 18676 34916
rect 18172 34242 18228 34244
rect 18172 34190 18174 34242
rect 18174 34190 18226 34242
rect 18226 34190 18228 34242
rect 18172 34188 18228 34190
rect 18396 34636 18452 34692
rect 18172 33852 18228 33908
rect 18060 32172 18116 32228
rect 18172 33068 18228 33124
rect 17836 31778 17892 31780
rect 17836 31726 17838 31778
rect 17838 31726 17890 31778
rect 17890 31726 17892 31778
rect 17836 31724 17892 31726
rect 17500 31388 17556 31444
rect 17836 31106 17892 31108
rect 17836 31054 17838 31106
rect 17838 31054 17890 31106
rect 17890 31054 17892 31106
rect 17836 31052 17892 31054
rect 17276 28924 17332 28980
rect 17388 28700 17444 28756
rect 17276 28476 17332 28532
rect 16940 26908 16996 26964
rect 17052 26684 17108 26740
rect 17276 26572 17332 26628
rect 16828 25116 16884 25172
rect 15596 24444 15652 24500
rect 15372 22876 15428 22932
rect 15820 22540 15876 22596
rect 15260 22204 15316 22260
rect 15596 21698 15652 21700
rect 15596 21646 15598 21698
rect 15598 21646 15650 21698
rect 15650 21646 15652 21698
rect 15596 21644 15652 21646
rect 15596 21084 15652 21140
rect 14812 20972 14868 21028
rect 14476 20690 14532 20692
rect 14476 20638 14478 20690
rect 14478 20638 14530 20690
rect 14530 20638 14532 20690
rect 14476 20636 14532 20638
rect 15932 21308 15988 21364
rect 14924 20636 14980 20692
rect 15036 20748 15092 20804
rect 14364 18396 14420 18452
rect 14476 20300 14532 20356
rect 14364 17778 14420 17780
rect 14364 17726 14366 17778
rect 14366 17726 14418 17778
rect 14418 17726 14420 17778
rect 14364 17724 14420 17726
rect 13804 16940 13860 16996
rect 13244 16156 13300 16212
rect 13580 16828 13636 16884
rect 13468 16098 13524 16100
rect 13468 16046 13470 16098
rect 13470 16046 13522 16098
rect 13522 16046 13524 16098
rect 13468 16044 13524 16046
rect 14140 16828 14196 16884
rect 14252 16940 14308 16996
rect 14700 20076 14756 20132
rect 14700 19740 14756 19796
rect 14588 19404 14644 19460
rect 15484 20748 15540 20804
rect 15036 18620 15092 18676
rect 15372 20690 15428 20692
rect 15372 20638 15374 20690
rect 15374 20638 15426 20690
rect 15426 20638 15428 20690
rect 15372 20636 15428 20638
rect 16156 22316 16212 22372
rect 16268 21362 16324 21364
rect 16268 21310 16270 21362
rect 16270 21310 16322 21362
rect 16322 21310 16324 21362
rect 16268 21308 16324 21310
rect 16044 20748 16100 20804
rect 15596 20524 15652 20580
rect 15484 20076 15540 20132
rect 15372 20018 15428 20020
rect 15372 19966 15374 20018
rect 15374 19966 15426 20018
rect 15426 19966 15428 20018
rect 15372 19964 15428 19966
rect 15148 18396 15204 18452
rect 16604 24946 16660 24948
rect 16604 24894 16606 24946
rect 16606 24894 16658 24946
rect 16658 24894 16660 24946
rect 16604 24892 16660 24894
rect 16828 24722 16884 24724
rect 16828 24670 16830 24722
rect 16830 24670 16882 24722
rect 16882 24670 16884 24722
rect 16828 24668 16884 24670
rect 16604 24556 16660 24612
rect 16492 23660 16548 23716
rect 16716 23660 16772 23716
rect 16716 23324 16772 23380
rect 17612 26236 17668 26292
rect 17724 26460 17780 26516
rect 17052 26124 17108 26180
rect 17052 25506 17108 25508
rect 17052 25454 17054 25506
rect 17054 25454 17106 25506
rect 17106 25454 17108 25506
rect 17052 25452 17108 25454
rect 17612 26012 17668 26068
rect 17724 25564 17780 25620
rect 16940 22876 16996 22932
rect 16940 22428 16996 22484
rect 16828 22204 16884 22260
rect 16940 22146 16996 22148
rect 16940 22094 16942 22146
rect 16942 22094 16994 22146
rect 16994 22094 16996 22146
rect 16940 22092 16996 22094
rect 15596 19964 15652 20020
rect 16492 21084 16548 21140
rect 16492 20524 16548 20580
rect 15708 19234 15764 19236
rect 15708 19182 15710 19234
rect 15710 19182 15762 19234
rect 15762 19182 15764 19234
rect 15708 19180 15764 19182
rect 15484 18620 15540 18676
rect 15260 17890 15316 17892
rect 15260 17838 15262 17890
rect 15262 17838 15314 17890
rect 15314 17838 15316 17890
rect 15260 17836 15316 17838
rect 16044 18172 16100 18228
rect 15596 17500 15652 17556
rect 15484 17106 15540 17108
rect 15484 17054 15486 17106
rect 15486 17054 15538 17106
rect 15538 17054 15540 17106
rect 15484 17052 15540 17054
rect 16044 17052 16100 17108
rect 14476 16380 14532 16436
rect 13916 16322 13972 16324
rect 13916 16270 13918 16322
rect 13918 16270 13970 16322
rect 13970 16270 13972 16322
rect 13916 16268 13972 16270
rect 14028 16098 14084 16100
rect 14028 16046 14030 16098
rect 14030 16046 14082 16098
rect 14082 16046 14084 16098
rect 14028 16044 14084 16046
rect 13132 13804 13188 13860
rect 13132 12290 13188 12292
rect 13132 12238 13134 12290
rect 13134 12238 13186 12290
rect 13186 12238 13188 12290
rect 13132 12236 13188 12238
rect 12684 11564 12740 11620
rect 12572 11452 12628 11508
rect 12460 10834 12516 10836
rect 12460 10782 12462 10834
rect 12462 10782 12514 10834
rect 12514 10782 12516 10834
rect 12460 10780 12516 10782
rect 12460 10610 12516 10612
rect 12460 10558 12462 10610
rect 12462 10558 12514 10610
rect 12514 10558 12516 10610
rect 12460 10556 12516 10558
rect 12236 10444 12292 10500
rect 12124 10220 12180 10276
rect 11564 8876 11620 8932
rect 11004 8258 11060 8260
rect 11004 8206 11006 8258
rect 11006 8206 11058 8258
rect 11058 8206 11060 8258
rect 11004 8204 11060 8206
rect 11564 8204 11620 8260
rect 10892 8092 10948 8148
rect 10892 6802 10948 6804
rect 10892 6750 10894 6802
rect 10894 6750 10946 6802
rect 10946 6750 10948 6802
rect 10892 6748 10948 6750
rect 12012 9212 12068 9268
rect 11676 7308 11732 7364
rect 11788 6748 11844 6804
rect 11676 6690 11732 6692
rect 11676 6638 11678 6690
rect 11678 6638 11730 6690
rect 11730 6638 11732 6690
rect 11676 6636 11732 6638
rect 12236 6636 12292 6692
rect 12572 8316 12628 8372
rect 12460 8258 12516 8260
rect 12460 8206 12462 8258
rect 12462 8206 12514 8258
rect 12514 8206 12516 8258
rect 12460 8204 12516 8206
rect 13020 11004 13076 11060
rect 13132 11340 13188 11396
rect 13020 10780 13076 10836
rect 13356 11394 13412 11396
rect 13356 11342 13358 11394
rect 13358 11342 13410 11394
rect 13410 11342 13412 11394
rect 13356 11340 13412 11342
rect 13244 11116 13300 11172
rect 13244 10892 13300 10948
rect 13580 14754 13636 14756
rect 13580 14702 13582 14754
rect 13582 14702 13634 14754
rect 13634 14702 13636 14754
rect 13580 14700 13636 14702
rect 13804 15426 13860 15428
rect 13804 15374 13806 15426
rect 13806 15374 13858 15426
rect 13858 15374 13860 15426
rect 13804 15372 13860 15374
rect 15484 16882 15540 16884
rect 15484 16830 15486 16882
rect 15486 16830 15538 16882
rect 15538 16830 15540 16882
rect 15484 16828 15540 16830
rect 15372 16716 15428 16772
rect 15708 15372 15764 15428
rect 13804 14924 13860 14980
rect 13804 14418 13860 14420
rect 13804 14366 13806 14418
rect 13806 14366 13858 14418
rect 13858 14366 13860 14418
rect 13804 14364 13860 14366
rect 14700 14700 14756 14756
rect 13692 13468 13748 13524
rect 13580 12290 13636 12292
rect 13580 12238 13582 12290
rect 13582 12238 13634 12290
rect 13634 12238 13636 12290
rect 13580 12236 13636 12238
rect 13132 10444 13188 10500
rect 12796 9884 12852 9940
rect 13020 10220 13076 10276
rect 13020 9266 13076 9268
rect 13020 9214 13022 9266
rect 13022 9214 13074 9266
rect 13074 9214 13076 9266
rect 13020 9212 13076 9214
rect 12796 8258 12852 8260
rect 12796 8206 12798 8258
rect 12798 8206 12850 8258
rect 12850 8206 12852 8258
rect 12796 8204 12852 8206
rect 12796 6524 12852 6580
rect 13580 11004 13636 11060
rect 14476 14476 14532 14532
rect 14588 13692 14644 13748
rect 14364 13468 14420 13524
rect 14252 12908 14308 12964
rect 14028 12850 14084 12852
rect 14028 12798 14030 12850
rect 14030 12798 14082 12850
rect 14082 12798 14084 12850
rect 14028 12796 14084 12798
rect 13804 12178 13860 12180
rect 13804 12126 13806 12178
rect 13806 12126 13858 12178
rect 13858 12126 13860 12178
rect 13804 12124 13860 12126
rect 14028 11564 14084 11620
rect 13692 10780 13748 10836
rect 13916 11340 13972 11396
rect 13580 10332 13636 10388
rect 13804 10108 13860 10164
rect 14588 12178 14644 12180
rect 14588 12126 14590 12178
rect 14590 12126 14642 12178
rect 14642 12126 14644 12178
rect 14588 12124 14644 12126
rect 14476 10556 14532 10612
rect 14364 9602 14420 9604
rect 14364 9550 14366 9602
rect 14366 9550 14418 9602
rect 14418 9550 14420 9602
rect 14364 9548 14420 9550
rect 14252 9212 14308 9268
rect 14924 14530 14980 14532
rect 14924 14478 14926 14530
rect 14926 14478 14978 14530
rect 14978 14478 14980 14530
rect 14924 14476 14980 14478
rect 14812 14364 14868 14420
rect 15596 14418 15652 14420
rect 15596 14366 15598 14418
rect 15598 14366 15650 14418
rect 15650 14366 15652 14418
rect 15596 14364 15652 14366
rect 15260 14306 15316 14308
rect 15260 14254 15262 14306
rect 15262 14254 15314 14306
rect 15314 14254 15316 14306
rect 15260 14252 15316 14254
rect 15036 13746 15092 13748
rect 15036 13694 15038 13746
rect 15038 13694 15090 13746
rect 15090 13694 15092 13746
rect 15036 13692 15092 13694
rect 15260 12290 15316 12292
rect 15260 12238 15262 12290
rect 15262 12238 15314 12290
rect 15314 12238 15316 12290
rect 15260 12236 15316 12238
rect 15036 12178 15092 12180
rect 15036 12126 15038 12178
rect 15038 12126 15090 12178
rect 15090 12126 15092 12178
rect 15036 12124 15092 12126
rect 14140 8316 14196 8372
rect 13580 6748 13636 6804
rect 13468 6690 13524 6692
rect 13468 6638 13470 6690
rect 13470 6638 13522 6690
rect 13522 6638 13524 6690
rect 13468 6636 13524 6638
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 13804 6578 13860 6580
rect 13804 6526 13806 6578
rect 13806 6526 13858 6578
rect 13858 6526 13860 6578
rect 13804 6524 13860 6526
rect 14700 9884 14756 9940
rect 14812 9100 14868 9156
rect 14588 6636 14644 6692
rect 14700 6972 14756 7028
rect 15148 11564 15204 11620
rect 15148 10668 15204 10724
rect 15036 9826 15092 9828
rect 15036 9774 15038 9826
rect 15038 9774 15090 9826
rect 15090 9774 15092 9826
rect 15036 9772 15092 9774
rect 15932 16156 15988 16212
rect 16044 14364 16100 14420
rect 16268 19964 16324 20020
rect 16604 20690 16660 20692
rect 16604 20638 16606 20690
rect 16606 20638 16658 20690
rect 16658 20638 16660 20690
rect 16604 20636 16660 20638
rect 16716 19964 16772 20020
rect 16828 20972 16884 21028
rect 16492 18396 16548 18452
rect 16268 18172 16324 18228
rect 16940 19346 16996 19348
rect 16940 19294 16942 19346
rect 16942 19294 16994 19346
rect 16994 19294 16996 19346
rect 16940 19292 16996 19294
rect 16828 19234 16884 19236
rect 16828 19182 16830 19234
rect 16830 19182 16882 19234
rect 16882 19182 16884 19234
rect 16828 19180 16884 19182
rect 16940 18338 16996 18340
rect 16940 18286 16942 18338
rect 16942 18286 16994 18338
rect 16994 18286 16996 18338
rect 16940 18284 16996 18286
rect 16604 17612 16660 17668
rect 18060 28476 18116 28532
rect 18172 28364 18228 28420
rect 18508 33740 18564 33796
rect 18508 32508 18564 32564
rect 19068 33458 19124 33460
rect 19068 33406 19070 33458
rect 19070 33406 19122 33458
rect 19122 33406 19124 33458
rect 19068 33404 19124 33406
rect 19068 33234 19124 33236
rect 19068 33182 19070 33234
rect 19070 33182 19122 33234
rect 19122 33182 19124 33234
rect 19068 33180 19124 33182
rect 18732 32396 18788 32452
rect 19068 32284 19124 32340
rect 18508 31612 18564 31668
rect 18732 31164 18788 31220
rect 19068 31164 19124 31220
rect 18508 30940 18564 30996
rect 18620 28700 18676 28756
rect 18060 28028 18116 28084
rect 17948 25676 18004 25732
rect 19292 33740 19348 33796
rect 19180 29484 19236 29540
rect 19068 28642 19124 28644
rect 19068 28590 19070 28642
rect 19070 28590 19122 28642
rect 19122 28590 19124 28642
rect 19068 28588 19124 28590
rect 18620 27916 18676 27972
rect 18732 27692 18788 27748
rect 18844 27020 18900 27076
rect 18732 26962 18788 26964
rect 18732 26910 18734 26962
rect 18734 26910 18786 26962
rect 18786 26910 18788 26962
rect 18732 26908 18788 26910
rect 18396 26460 18452 26516
rect 18732 25900 18788 25956
rect 18060 25340 18116 25396
rect 18508 25564 18564 25620
rect 18060 25116 18116 25172
rect 17500 24722 17556 24724
rect 17500 24670 17502 24722
rect 17502 24670 17554 24722
rect 17554 24670 17556 24722
rect 17500 24668 17556 24670
rect 17388 23436 17444 23492
rect 17724 24108 17780 24164
rect 17276 22428 17332 22484
rect 17612 22204 17668 22260
rect 18396 25452 18452 25508
rect 18396 25116 18452 25172
rect 17836 23324 17892 23380
rect 18060 23212 18116 23268
rect 18284 23154 18340 23156
rect 18284 23102 18286 23154
rect 18286 23102 18338 23154
rect 18338 23102 18340 23154
rect 18284 23100 18340 23102
rect 18060 22876 18116 22932
rect 17612 21698 17668 21700
rect 17612 21646 17614 21698
rect 17614 21646 17666 21698
rect 17666 21646 17668 21698
rect 17612 21644 17668 21646
rect 17388 21026 17444 21028
rect 17388 20974 17390 21026
rect 17390 20974 17442 21026
rect 17442 20974 17444 21026
rect 17388 20972 17444 20974
rect 17276 20860 17332 20916
rect 17276 20412 17332 20468
rect 16492 17500 16548 17556
rect 16268 16994 16324 16996
rect 16268 16942 16270 16994
rect 16270 16942 16322 16994
rect 16322 16942 16324 16994
rect 16268 16940 16324 16942
rect 16716 16994 16772 16996
rect 16716 16942 16718 16994
rect 16718 16942 16770 16994
rect 16770 16942 16772 16994
rect 16716 16940 16772 16942
rect 16492 16156 16548 16212
rect 16268 15372 16324 15428
rect 15820 13804 15876 13860
rect 16268 14252 16324 14308
rect 15596 13580 15652 13636
rect 15484 13132 15540 13188
rect 15596 12348 15652 12404
rect 15484 9996 15540 10052
rect 15260 8652 15316 8708
rect 14924 6524 14980 6580
rect 13916 5964 13972 6020
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 15260 8316 15316 8372
rect 15260 7420 15316 7476
rect 15372 6578 15428 6580
rect 15372 6526 15374 6578
rect 15374 6526 15426 6578
rect 15426 6526 15428 6578
rect 15372 6524 15428 6526
rect 15932 11900 15988 11956
rect 16380 13692 16436 13748
rect 16940 13804 16996 13860
rect 16380 13468 16436 13524
rect 16604 12962 16660 12964
rect 16604 12910 16606 12962
rect 16606 12910 16658 12962
rect 16658 12910 16660 12962
rect 16604 12908 16660 12910
rect 16492 12796 16548 12852
rect 16492 12236 16548 12292
rect 16268 12178 16324 12180
rect 16268 12126 16270 12178
rect 16270 12126 16322 12178
rect 16322 12126 16324 12178
rect 16268 12124 16324 12126
rect 17836 21308 17892 21364
rect 17948 20524 18004 20580
rect 19292 29372 19348 29428
rect 19180 27804 19236 27860
rect 19068 27186 19124 27188
rect 19068 27134 19070 27186
rect 19070 27134 19122 27186
rect 19122 27134 19124 27186
rect 19068 27132 19124 27134
rect 18956 25676 19012 25732
rect 19292 27020 19348 27076
rect 19964 34972 20020 35028
rect 20524 36594 20580 36596
rect 20524 36542 20526 36594
rect 20526 36542 20578 36594
rect 20578 36542 20580 36594
rect 20524 36540 20580 36542
rect 21308 39452 21364 39508
rect 21084 37996 21140 38052
rect 21196 38780 21252 38836
rect 22652 40796 22708 40852
rect 22428 40012 22484 40068
rect 22316 39506 22372 39508
rect 22316 39454 22318 39506
rect 22318 39454 22370 39506
rect 22370 39454 22372 39506
rect 22316 39452 22372 39454
rect 22204 38668 22260 38724
rect 21532 38332 21588 38388
rect 21532 38050 21588 38052
rect 21532 37998 21534 38050
rect 21534 37998 21586 38050
rect 21586 37998 21588 38050
rect 21532 37996 21588 37998
rect 21420 37938 21476 37940
rect 21420 37886 21422 37938
rect 21422 37886 21474 37938
rect 21474 37886 21476 37938
rect 21420 37884 21476 37886
rect 20748 36876 20804 36932
rect 20636 36316 20692 36372
rect 22652 38722 22708 38724
rect 22652 38670 22654 38722
rect 22654 38670 22706 38722
rect 22706 38670 22708 38722
rect 22652 38668 22708 38670
rect 22540 38332 22596 38388
rect 21644 36482 21700 36484
rect 21644 36430 21646 36482
rect 21646 36430 21698 36482
rect 21698 36430 21700 36482
rect 21644 36428 21700 36430
rect 21532 36258 21588 36260
rect 21532 36206 21534 36258
rect 21534 36206 21586 36258
rect 21586 36206 21588 36258
rect 21532 36204 21588 36206
rect 20860 35532 20916 35588
rect 20076 34690 20132 34692
rect 20076 34638 20078 34690
rect 20078 34638 20130 34690
rect 20130 34638 20132 34690
rect 20076 34636 20132 34638
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19852 33628 19908 33684
rect 20748 34802 20804 34804
rect 20748 34750 20750 34802
rect 20750 34750 20802 34802
rect 20802 34750 20804 34802
rect 20748 34748 20804 34750
rect 20972 35644 21028 35700
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20412 31948 20468 32004
rect 20300 31724 20356 31780
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19516 30268 19572 30324
rect 20300 30492 20356 30548
rect 19852 30210 19908 30212
rect 19852 30158 19854 30210
rect 19854 30158 19906 30210
rect 19906 30158 19908 30210
rect 19852 30156 19908 30158
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20524 29820 20580 29876
rect 20044 29764 20100 29766
rect 19516 28812 19572 28868
rect 19740 29036 19796 29092
rect 20300 28866 20356 28868
rect 20300 28814 20302 28866
rect 20302 28814 20354 28866
rect 20354 28814 20356 28866
rect 20300 28812 20356 28814
rect 20524 28812 20580 28868
rect 19964 28700 20020 28756
rect 19628 28588 19684 28644
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20748 33068 20804 33124
rect 20860 32396 20916 32452
rect 23660 44322 23716 44324
rect 23660 44270 23662 44322
rect 23662 44270 23714 44322
rect 23714 44270 23716 44322
rect 23660 44268 23716 44270
rect 23436 42642 23492 42644
rect 23436 42590 23438 42642
rect 23438 42590 23490 42642
rect 23490 42590 23492 42642
rect 23436 42588 23492 42590
rect 23772 43036 23828 43092
rect 24108 44268 24164 44324
rect 24108 43260 24164 43316
rect 23996 42924 24052 42980
rect 23436 41970 23492 41972
rect 23436 41918 23438 41970
rect 23438 41918 23490 41970
rect 23490 41918 23492 41970
rect 23436 41916 23492 41918
rect 23100 41356 23156 41412
rect 22988 41074 23044 41076
rect 22988 41022 22990 41074
rect 22990 41022 23042 41074
rect 23042 41022 23044 41074
rect 22988 41020 23044 41022
rect 23212 40012 23268 40068
rect 24108 42140 24164 42196
rect 24668 45106 24724 45108
rect 24668 45054 24670 45106
rect 24670 45054 24722 45106
rect 24722 45054 24724 45106
rect 24668 45052 24724 45054
rect 24780 44604 24836 44660
rect 24556 44434 24612 44436
rect 24556 44382 24558 44434
rect 24558 44382 24610 44434
rect 24610 44382 24612 44434
rect 24556 44380 24612 44382
rect 24444 44268 24500 44324
rect 24556 43426 24612 43428
rect 24556 43374 24558 43426
rect 24558 43374 24610 43426
rect 24610 43374 24612 43426
rect 24556 43372 24612 43374
rect 24556 42252 24612 42308
rect 24220 41692 24276 41748
rect 23884 41468 23940 41524
rect 24444 41580 24500 41636
rect 24332 41186 24388 41188
rect 24332 41134 24334 41186
rect 24334 41134 24386 41186
rect 24386 41134 24388 41186
rect 24332 41132 24388 41134
rect 23660 40572 23716 40628
rect 23996 40908 24052 40964
rect 23884 40124 23940 40180
rect 24108 40796 24164 40852
rect 24220 40684 24276 40740
rect 23548 38946 23604 38948
rect 23548 38894 23550 38946
rect 23550 38894 23602 38946
rect 23602 38894 23604 38946
rect 23548 38892 23604 38894
rect 23996 38780 24052 38836
rect 23324 38556 23380 38612
rect 22764 37772 22820 37828
rect 22428 36876 22484 36932
rect 22652 37100 22708 37156
rect 22316 36482 22372 36484
rect 22316 36430 22318 36482
rect 22318 36430 22370 36482
rect 22370 36430 22372 36482
rect 22316 36428 22372 36430
rect 21980 36316 22036 36372
rect 22428 35644 22484 35700
rect 21868 35532 21924 35588
rect 21420 34636 21476 34692
rect 21084 33628 21140 33684
rect 21420 32620 21476 32676
rect 22092 33852 22148 33908
rect 21868 33234 21924 33236
rect 21868 33182 21870 33234
rect 21870 33182 21922 33234
rect 21922 33182 21924 33234
rect 21868 33180 21924 33182
rect 21196 32338 21252 32340
rect 21196 32286 21198 32338
rect 21198 32286 21250 32338
rect 21250 32286 21252 32338
rect 21196 32284 21252 32286
rect 20748 30716 20804 30772
rect 21084 30994 21140 30996
rect 21084 30942 21086 30994
rect 21086 30942 21138 30994
rect 21138 30942 21140 30994
rect 21084 30940 21140 30942
rect 20860 29986 20916 29988
rect 20860 29934 20862 29986
rect 20862 29934 20914 29986
rect 20914 29934 20916 29986
rect 20860 29932 20916 29934
rect 20748 29426 20804 29428
rect 20748 29374 20750 29426
rect 20750 29374 20802 29426
rect 20802 29374 20804 29426
rect 20748 29372 20804 29374
rect 20860 28642 20916 28644
rect 20860 28590 20862 28642
rect 20862 28590 20914 28642
rect 20914 28590 20916 28642
rect 20860 28588 20916 28590
rect 21084 27916 21140 27972
rect 20524 27244 20580 27300
rect 19404 25900 19460 25956
rect 19516 27132 19572 27188
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19628 25676 19684 25732
rect 19516 25394 19572 25396
rect 19516 25342 19518 25394
rect 19518 25342 19570 25394
rect 19570 25342 19572 25394
rect 19516 25340 19572 25342
rect 20300 25730 20356 25732
rect 20300 25678 20302 25730
rect 20302 25678 20354 25730
rect 20354 25678 20356 25730
rect 20300 25676 20356 25678
rect 18844 24892 18900 24948
rect 18732 23884 18788 23940
rect 18844 23772 18900 23828
rect 18956 24108 19012 24164
rect 18956 23548 19012 23604
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19292 24332 19348 24388
rect 19404 24892 19460 24948
rect 19180 24108 19236 24164
rect 19404 23996 19460 24052
rect 19180 23772 19236 23828
rect 19180 23436 19236 23492
rect 19068 23100 19124 23156
rect 18956 22652 19012 22708
rect 18620 21756 18676 21812
rect 18732 22092 18788 22148
rect 18060 19906 18116 19908
rect 18060 19854 18062 19906
rect 18062 19854 18114 19906
rect 18114 19854 18116 19906
rect 18060 19852 18116 19854
rect 18620 19852 18676 19908
rect 18284 19068 18340 19124
rect 17388 17836 17444 17892
rect 17612 17106 17668 17108
rect 17612 17054 17614 17106
rect 17614 17054 17666 17106
rect 17666 17054 17668 17106
rect 17612 17052 17668 17054
rect 17388 16940 17444 16996
rect 17388 15426 17444 15428
rect 17388 15374 17390 15426
rect 17390 15374 17442 15426
rect 17442 15374 17444 15426
rect 17388 15372 17444 15374
rect 17276 14252 17332 14308
rect 17612 13746 17668 13748
rect 17612 13694 17614 13746
rect 17614 13694 17666 13746
rect 17666 13694 17668 13746
rect 17612 13692 17668 13694
rect 17052 12796 17108 12852
rect 18060 17836 18116 17892
rect 18172 17666 18228 17668
rect 18172 17614 18174 17666
rect 18174 17614 18226 17666
rect 18226 17614 18228 17666
rect 18172 17612 18228 17614
rect 17948 16994 18004 16996
rect 17948 16942 17950 16994
rect 17950 16942 18002 16994
rect 18002 16942 18004 16994
rect 17948 16940 18004 16942
rect 18508 18226 18564 18228
rect 18508 18174 18510 18226
rect 18510 18174 18562 18226
rect 18562 18174 18564 18226
rect 18508 18172 18564 18174
rect 18844 20860 18900 20916
rect 18732 19740 18788 19796
rect 19068 20972 19124 21028
rect 18732 17890 18788 17892
rect 18732 17838 18734 17890
rect 18734 17838 18786 17890
rect 18786 17838 18788 17890
rect 18732 17836 18788 17838
rect 18620 17724 18676 17780
rect 18956 18450 19012 18452
rect 18956 18398 18958 18450
rect 18958 18398 19010 18450
rect 19010 18398 19012 18450
rect 18956 18396 19012 18398
rect 19964 24722 20020 24724
rect 19964 24670 19966 24722
rect 19966 24670 20018 24722
rect 20018 24670 20020 24722
rect 19964 24668 20020 24670
rect 19628 24332 19684 24388
rect 19628 24108 19684 24164
rect 20188 23996 20244 24052
rect 20076 23938 20132 23940
rect 20076 23886 20078 23938
rect 20078 23886 20130 23938
rect 20130 23886 20132 23938
rect 20076 23884 20132 23886
rect 19964 23772 20020 23828
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19628 23324 19684 23380
rect 19516 22316 19572 22372
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19628 21810 19684 21812
rect 19628 21758 19630 21810
rect 19630 21758 19682 21810
rect 19682 21758 19684 21810
rect 19628 21756 19684 21758
rect 20076 21756 20132 21812
rect 19404 21698 19460 21700
rect 19404 21646 19406 21698
rect 19406 21646 19458 21698
rect 19458 21646 19460 21698
rect 19404 21644 19460 21646
rect 19964 21698 20020 21700
rect 19964 21646 19966 21698
rect 19966 21646 20018 21698
rect 20018 21646 20020 21698
rect 19964 21644 20020 21646
rect 19292 21420 19348 21476
rect 20076 21420 20132 21476
rect 19628 20860 19684 20916
rect 19516 19404 19572 19460
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20748 25564 20804 25620
rect 20860 25452 20916 25508
rect 20524 23660 20580 23716
rect 20972 24668 21028 24724
rect 21868 31948 21924 32004
rect 22540 35026 22596 35028
rect 22540 34974 22542 35026
rect 22542 34974 22594 35026
rect 22594 34974 22596 35026
rect 22540 34972 22596 34974
rect 22876 36258 22932 36260
rect 22876 36206 22878 36258
rect 22878 36206 22930 36258
rect 22930 36206 22932 36258
rect 22876 36204 22932 36206
rect 23548 37212 23604 37268
rect 23212 35698 23268 35700
rect 23212 35646 23214 35698
rect 23214 35646 23266 35698
rect 23266 35646 23268 35698
rect 23212 35644 23268 35646
rect 23548 35644 23604 35700
rect 23660 36876 23716 36932
rect 24668 40796 24724 40852
rect 24892 44322 24948 44324
rect 24892 44270 24894 44322
rect 24894 44270 24946 44322
rect 24946 44270 24948 44322
rect 24892 44268 24948 44270
rect 24892 41916 24948 41972
rect 24780 40684 24836 40740
rect 24668 40626 24724 40628
rect 24668 40574 24670 40626
rect 24670 40574 24722 40626
rect 24722 40574 24724 40626
rect 24668 40572 24724 40574
rect 25116 45276 25172 45332
rect 25564 46786 25620 46788
rect 25564 46734 25566 46786
rect 25566 46734 25618 46786
rect 25618 46734 25620 46786
rect 25564 46732 25620 46734
rect 25340 45500 25396 45556
rect 25452 45276 25508 45332
rect 25116 44380 25172 44436
rect 25452 44604 25508 44660
rect 25340 44268 25396 44324
rect 25452 43372 25508 43428
rect 25228 42754 25284 42756
rect 25228 42702 25230 42754
rect 25230 42702 25282 42754
rect 25282 42702 25284 42754
rect 25228 42700 25284 42702
rect 25340 41580 25396 41636
rect 25228 40572 25284 40628
rect 25900 48018 25956 48020
rect 25900 47966 25902 48018
rect 25902 47966 25954 48018
rect 25954 47966 25956 48018
rect 25900 47964 25956 47966
rect 28476 57820 28532 57876
rect 28476 57538 28532 57540
rect 28476 57486 28478 57538
rect 28478 57486 28530 57538
rect 28530 57486 28532 57538
rect 28476 57484 28532 57486
rect 28252 55356 28308 55412
rect 28476 57148 28532 57204
rect 28588 56252 28644 56308
rect 28812 58156 28868 58212
rect 28812 56364 28868 56420
rect 28252 55074 28308 55076
rect 28252 55022 28254 55074
rect 28254 55022 28306 55074
rect 28306 55022 28308 55074
rect 28252 55020 28308 55022
rect 28476 54626 28532 54628
rect 28476 54574 28478 54626
rect 28478 54574 28530 54626
rect 28530 54574 28532 54626
rect 28476 54572 28532 54574
rect 28140 53564 28196 53620
rect 28588 53676 28644 53732
rect 28252 53506 28308 53508
rect 28252 53454 28254 53506
rect 28254 53454 28306 53506
rect 28306 53454 28308 53506
rect 28252 53452 28308 53454
rect 28028 52668 28084 52724
rect 27132 52108 27188 52164
rect 27020 49196 27076 49252
rect 27132 49756 27188 49812
rect 26684 48914 26740 48916
rect 26684 48862 26686 48914
rect 26686 48862 26738 48914
rect 26738 48862 26740 48914
rect 26684 48860 26740 48862
rect 26572 47682 26628 47684
rect 26572 47630 26574 47682
rect 26574 47630 26626 47682
rect 26626 47630 26628 47682
rect 26572 47628 26628 47630
rect 26012 47404 26068 47460
rect 25788 45724 25844 45780
rect 25900 47180 25956 47236
rect 26012 45890 26068 45892
rect 26012 45838 26014 45890
rect 26014 45838 26066 45890
rect 26066 45838 26068 45890
rect 26012 45836 26068 45838
rect 26012 45666 26068 45668
rect 26012 45614 26014 45666
rect 26014 45614 26066 45666
rect 26066 45614 26068 45666
rect 26012 45612 26068 45614
rect 25676 45276 25732 45332
rect 25900 45164 25956 45220
rect 25676 44716 25732 44772
rect 26908 47346 26964 47348
rect 26908 47294 26910 47346
rect 26910 47294 26962 47346
rect 26962 47294 26964 47346
rect 26908 47292 26964 47294
rect 26236 46620 26292 46676
rect 26796 45890 26852 45892
rect 26796 45838 26798 45890
rect 26798 45838 26850 45890
rect 26850 45838 26852 45890
rect 26796 45836 26852 45838
rect 26236 45500 26292 45556
rect 26908 45724 26964 45780
rect 26684 45500 26740 45556
rect 26796 45612 26852 45668
rect 26572 45164 26628 45220
rect 26012 44940 26068 44996
rect 25900 44716 25956 44772
rect 26236 44604 26292 44660
rect 26124 43538 26180 43540
rect 26124 43486 26126 43538
rect 26126 43486 26178 43538
rect 26178 43486 26180 43538
rect 26124 43484 26180 43486
rect 26460 44156 26516 44212
rect 28700 53116 28756 53172
rect 28588 53004 28644 53060
rect 27580 52220 27636 52276
rect 27804 52108 27860 52164
rect 28924 51996 28980 52052
rect 28028 50594 28084 50596
rect 28028 50542 28030 50594
rect 28030 50542 28082 50594
rect 28082 50542 28084 50594
rect 28028 50540 28084 50542
rect 29148 58716 29204 58772
rect 29596 58716 29652 58772
rect 29484 58658 29540 58660
rect 29484 58606 29486 58658
rect 29486 58606 29538 58658
rect 29538 58606 29540 58658
rect 29484 58604 29540 58606
rect 29596 58434 29652 58436
rect 29596 58382 29598 58434
rect 29598 58382 29650 58434
rect 29650 58382 29652 58434
rect 29596 58380 29652 58382
rect 29260 57650 29316 57652
rect 29260 57598 29262 57650
rect 29262 57598 29314 57650
rect 29314 57598 29316 57650
rect 29260 57596 29316 57598
rect 31164 59890 31220 59892
rect 31164 59838 31166 59890
rect 31166 59838 31218 59890
rect 31218 59838 31220 59890
rect 31164 59836 31220 59838
rect 32732 59836 32788 59892
rect 30044 59724 30100 59780
rect 29820 59276 29876 59332
rect 29820 59052 29876 59108
rect 30268 58828 30324 58884
rect 30156 58380 30212 58436
rect 30156 57650 30212 57652
rect 30156 57598 30158 57650
rect 30158 57598 30210 57650
rect 30210 57598 30212 57650
rect 30156 57596 30212 57598
rect 29148 57148 29204 57204
rect 29484 57484 29540 57540
rect 29148 56252 29204 56308
rect 29820 57148 29876 57204
rect 29596 56140 29652 56196
rect 29708 56476 29764 56532
rect 29932 56082 29988 56084
rect 29932 56030 29934 56082
rect 29934 56030 29986 56082
rect 29986 56030 29988 56082
rect 29932 56028 29988 56030
rect 29484 54738 29540 54740
rect 29484 54686 29486 54738
rect 29486 54686 29538 54738
rect 29538 54686 29540 54738
rect 29484 54684 29540 54686
rect 29148 54460 29204 54516
rect 29932 54460 29988 54516
rect 30380 58716 30436 58772
rect 31164 58940 31220 58996
rect 32284 59164 32340 59220
rect 32396 59778 32452 59780
rect 32396 59726 32398 59778
rect 32398 59726 32450 59778
rect 32450 59726 32452 59778
rect 32396 59724 32452 59726
rect 32172 58940 32228 58996
rect 31276 58716 31332 58772
rect 30492 56588 30548 56644
rect 32172 58380 32228 58436
rect 31388 56754 31444 56756
rect 31388 56702 31390 56754
rect 31390 56702 31442 56754
rect 31442 56702 31444 56754
rect 31388 56700 31444 56702
rect 31276 56588 31332 56644
rect 31052 56476 31108 56532
rect 30604 56140 30660 56196
rect 30156 55410 30212 55412
rect 30156 55358 30158 55410
rect 30158 55358 30210 55410
rect 30210 55358 30212 55410
rect 30156 55356 30212 55358
rect 30156 54684 30212 54740
rect 30380 54236 30436 54292
rect 29708 53506 29764 53508
rect 29708 53454 29710 53506
rect 29710 53454 29762 53506
rect 29762 53454 29764 53506
rect 29708 53452 29764 53454
rect 29260 53170 29316 53172
rect 29260 53118 29262 53170
rect 29262 53118 29314 53170
rect 29314 53118 29316 53170
rect 29260 53116 29316 53118
rect 29372 52780 29428 52836
rect 29260 52108 29316 52164
rect 29148 52050 29204 52052
rect 29148 51998 29150 52050
rect 29150 51998 29202 52050
rect 29202 51998 29204 52050
rect 29148 51996 29204 51998
rect 29708 53170 29764 53172
rect 29708 53118 29710 53170
rect 29710 53118 29762 53170
rect 29762 53118 29764 53170
rect 29708 53116 29764 53118
rect 27804 49756 27860 49812
rect 27692 49644 27748 49700
rect 29036 49586 29092 49588
rect 29036 49534 29038 49586
rect 29038 49534 29090 49586
rect 29090 49534 29092 49586
rect 29036 49532 29092 49534
rect 27244 48860 27300 48916
rect 27132 45388 27188 45444
rect 27020 45052 27076 45108
rect 26236 43372 26292 43428
rect 26796 43260 26852 43316
rect 26124 42194 26180 42196
rect 26124 42142 26126 42194
rect 26126 42142 26178 42194
rect 26178 42142 26180 42194
rect 26124 42140 26180 42142
rect 25676 41356 25732 41412
rect 25676 40514 25732 40516
rect 25676 40462 25678 40514
rect 25678 40462 25730 40514
rect 25730 40462 25732 40514
rect 25676 40460 25732 40462
rect 26012 41970 26068 41972
rect 26012 41918 26014 41970
rect 26014 41918 26066 41970
rect 26066 41918 26068 41970
rect 26012 41916 26068 41918
rect 26348 41468 26404 41524
rect 26012 40684 26068 40740
rect 24220 38444 24276 38500
rect 25228 39452 25284 39508
rect 24668 37154 24724 37156
rect 24668 37102 24670 37154
rect 24670 37102 24722 37154
rect 24722 37102 24724 37154
rect 24668 37100 24724 37102
rect 23996 36540 24052 36596
rect 24332 36370 24388 36372
rect 24332 36318 24334 36370
rect 24334 36318 24386 36370
rect 24386 36318 24388 36370
rect 24332 36316 24388 36318
rect 24444 35586 24500 35588
rect 24444 35534 24446 35586
rect 24446 35534 24498 35586
rect 24498 35534 24500 35586
rect 24444 35532 24500 35534
rect 23548 35474 23604 35476
rect 23548 35422 23550 35474
rect 23550 35422 23602 35474
rect 23602 35422 23604 35474
rect 23548 35420 23604 35422
rect 23324 34188 23380 34244
rect 22876 33906 22932 33908
rect 22876 33854 22878 33906
rect 22878 33854 22930 33906
rect 22930 33854 22932 33906
rect 22876 33852 22932 33854
rect 22316 32620 22372 32676
rect 22316 32002 22372 32004
rect 22316 31950 22318 32002
rect 22318 31950 22370 32002
rect 22370 31950 22372 32002
rect 22316 31948 22372 31950
rect 22540 31948 22596 32004
rect 21532 31778 21588 31780
rect 21532 31726 21534 31778
rect 21534 31726 21586 31778
rect 21586 31726 21588 31778
rect 21532 31724 21588 31726
rect 22092 31724 22148 31780
rect 21308 31666 21364 31668
rect 21308 31614 21310 31666
rect 21310 31614 21362 31666
rect 21362 31614 21364 31666
rect 21308 31612 21364 31614
rect 21980 31612 22036 31668
rect 21308 30828 21364 30884
rect 21420 30268 21476 30324
rect 21868 30044 21924 30100
rect 21644 29372 21700 29428
rect 21756 27916 21812 27972
rect 21196 27020 21252 27076
rect 21644 25788 21700 25844
rect 21532 25394 21588 25396
rect 21532 25342 21534 25394
rect 21534 25342 21586 25394
rect 21586 25342 21588 25394
rect 21532 25340 21588 25342
rect 21308 24668 21364 24724
rect 21084 24556 21140 24612
rect 20972 24332 21028 24388
rect 21420 23772 21476 23828
rect 20412 21644 20468 21700
rect 20636 21586 20692 21588
rect 20636 21534 20638 21586
rect 20638 21534 20690 21586
rect 20690 21534 20692 21586
rect 20636 21532 20692 21534
rect 20636 20802 20692 20804
rect 20636 20750 20638 20802
rect 20638 20750 20690 20802
rect 20690 20750 20692 20802
rect 20636 20748 20692 20750
rect 20188 20188 20244 20244
rect 20076 19404 20132 19460
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19068 18284 19124 18340
rect 18396 16716 18452 16772
rect 18956 17612 19012 17668
rect 18172 16044 18228 16100
rect 17836 14476 17892 14532
rect 17836 13020 17892 13076
rect 18396 14252 18452 14308
rect 18284 14140 18340 14196
rect 16492 11340 16548 11396
rect 16716 11676 16772 11732
rect 16828 11618 16884 11620
rect 16828 11566 16830 11618
rect 16830 11566 16882 11618
rect 16882 11566 16884 11618
rect 16828 11564 16884 11566
rect 17724 12124 17780 12180
rect 17500 12012 17556 12068
rect 16604 11116 16660 11172
rect 16156 10668 16212 10724
rect 16044 10498 16100 10500
rect 16044 10446 16046 10498
rect 16046 10446 16098 10498
rect 16098 10446 16100 10498
rect 16044 10444 16100 10446
rect 16380 9772 16436 9828
rect 16492 9996 16548 10052
rect 15708 9436 15764 9492
rect 15708 8540 15764 8596
rect 15596 6972 15652 7028
rect 16044 8204 16100 8260
rect 15932 8034 15988 8036
rect 15932 7982 15934 8034
rect 15934 7982 15986 8034
rect 15986 7982 15988 8034
rect 15932 7980 15988 7982
rect 16156 8876 16212 8932
rect 15932 7474 15988 7476
rect 15932 7422 15934 7474
rect 15934 7422 15986 7474
rect 15986 7422 15988 7474
rect 15932 7420 15988 7422
rect 15820 6690 15876 6692
rect 15820 6638 15822 6690
rect 15822 6638 15874 6690
rect 15874 6638 15876 6690
rect 15820 6636 15876 6638
rect 16044 6076 16100 6132
rect 16492 8876 16548 8932
rect 16380 8316 16436 8372
rect 16492 8652 16548 8708
rect 16268 6690 16324 6692
rect 16268 6638 16270 6690
rect 16270 6638 16322 6690
rect 16322 6638 16324 6690
rect 16268 6636 16324 6638
rect 17052 10220 17108 10276
rect 16940 9996 16996 10052
rect 16716 8316 16772 8372
rect 16940 9772 16996 9828
rect 17612 11564 17668 11620
rect 17948 12012 18004 12068
rect 17836 11676 17892 11732
rect 20636 20076 20692 20132
rect 20524 20018 20580 20020
rect 20524 19966 20526 20018
rect 20526 19966 20578 20018
rect 20578 19966 20580 20018
rect 20524 19964 20580 19966
rect 20300 18396 20356 18452
rect 20524 18450 20580 18452
rect 20524 18398 20526 18450
rect 20526 18398 20578 18450
rect 20578 18398 20580 18450
rect 20524 18396 20580 18398
rect 18732 15036 18788 15092
rect 18620 14700 18676 14756
rect 18732 14140 18788 14196
rect 18956 14364 19012 14420
rect 18620 13858 18676 13860
rect 18620 13806 18622 13858
rect 18622 13806 18674 13858
rect 18674 13806 18676 13858
rect 18620 13804 18676 13806
rect 19516 16156 19572 16212
rect 19292 15036 19348 15092
rect 19516 14924 19572 14980
rect 19068 13692 19124 13748
rect 20076 17778 20132 17780
rect 20076 17726 20078 17778
rect 20078 17726 20130 17778
rect 20130 17726 20132 17778
rect 20076 17724 20132 17726
rect 20188 17666 20244 17668
rect 20188 17614 20190 17666
rect 20190 17614 20242 17666
rect 20242 17614 20244 17666
rect 20188 17612 20244 17614
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20524 17836 20580 17892
rect 20412 16994 20468 16996
rect 20412 16942 20414 16994
rect 20414 16942 20466 16994
rect 20466 16942 20468 16994
rect 20412 16940 20468 16942
rect 20636 17724 20692 17780
rect 20972 21698 21028 21700
rect 20972 21646 20974 21698
rect 20974 21646 21026 21698
rect 21026 21646 21028 21698
rect 20972 21644 21028 21646
rect 21084 21532 21140 21588
rect 21532 23660 21588 23716
rect 21420 21980 21476 22036
rect 21308 21756 21364 21812
rect 21420 20018 21476 20020
rect 21420 19966 21422 20018
rect 21422 19966 21474 20018
rect 21474 19966 21476 20018
rect 21420 19964 21476 19966
rect 21420 19458 21476 19460
rect 21420 19406 21422 19458
rect 21422 19406 21474 19458
rect 21474 19406 21476 19458
rect 21420 19404 21476 19406
rect 21644 22428 21700 22484
rect 22428 30882 22484 30884
rect 22428 30830 22430 30882
rect 22430 30830 22482 30882
rect 22482 30830 22484 30882
rect 22428 30828 22484 30830
rect 22876 32674 22932 32676
rect 22876 32622 22878 32674
rect 22878 32622 22930 32674
rect 22930 32622 22932 32674
rect 22876 32620 22932 32622
rect 22764 31778 22820 31780
rect 22764 31726 22766 31778
rect 22766 31726 22818 31778
rect 22818 31726 22820 31778
rect 22764 31724 22820 31726
rect 23436 34130 23492 34132
rect 23436 34078 23438 34130
rect 23438 34078 23490 34130
rect 23490 34078 23492 34130
rect 23436 34076 23492 34078
rect 23660 33906 23716 33908
rect 23660 33854 23662 33906
rect 23662 33854 23714 33906
rect 23714 33854 23716 33906
rect 23660 33852 23716 33854
rect 23436 33628 23492 33684
rect 23212 31836 23268 31892
rect 22204 29932 22260 29988
rect 23100 31500 23156 31556
rect 23772 32060 23828 32116
rect 23548 31666 23604 31668
rect 23548 31614 23550 31666
rect 23550 31614 23602 31666
rect 23602 31614 23604 31666
rect 23548 31612 23604 31614
rect 23212 31164 23268 31220
rect 22316 29148 22372 29204
rect 23100 30940 23156 30996
rect 22204 29036 22260 29092
rect 23212 30716 23268 30772
rect 23212 30268 23268 30324
rect 22652 29372 22708 29428
rect 22428 27074 22484 27076
rect 22428 27022 22430 27074
rect 22430 27022 22482 27074
rect 22482 27022 22484 27074
rect 22428 27020 22484 27022
rect 22764 27858 22820 27860
rect 22764 27806 22766 27858
rect 22766 27806 22818 27858
rect 22818 27806 22820 27858
rect 22764 27804 22820 27806
rect 22204 26290 22260 26292
rect 22204 26238 22206 26290
rect 22206 26238 22258 26290
rect 22258 26238 22260 26290
rect 22204 26236 22260 26238
rect 22092 25564 22148 25620
rect 21868 25506 21924 25508
rect 21868 25454 21870 25506
rect 21870 25454 21922 25506
rect 21922 25454 21924 25506
rect 21868 25452 21924 25454
rect 22316 25564 22372 25620
rect 22540 25452 22596 25508
rect 22204 25394 22260 25396
rect 22204 25342 22206 25394
rect 22206 25342 22258 25394
rect 22258 25342 22260 25394
rect 22204 25340 22260 25342
rect 21868 23660 21924 23716
rect 21980 23548 22036 23604
rect 21756 22316 21812 22372
rect 21868 21980 21924 22036
rect 21980 22092 22036 22148
rect 21644 21420 21700 21476
rect 21980 21308 22036 21364
rect 21756 20188 21812 20244
rect 21756 18284 21812 18340
rect 22764 26348 22820 26404
rect 22764 25228 22820 25284
rect 23436 30716 23492 30772
rect 26124 40012 26180 40068
rect 25564 38892 25620 38948
rect 25788 38780 25844 38836
rect 25676 38722 25732 38724
rect 25676 38670 25678 38722
rect 25678 38670 25730 38722
rect 25730 38670 25732 38722
rect 25676 38668 25732 38670
rect 25564 38444 25620 38500
rect 25340 37772 25396 37828
rect 25676 38332 25732 38388
rect 25452 36652 25508 36708
rect 25228 35698 25284 35700
rect 25228 35646 25230 35698
rect 25230 35646 25282 35698
rect 25282 35646 25284 35698
rect 25228 35644 25284 35646
rect 24556 34188 24612 34244
rect 24332 34018 24388 34020
rect 24332 33966 24334 34018
rect 24334 33966 24386 34018
rect 24386 33966 24388 34018
rect 24332 33964 24388 33966
rect 24108 33068 24164 33124
rect 24444 33740 24500 33796
rect 24780 33628 24836 33684
rect 24668 31948 24724 32004
rect 24332 31836 24388 31892
rect 23996 31778 24052 31780
rect 23996 31726 23998 31778
rect 23998 31726 24050 31778
rect 24050 31726 24052 31778
rect 23996 31724 24052 31726
rect 24556 31666 24612 31668
rect 24556 31614 24558 31666
rect 24558 31614 24610 31666
rect 24610 31614 24612 31666
rect 24556 31612 24612 31614
rect 23772 30940 23828 30996
rect 23660 30882 23716 30884
rect 23660 30830 23662 30882
rect 23662 30830 23714 30882
rect 23714 30830 23716 30882
rect 23660 30828 23716 30830
rect 23548 30492 23604 30548
rect 23436 27970 23492 27972
rect 23436 27918 23438 27970
rect 23438 27918 23490 27970
rect 23490 27918 23492 27970
rect 23436 27916 23492 27918
rect 23660 27468 23716 27524
rect 23660 27244 23716 27300
rect 22876 24780 22932 24836
rect 23324 27020 23380 27076
rect 23324 26402 23380 26404
rect 23324 26350 23326 26402
rect 23326 26350 23378 26402
rect 23378 26350 23380 26402
rect 23324 26348 23380 26350
rect 24332 31500 24388 31556
rect 23996 30380 24052 30436
rect 23884 30098 23940 30100
rect 23884 30046 23886 30098
rect 23886 30046 23938 30098
rect 23938 30046 23940 30098
rect 23884 30044 23940 30046
rect 23884 29820 23940 29876
rect 23996 29426 24052 29428
rect 23996 29374 23998 29426
rect 23998 29374 24050 29426
rect 24050 29374 24052 29426
rect 23996 29372 24052 29374
rect 24332 29596 24388 29652
rect 24220 29426 24276 29428
rect 24220 29374 24222 29426
rect 24222 29374 24274 29426
rect 24274 29374 24276 29426
rect 24220 29372 24276 29374
rect 23772 26124 23828 26180
rect 24220 27858 24276 27860
rect 24220 27806 24222 27858
rect 24222 27806 24274 27858
rect 24274 27806 24276 27858
rect 24220 27804 24276 27806
rect 24332 27692 24388 27748
rect 24556 31218 24612 31220
rect 24556 31166 24558 31218
rect 24558 31166 24610 31218
rect 24610 31166 24612 31218
rect 24556 31164 24612 31166
rect 24668 30994 24724 30996
rect 24668 30942 24670 30994
rect 24670 30942 24722 30994
rect 24722 30942 24724 30994
rect 24668 30940 24724 30942
rect 24668 30492 24724 30548
rect 24556 30210 24612 30212
rect 24556 30158 24558 30210
rect 24558 30158 24610 30210
rect 24610 30158 24612 30210
rect 24556 30156 24612 30158
rect 24668 29260 24724 29316
rect 24556 28754 24612 28756
rect 24556 28702 24558 28754
rect 24558 28702 24610 28754
rect 24610 28702 24612 28754
rect 24556 28700 24612 28702
rect 24668 27970 24724 27972
rect 24668 27918 24670 27970
rect 24670 27918 24722 27970
rect 24722 27918 24724 27970
rect 24668 27916 24724 27918
rect 24444 27356 24500 27412
rect 24220 26236 24276 26292
rect 25004 33628 25060 33684
rect 25900 38892 25956 38948
rect 25676 36204 25732 36260
rect 26124 39228 26180 39284
rect 26908 42812 26964 42868
rect 27468 46956 27524 47012
rect 27468 46060 27524 46116
rect 27804 46674 27860 46676
rect 27804 46622 27806 46674
rect 27806 46622 27858 46674
rect 27858 46622 27860 46674
rect 27804 46620 27860 46622
rect 27916 46172 27972 46228
rect 28028 48300 28084 48356
rect 28252 48188 28308 48244
rect 28028 47068 28084 47124
rect 28140 47516 28196 47572
rect 29036 48242 29092 48244
rect 29036 48190 29038 48242
rect 29038 48190 29090 48242
rect 29090 48190 29092 48242
rect 29036 48188 29092 48190
rect 28476 47964 28532 48020
rect 28364 47852 28420 47908
rect 28700 47404 28756 47460
rect 27804 44380 27860 44436
rect 27804 44210 27860 44212
rect 27804 44158 27806 44210
rect 27806 44158 27858 44210
rect 27858 44158 27860 44210
rect 27804 44156 27860 44158
rect 28252 45164 28308 45220
rect 27804 43484 27860 43540
rect 27580 43260 27636 43316
rect 27132 42252 27188 42308
rect 27244 42364 27300 42420
rect 27020 42140 27076 42196
rect 27244 42028 27300 42084
rect 27356 41692 27412 41748
rect 27468 42476 27524 42532
rect 26572 41356 26628 41412
rect 27020 40572 27076 40628
rect 26460 39452 26516 39508
rect 26796 39228 26852 39284
rect 26908 38780 26964 38836
rect 26124 38556 26180 38612
rect 26796 37660 26852 37716
rect 26236 37212 26292 37268
rect 26908 37436 26964 37492
rect 27580 40460 27636 40516
rect 28028 43372 28084 43428
rect 27916 43260 27972 43316
rect 27916 42476 27972 42532
rect 28700 44098 28756 44100
rect 28700 44046 28702 44098
rect 28702 44046 28754 44098
rect 28754 44046 28756 44098
rect 28700 44044 28756 44046
rect 28364 43426 28420 43428
rect 28364 43374 28366 43426
rect 28366 43374 28418 43426
rect 28418 43374 28420 43426
rect 28364 43372 28420 43374
rect 27916 42082 27972 42084
rect 27916 42030 27918 42082
rect 27918 42030 27970 42082
rect 27970 42030 27972 42082
rect 27916 42028 27972 42030
rect 28476 42530 28532 42532
rect 28476 42478 28478 42530
rect 28478 42478 28530 42530
rect 28530 42478 28532 42530
rect 28476 42476 28532 42478
rect 28924 45836 28980 45892
rect 29148 47180 29204 47236
rect 29708 52892 29764 52948
rect 30380 53452 30436 53508
rect 30156 52834 30212 52836
rect 30156 52782 30158 52834
rect 30158 52782 30210 52834
rect 30210 52782 30212 52834
rect 30156 52780 30212 52782
rect 30716 56364 30772 56420
rect 31276 56364 31332 56420
rect 30828 55692 30884 55748
rect 30716 55468 30772 55524
rect 31052 55522 31108 55524
rect 31052 55470 31054 55522
rect 31054 55470 31106 55522
rect 31106 55470 31108 55522
rect 31052 55468 31108 55470
rect 31500 55468 31556 55524
rect 31612 56476 31668 56532
rect 30604 55020 30660 55076
rect 30716 55298 30772 55300
rect 30716 55246 30718 55298
rect 30718 55246 30770 55298
rect 30770 55246 30772 55298
rect 30716 55244 30772 55246
rect 30604 54572 30660 54628
rect 30492 53228 30548 53284
rect 30604 53676 30660 53732
rect 30492 52946 30548 52948
rect 30492 52894 30494 52946
rect 30494 52894 30546 52946
rect 30546 52894 30548 52946
rect 30492 52892 30548 52894
rect 30380 52220 30436 52276
rect 29596 49196 29652 49252
rect 30156 52108 30212 52164
rect 30268 52050 30324 52052
rect 30268 51998 30270 52050
rect 30270 51998 30322 52050
rect 30322 51998 30324 52050
rect 30268 51996 30324 51998
rect 31276 54514 31332 54516
rect 31276 54462 31278 54514
rect 31278 54462 31330 54514
rect 31330 54462 31332 54514
rect 31276 54460 31332 54462
rect 30940 54236 30996 54292
rect 30828 54124 30884 54180
rect 30828 53954 30884 53956
rect 30828 53902 30830 53954
rect 30830 53902 30882 53954
rect 30882 53902 30884 53954
rect 30828 53900 30884 53902
rect 31276 53954 31332 53956
rect 31276 53902 31278 53954
rect 31278 53902 31330 53954
rect 31330 53902 31332 53954
rect 31276 53900 31332 53902
rect 30940 53228 30996 53284
rect 31612 54460 31668 54516
rect 32620 58716 32676 58772
rect 32508 58380 32564 58436
rect 33068 59890 33124 59892
rect 33068 59838 33070 59890
rect 33070 59838 33122 59890
rect 33122 59838 33124 59890
rect 33068 59836 33124 59838
rect 47740 60172 47796 60228
rect 33180 59778 33236 59780
rect 33180 59726 33182 59778
rect 33182 59726 33234 59778
rect 33234 59726 33236 59778
rect 33180 59724 33236 59726
rect 33740 59612 33796 59668
rect 33180 58994 33236 58996
rect 33180 58942 33182 58994
rect 33182 58942 33234 58994
rect 33234 58942 33236 58994
rect 33180 58940 33236 58942
rect 33516 58716 33572 58772
rect 34188 59330 34244 59332
rect 34188 59278 34190 59330
rect 34190 59278 34242 59330
rect 34242 59278 34244 59330
rect 34188 59276 34244 59278
rect 32844 57596 32900 57652
rect 32060 56700 32116 56756
rect 32396 56588 32452 56644
rect 32172 56194 32228 56196
rect 32172 56142 32174 56194
rect 32174 56142 32226 56194
rect 32226 56142 32228 56194
rect 32172 56140 32228 56142
rect 31948 56082 32004 56084
rect 31948 56030 31950 56082
rect 31950 56030 32002 56082
rect 32002 56030 32004 56082
rect 31948 56028 32004 56030
rect 32172 55916 32228 55972
rect 31948 55186 32004 55188
rect 31948 55134 31950 55186
rect 31950 55134 32002 55186
rect 32002 55134 32004 55186
rect 31948 55132 32004 55134
rect 32732 57148 32788 57204
rect 33740 57650 33796 57652
rect 33740 57598 33742 57650
rect 33742 57598 33794 57650
rect 33794 57598 33796 57650
rect 33740 57596 33796 57598
rect 34076 59052 34132 59108
rect 32620 55468 32676 55524
rect 33068 56588 33124 56644
rect 32732 55692 32788 55748
rect 33068 55356 33124 55412
rect 32620 55298 32676 55300
rect 32620 55246 32622 55298
rect 32622 55246 32674 55298
rect 32674 55246 32676 55298
rect 32620 55244 32676 55246
rect 33292 55916 33348 55972
rect 33180 55244 33236 55300
rect 33292 55356 33348 55412
rect 32508 54796 32564 54852
rect 32172 54626 32228 54628
rect 32172 54574 32174 54626
rect 32174 54574 32226 54626
rect 32226 54574 32228 54626
rect 32172 54572 32228 54574
rect 31836 54348 31892 54404
rect 31948 54124 32004 54180
rect 31724 53676 31780 53732
rect 33180 53788 33236 53844
rect 31724 53506 31780 53508
rect 31724 53454 31726 53506
rect 31726 53454 31778 53506
rect 31778 53454 31780 53506
rect 31724 53452 31780 53454
rect 31276 52780 31332 52836
rect 30604 52332 30660 52388
rect 30492 51548 30548 51604
rect 29932 50540 29988 50596
rect 30156 50652 30212 50708
rect 29820 50428 29876 50484
rect 29932 50092 29988 50148
rect 29820 49698 29876 49700
rect 29820 49646 29822 49698
rect 29822 49646 29874 49698
rect 29874 49646 29876 49698
rect 29820 49644 29876 49646
rect 29708 49532 29764 49588
rect 29596 48748 29652 48804
rect 30044 49026 30100 49028
rect 30044 48974 30046 49026
rect 30046 48974 30098 49026
rect 30098 48974 30100 49026
rect 30044 48972 30100 48974
rect 29932 48636 29988 48692
rect 29820 48412 29876 48468
rect 29596 48300 29652 48356
rect 29372 47292 29428 47348
rect 29820 47852 29876 47908
rect 32620 53676 32676 53732
rect 32396 53618 32452 53620
rect 32396 53566 32398 53618
rect 32398 53566 32450 53618
rect 32450 53566 32452 53618
rect 32396 53564 32452 53566
rect 32508 53506 32564 53508
rect 32508 53454 32510 53506
rect 32510 53454 32562 53506
rect 32562 53454 32564 53506
rect 32508 53452 32564 53454
rect 31948 52780 32004 52836
rect 31612 52722 31668 52724
rect 31612 52670 31614 52722
rect 31614 52670 31666 52722
rect 31666 52670 31668 52722
rect 31612 52668 31668 52670
rect 31612 52332 31668 52388
rect 30492 50876 30548 50932
rect 31948 52220 32004 52276
rect 31836 52050 31892 52052
rect 31836 51998 31838 52050
rect 31838 51998 31890 52050
rect 31890 51998 31892 52050
rect 31836 51996 31892 51998
rect 30940 50594 30996 50596
rect 30940 50542 30942 50594
rect 30942 50542 30994 50594
rect 30994 50542 30996 50594
rect 30940 50540 30996 50542
rect 30828 50092 30884 50148
rect 31164 50092 31220 50148
rect 30380 49868 30436 49924
rect 30940 49250 30996 49252
rect 30940 49198 30942 49250
rect 30942 49198 30994 49250
rect 30994 49198 30996 49250
rect 30940 49196 30996 49198
rect 30604 48972 30660 49028
rect 30604 48354 30660 48356
rect 30604 48302 30606 48354
rect 30606 48302 30658 48354
rect 30658 48302 30660 48354
rect 30604 48300 30660 48302
rect 30380 48076 30436 48132
rect 31052 48748 31108 48804
rect 30044 47404 30100 47460
rect 30604 47516 30660 47572
rect 31500 50540 31556 50596
rect 31500 49868 31556 49924
rect 31724 50428 31780 50484
rect 32172 52162 32228 52164
rect 32172 52110 32174 52162
rect 32174 52110 32226 52162
rect 32226 52110 32228 52162
rect 32172 52108 32228 52110
rect 32396 52780 32452 52836
rect 32172 51378 32228 51380
rect 32172 51326 32174 51378
rect 32174 51326 32226 51378
rect 32226 51326 32228 51378
rect 32172 51324 32228 51326
rect 32060 50764 32116 50820
rect 31948 49644 32004 49700
rect 31836 49532 31892 49588
rect 31836 49196 31892 49252
rect 31052 47404 31108 47460
rect 29708 47292 29764 47348
rect 30940 46956 30996 47012
rect 29484 45890 29540 45892
rect 29484 45838 29486 45890
rect 29486 45838 29538 45890
rect 29538 45838 29540 45890
rect 29484 45836 29540 45838
rect 29932 46674 29988 46676
rect 29932 46622 29934 46674
rect 29934 46622 29986 46674
rect 29986 46622 29988 46674
rect 29932 46620 29988 46622
rect 29932 45836 29988 45892
rect 30380 46172 30436 46228
rect 30268 45500 30324 45556
rect 29260 45388 29316 45444
rect 29484 45388 29540 45444
rect 29036 44380 29092 44436
rect 28812 42588 28868 42644
rect 29036 44044 29092 44100
rect 28140 41692 28196 41748
rect 27356 40290 27412 40292
rect 27356 40238 27358 40290
rect 27358 40238 27410 40290
rect 27410 40238 27412 40290
rect 27356 40236 27412 40238
rect 27468 39618 27524 39620
rect 27468 39566 27470 39618
rect 27470 39566 27522 39618
rect 27522 39566 27524 39618
rect 27468 39564 27524 39566
rect 27356 39506 27412 39508
rect 27356 39454 27358 39506
rect 27358 39454 27410 39506
rect 27410 39454 27412 39506
rect 27356 39452 27412 39454
rect 27244 37884 27300 37940
rect 27132 37548 27188 37604
rect 26684 37042 26740 37044
rect 26684 36990 26686 37042
rect 26686 36990 26738 37042
rect 26738 36990 26740 37042
rect 26684 36988 26740 36990
rect 26572 36876 26628 36932
rect 26572 34972 26628 35028
rect 25676 34188 25732 34244
rect 25788 33964 25844 34020
rect 25004 33122 25060 33124
rect 25004 33070 25006 33122
rect 25006 33070 25058 33122
rect 25058 33070 25060 33122
rect 25004 33068 25060 33070
rect 25228 32620 25284 32676
rect 25228 30322 25284 30324
rect 25228 30270 25230 30322
rect 25230 30270 25282 30322
rect 25282 30270 25284 30322
rect 25228 30268 25284 30270
rect 25564 31836 25620 31892
rect 25788 32732 25844 32788
rect 26012 33234 26068 33236
rect 26012 33182 26014 33234
rect 26014 33182 26066 33234
rect 26066 33182 26068 33234
rect 26012 33180 26068 33182
rect 26012 32060 26068 32116
rect 26460 33628 26516 33684
rect 26684 33404 26740 33460
rect 26236 31836 26292 31892
rect 25900 31666 25956 31668
rect 25900 31614 25902 31666
rect 25902 31614 25954 31666
rect 25954 31614 25956 31666
rect 25900 31612 25956 31614
rect 26012 31500 26068 31556
rect 25676 30770 25732 30772
rect 25676 30718 25678 30770
rect 25678 30718 25730 30770
rect 25730 30718 25732 30770
rect 25676 30716 25732 30718
rect 25452 30268 25508 30324
rect 25004 29372 25060 29428
rect 25564 30156 25620 30212
rect 25564 29708 25620 29764
rect 25564 29372 25620 29428
rect 26012 30268 26068 30324
rect 26236 30044 26292 30100
rect 26348 29372 26404 29428
rect 26124 29036 26180 29092
rect 26236 28700 26292 28756
rect 26124 28588 26180 28644
rect 25676 28476 25732 28532
rect 25452 27804 25508 27860
rect 25228 27132 25284 27188
rect 22428 23996 22484 24052
rect 22988 24108 23044 24164
rect 22876 23772 22932 23828
rect 22428 22370 22484 22372
rect 22428 22318 22430 22370
rect 22430 22318 22482 22370
rect 22482 22318 22484 22370
rect 22428 22316 22484 22318
rect 22316 22258 22372 22260
rect 22316 22206 22318 22258
rect 22318 22206 22370 22258
rect 22370 22206 22372 22258
rect 22316 22204 22372 22206
rect 22316 21586 22372 21588
rect 22316 21534 22318 21586
rect 22318 21534 22370 21586
rect 22370 21534 22372 21586
rect 22316 21532 22372 21534
rect 23100 23996 23156 24052
rect 23324 23996 23380 24052
rect 23100 23548 23156 23604
rect 23660 24722 23716 24724
rect 23660 24670 23662 24722
rect 23662 24670 23714 24722
rect 23714 24670 23716 24722
rect 23660 24668 23716 24670
rect 23660 24444 23716 24500
rect 23660 23996 23716 24052
rect 23324 23660 23380 23716
rect 23548 23772 23604 23828
rect 23324 23436 23380 23492
rect 23212 23154 23268 23156
rect 23212 23102 23214 23154
rect 23214 23102 23266 23154
rect 23266 23102 23268 23154
rect 23212 23100 23268 23102
rect 23324 22316 23380 22372
rect 23884 23548 23940 23604
rect 23100 21756 23156 21812
rect 22876 21644 22932 21700
rect 23436 21644 23492 21700
rect 22428 21084 22484 21140
rect 22092 20130 22148 20132
rect 22092 20078 22094 20130
rect 22094 20078 22146 20130
rect 22146 20078 22148 20130
rect 22092 20076 22148 20078
rect 21868 19964 21924 20020
rect 22316 19122 22372 19124
rect 22316 19070 22318 19122
rect 22318 19070 22370 19122
rect 22370 19070 22372 19122
rect 22316 19068 22372 19070
rect 22428 18562 22484 18564
rect 22428 18510 22430 18562
rect 22430 18510 22482 18562
rect 22482 18510 22484 18562
rect 22428 18508 22484 18510
rect 21980 18396 22036 18452
rect 22204 18450 22260 18452
rect 22204 18398 22206 18450
rect 22206 18398 22258 18450
rect 22258 18398 22260 18450
rect 22204 18396 22260 18398
rect 20636 16210 20692 16212
rect 20636 16158 20638 16210
rect 20638 16158 20690 16210
rect 20690 16158 20692 16210
rect 20636 16156 20692 16158
rect 20300 16098 20356 16100
rect 20300 16046 20302 16098
rect 20302 16046 20354 16098
rect 20354 16046 20356 16098
rect 20300 16044 20356 16046
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20524 15260 20580 15316
rect 20076 14924 20132 14980
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19628 13356 19684 13412
rect 19740 13244 19796 13300
rect 20412 13132 20468 13188
rect 17612 10722 17668 10724
rect 17612 10670 17614 10722
rect 17614 10670 17666 10722
rect 17666 10670 17668 10722
rect 17612 10668 17668 10670
rect 17164 9548 17220 9604
rect 17500 10220 17556 10276
rect 17388 8258 17444 8260
rect 17388 8206 17390 8258
rect 17390 8206 17442 8258
rect 17442 8206 17444 8258
rect 17388 8204 17444 8206
rect 17388 7644 17444 7700
rect 17948 11394 18004 11396
rect 17948 11342 17950 11394
rect 17950 11342 18002 11394
rect 18002 11342 18004 11394
rect 17948 11340 18004 11342
rect 17612 7644 17668 7700
rect 17500 7084 17556 7140
rect 16492 6076 16548 6132
rect 17500 6466 17556 6468
rect 17500 6414 17502 6466
rect 17502 6414 17554 6466
rect 17554 6414 17556 6466
rect 17500 6412 17556 6414
rect 16828 6130 16884 6132
rect 16828 6078 16830 6130
rect 16830 6078 16882 6130
rect 16882 6078 16884 6130
rect 16828 6076 16884 6078
rect 18732 12684 18788 12740
rect 18508 12236 18564 12292
rect 18284 10444 18340 10500
rect 18620 11004 18676 11060
rect 18060 9772 18116 9828
rect 18732 10332 18788 10388
rect 18060 9212 18116 9268
rect 19516 12850 19572 12852
rect 19516 12798 19518 12850
rect 19518 12798 19570 12850
rect 19570 12798 19572 12850
rect 19516 12796 19572 12798
rect 20188 12684 20244 12740
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 18956 12124 19012 12180
rect 21644 16940 21700 16996
rect 21532 16828 21588 16884
rect 21308 16098 21364 16100
rect 21308 16046 21310 16098
rect 21310 16046 21362 16098
rect 21362 16046 21364 16098
rect 21308 16044 21364 16046
rect 21868 16770 21924 16772
rect 21868 16718 21870 16770
rect 21870 16718 21922 16770
rect 21922 16718 21924 16770
rect 21868 16716 21924 16718
rect 21868 15820 21924 15876
rect 23436 21420 23492 21476
rect 23772 21308 23828 21364
rect 23324 20188 23380 20244
rect 23436 20300 23492 20356
rect 23660 19010 23716 19012
rect 23660 18958 23662 19010
rect 23662 18958 23714 19010
rect 23714 18958 23716 19010
rect 23660 18956 23716 18958
rect 23212 16940 23268 16996
rect 22764 16716 22820 16772
rect 22764 16268 22820 16324
rect 21980 16156 22036 16212
rect 20636 14476 20692 14532
rect 20636 13804 20692 13860
rect 21084 12908 21140 12964
rect 20524 12684 20580 12740
rect 18956 11282 19012 11284
rect 18956 11230 18958 11282
rect 18958 11230 19010 11282
rect 19010 11230 19012 11282
rect 18956 11228 19012 11230
rect 19292 10444 19348 10500
rect 18956 9996 19012 10052
rect 19292 9826 19348 9828
rect 19292 9774 19294 9826
rect 19294 9774 19346 9826
rect 19346 9774 19348 9826
rect 19292 9772 19348 9774
rect 19516 11394 19572 11396
rect 19516 11342 19518 11394
rect 19518 11342 19570 11394
rect 19570 11342 19572 11394
rect 19516 11340 19572 11342
rect 20076 12178 20132 12180
rect 20076 12126 20078 12178
rect 20078 12126 20130 12178
rect 20130 12126 20132 12178
rect 20076 12124 20132 12126
rect 20300 12236 20356 12292
rect 20188 11340 20244 11396
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19628 10780 19684 10836
rect 19516 10332 19572 10388
rect 19740 10220 19796 10276
rect 18844 9100 18900 9156
rect 19068 8988 19124 9044
rect 18620 8540 18676 8596
rect 17948 8316 18004 8372
rect 18732 7644 18788 7700
rect 17836 6636 17892 6692
rect 18956 6636 19012 6692
rect 16716 5852 16772 5908
rect 16380 5794 16436 5796
rect 16380 5742 16382 5794
rect 16382 5742 16434 5794
rect 16434 5742 16436 5794
rect 16380 5740 16436 5742
rect 19740 9548 19796 9604
rect 20860 12236 20916 12292
rect 20748 12178 20804 12180
rect 20748 12126 20750 12178
rect 20750 12126 20802 12178
rect 20802 12126 20804 12178
rect 20748 12124 20804 12126
rect 20524 11564 20580 11620
rect 20636 11170 20692 11172
rect 20636 11118 20638 11170
rect 20638 11118 20690 11170
rect 20690 11118 20692 11170
rect 20636 11116 20692 11118
rect 20300 9996 20356 10052
rect 20412 9660 20468 9716
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19740 9042 19796 9044
rect 19740 8990 19742 9042
rect 19742 8990 19794 9042
rect 19794 8990 19796 9042
rect 19740 8988 19796 8990
rect 20300 9548 20356 9604
rect 19964 8988 20020 9044
rect 20412 9100 20468 9156
rect 20636 9772 20692 9828
rect 20636 8988 20692 9044
rect 20860 9212 20916 9268
rect 21308 14812 21364 14868
rect 21420 14476 21476 14532
rect 21420 14306 21476 14308
rect 21420 14254 21422 14306
rect 21422 14254 21474 14306
rect 21474 14254 21476 14306
rect 21420 14252 21476 14254
rect 21420 13692 21476 13748
rect 21308 13244 21364 13300
rect 21868 15148 21924 15204
rect 22092 15036 22148 15092
rect 22204 14924 22260 14980
rect 21532 13634 21588 13636
rect 21532 13582 21534 13634
rect 21534 13582 21586 13634
rect 21586 13582 21588 13634
rect 21532 13580 21588 13582
rect 21756 13020 21812 13076
rect 21644 12796 21700 12852
rect 21308 12684 21364 12740
rect 21196 11004 21252 11060
rect 21308 10220 21364 10276
rect 22540 15820 22596 15876
rect 22652 15148 22708 15204
rect 24108 23660 24164 23716
rect 24108 23324 24164 23380
rect 24892 26124 24948 26180
rect 24668 25900 24724 25956
rect 24556 25564 24612 25620
rect 24556 25228 24612 25284
rect 24332 24556 24388 24612
rect 24332 24050 24388 24052
rect 24332 23998 24334 24050
rect 24334 23998 24386 24050
rect 24386 23998 24388 24050
rect 24332 23996 24388 23998
rect 24444 23938 24500 23940
rect 24444 23886 24446 23938
rect 24446 23886 24498 23938
rect 24498 23886 24500 23938
rect 24444 23884 24500 23886
rect 24668 24108 24724 24164
rect 24220 21644 24276 21700
rect 24892 23826 24948 23828
rect 24892 23774 24894 23826
rect 24894 23774 24946 23826
rect 24946 23774 24948 23826
rect 24892 23772 24948 23774
rect 24780 23324 24836 23380
rect 24556 23154 24612 23156
rect 24556 23102 24558 23154
rect 24558 23102 24610 23154
rect 24610 23102 24612 23154
rect 24556 23100 24612 23102
rect 24444 22316 24500 22372
rect 25340 27074 25396 27076
rect 25340 27022 25342 27074
rect 25342 27022 25394 27074
rect 25394 27022 25396 27074
rect 25340 27020 25396 27022
rect 26012 27970 26068 27972
rect 26012 27918 26014 27970
rect 26014 27918 26066 27970
rect 26066 27918 26068 27970
rect 26012 27916 26068 27918
rect 25676 27692 25732 27748
rect 26236 27916 26292 27972
rect 26348 27692 26404 27748
rect 26124 27356 26180 27412
rect 27020 36540 27076 36596
rect 28140 41132 28196 41188
rect 27916 40290 27972 40292
rect 27916 40238 27918 40290
rect 27918 40238 27970 40290
rect 27970 40238 27972 40290
rect 27916 40236 27972 40238
rect 28252 39900 28308 39956
rect 28252 39452 28308 39508
rect 27692 38332 27748 38388
rect 28140 38332 28196 38388
rect 28252 37996 28308 38052
rect 27692 37660 27748 37716
rect 27692 36988 27748 37044
rect 28476 41186 28532 41188
rect 28476 41134 28478 41186
rect 28478 41134 28530 41186
rect 28530 41134 28532 41186
rect 28476 41132 28532 41134
rect 28588 40796 28644 40852
rect 28700 40684 28756 40740
rect 28588 39900 28644 39956
rect 28476 39842 28532 39844
rect 28476 39790 28478 39842
rect 28478 39790 28530 39842
rect 28530 39790 28532 39842
rect 28476 39788 28532 39790
rect 28476 38220 28532 38276
rect 27804 37100 27860 37156
rect 27132 34636 27188 34692
rect 27356 34748 27412 34804
rect 27916 36594 27972 36596
rect 27916 36542 27918 36594
rect 27918 36542 27970 36594
rect 27970 36542 27972 36594
rect 27916 36540 27972 36542
rect 27804 36092 27860 36148
rect 28252 36482 28308 36484
rect 28252 36430 28254 36482
rect 28254 36430 28306 36482
rect 28306 36430 28308 36482
rect 28252 36428 28308 36430
rect 28140 35586 28196 35588
rect 28140 35534 28142 35586
rect 28142 35534 28194 35586
rect 28194 35534 28196 35586
rect 28140 35532 28196 35534
rect 28588 37266 28644 37268
rect 28588 37214 28590 37266
rect 28590 37214 28642 37266
rect 28642 37214 28644 37266
rect 28588 37212 28644 37214
rect 28028 35196 28084 35252
rect 27580 34802 27636 34804
rect 27580 34750 27582 34802
rect 27582 34750 27634 34802
rect 27634 34750 27636 34802
rect 27580 34748 27636 34750
rect 28140 34748 28196 34804
rect 28476 35026 28532 35028
rect 28476 34974 28478 35026
rect 28478 34974 28530 35026
rect 28530 34974 28532 35026
rect 28476 34972 28532 34974
rect 28588 34914 28644 34916
rect 28588 34862 28590 34914
rect 28590 34862 28642 34914
rect 28642 34862 28644 34914
rect 28588 34860 28644 34862
rect 27804 33404 27860 33460
rect 28140 34018 28196 34020
rect 28140 33966 28142 34018
rect 28142 33966 28194 34018
rect 28194 33966 28196 34018
rect 28140 33964 28196 33966
rect 28028 33906 28084 33908
rect 28028 33854 28030 33906
rect 28030 33854 28082 33906
rect 28082 33854 28084 33906
rect 28028 33852 28084 33854
rect 27916 32674 27972 32676
rect 27916 32622 27918 32674
rect 27918 32622 27970 32674
rect 27970 32622 27972 32674
rect 27916 32620 27972 32622
rect 27692 31500 27748 31556
rect 27244 31164 27300 31220
rect 27356 30994 27412 30996
rect 27356 30942 27358 30994
rect 27358 30942 27410 30994
rect 27410 30942 27412 30994
rect 27356 30940 27412 30942
rect 27692 30380 27748 30436
rect 27244 29708 27300 29764
rect 27356 29260 27412 29316
rect 26796 29148 26852 29204
rect 27580 29708 27636 29764
rect 27468 27916 27524 27972
rect 26684 27804 26740 27860
rect 25452 24892 25508 24948
rect 25116 23772 25172 23828
rect 26348 26796 26404 26852
rect 26236 26514 26292 26516
rect 26236 26462 26238 26514
rect 26238 26462 26290 26514
rect 26290 26462 26292 26514
rect 26236 26460 26292 26462
rect 25900 26012 25956 26068
rect 26124 26236 26180 26292
rect 26124 25900 26180 25956
rect 25676 24780 25732 24836
rect 25900 24892 25956 24948
rect 25676 24610 25732 24612
rect 25676 24558 25678 24610
rect 25678 24558 25730 24610
rect 25730 24558 25732 24610
rect 25676 24556 25732 24558
rect 25900 24444 25956 24500
rect 25228 23100 25284 23156
rect 26572 27132 26628 27188
rect 27580 27804 27636 27860
rect 27804 30044 27860 30100
rect 28252 33458 28308 33460
rect 28252 33406 28254 33458
rect 28254 33406 28306 33458
rect 28306 33406 28308 33458
rect 28252 33404 28308 33406
rect 28252 32786 28308 32788
rect 28252 32734 28254 32786
rect 28254 32734 28306 32786
rect 28306 32734 28308 32786
rect 28252 32732 28308 32734
rect 29372 43538 29428 43540
rect 29372 43486 29374 43538
rect 29374 43486 29426 43538
rect 29426 43486 29428 43538
rect 29372 43484 29428 43486
rect 29820 43708 29876 43764
rect 30156 44940 30212 44996
rect 30156 44044 30212 44100
rect 31276 46844 31332 46900
rect 31500 47458 31556 47460
rect 31500 47406 31502 47458
rect 31502 47406 31554 47458
rect 31554 47406 31556 47458
rect 31500 47404 31556 47406
rect 32844 53676 32900 53732
rect 32844 52556 32900 52612
rect 33964 56364 34020 56420
rect 33740 55132 33796 55188
rect 33964 55132 34020 55188
rect 33852 54402 33908 54404
rect 33852 54350 33854 54402
rect 33854 54350 33906 54402
rect 33906 54350 33908 54402
rect 33852 54348 33908 54350
rect 34748 59330 34804 59332
rect 34748 59278 34750 59330
rect 34750 59278 34802 59330
rect 34802 59278 34804 59330
rect 34748 59276 34804 59278
rect 35532 59106 35588 59108
rect 35532 59054 35534 59106
rect 35534 59054 35586 59106
rect 35586 59054 35588 59106
rect 35532 59052 35588 59054
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 34524 56588 34580 56644
rect 34076 54124 34132 54180
rect 34188 56476 34244 56532
rect 32844 52220 32900 52276
rect 43708 58380 43764 58436
rect 36092 58156 36148 58212
rect 36428 57762 36484 57764
rect 36428 57710 36430 57762
rect 36430 57710 36482 57762
rect 36482 57710 36484 57762
rect 36428 57708 36484 57710
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 34636 56364 34692 56420
rect 35420 56082 35476 56084
rect 35420 56030 35422 56082
rect 35422 56030 35474 56082
rect 35474 56030 35476 56082
rect 35420 56028 35476 56030
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35308 55522 35364 55524
rect 35308 55470 35310 55522
rect 35310 55470 35362 55522
rect 35362 55470 35364 55522
rect 35308 55468 35364 55470
rect 35644 55356 35700 55412
rect 34636 54348 34692 54404
rect 36092 56028 36148 56084
rect 35868 55074 35924 55076
rect 35868 55022 35870 55074
rect 35870 55022 35922 55074
rect 35922 55022 35924 55074
rect 35868 55020 35924 55022
rect 35868 54572 35924 54628
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35084 53788 35140 53844
rect 34300 53618 34356 53620
rect 34300 53566 34302 53618
rect 34302 53566 34354 53618
rect 34354 53566 34356 53618
rect 34300 53564 34356 53566
rect 34188 53004 34244 53060
rect 34524 53452 34580 53508
rect 33292 52780 33348 52836
rect 32396 51602 32452 51604
rect 32396 51550 32398 51602
rect 32398 51550 32450 51602
rect 32450 51550 32452 51602
rect 32396 51548 32452 51550
rect 32396 51324 32452 51380
rect 32508 50876 32564 50932
rect 32620 50540 32676 50596
rect 32732 50092 32788 50148
rect 32060 47628 32116 47684
rect 32172 48972 32228 49028
rect 31948 47180 32004 47236
rect 32284 47404 32340 47460
rect 32172 47180 32228 47236
rect 30940 45778 30996 45780
rect 30940 45726 30942 45778
rect 30942 45726 30994 45778
rect 30994 45726 30996 45778
rect 30940 45724 30996 45726
rect 31164 45890 31220 45892
rect 31164 45838 31166 45890
rect 31166 45838 31218 45890
rect 31218 45838 31220 45890
rect 31164 45836 31220 45838
rect 30380 45388 30436 45444
rect 31388 45500 31444 45556
rect 31164 44604 31220 44660
rect 30268 43820 30324 43876
rect 29596 43484 29652 43540
rect 29708 42812 29764 42868
rect 29932 43260 29988 43316
rect 30044 43484 30100 43540
rect 29708 42588 29764 42644
rect 29036 40908 29092 40964
rect 29036 40348 29092 40404
rect 29148 40012 29204 40068
rect 28924 39900 28980 39956
rect 29372 40684 29428 40740
rect 29484 40626 29540 40628
rect 29484 40574 29486 40626
rect 29486 40574 29538 40626
rect 29538 40574 29540 40626
rect 29484 40572 29540 40574
rect 29148 39452 29204 39508
rect 28924 38444 28980 38500
rect 28924 38108 28980 38164
rect 29596 39618 29652 39620
rect 29596 39566 29598 39618
rect 29598 39566 29650 39618
rect 29650 39566 29652 39618
rect 29596 39564 29652 39566
rect 29484 38892 29540 38948
rect 29148 37938 29204 37940
rect 29148 37886 29150 37938
rect 29150 37886 29202 37938
rect 29202 37886 29204 37938
rect 29148 37884 29204 37886
rect 29036 37212 29092 37268
rect 29148 37660 29204 37716
rect 29372 35532 29428 35588
rect 29372 34690 29428 34692
rect 29372 34638 29374 34690
rect 29374 34638 29426 34690
rect 29426 34638 29428 34690
rect 29372 34636 29428 34638
rect 29260 34300 29316 34356
rect 29596 34972 29652 35028
rect 29372 33404 29428 33460
rect 28812 33180 28868 33236
rect 28812 32786 28868 32788
rect 28812 32734 28814 32786
rect 28814 32734 28866 32786
rect 28866 32734 28868 32786
rect 28812 32732 28868 32734
rect 28476 32620 28532 32676
rect 28364 31890 28420 31892
rect 28364 31838 28366 31890
rect 28366 31838 28418 31890
rect 28418 31838 28420 31890
rect 28364 31836 28420 31838
rect 28924 32562 28980 32564
rect 28924 32510 28926 32562
rect 28926 32510 28978 32562
rect 28978 32510 28980 32562
rect 28924 32508 28980 32510
rect 28700 31836 28756 31892
rect 28252 31164 28308 31220
rect 26796 27020 26852 27076
rect 26908 27132 26964 27188
rect 26684 26796 26740 26852
rect 26236 25506 26292 25508
rect 26236 25454 26238 25506
rect 26238 25454 26290 25506
rect 26290 25454 26292 25506
rect 26236 25452 26292 25454
rect 25788 23772 25844 23828
rect 26684 25116 26740 25172
rect 26348 24162 26404 24164
rect 26348 24110 26350 24162
rect 26350 24110 26402 24162
rect 26402 24110 26404 24162
rect 26348 24108 26404 24110
rect 26236 23772 26292 23828
rect 26124 23548 26180 23604
rect 26460 23212 26516 23268
rect 25228 22428 25284 22484
rect 26460 22370 26516 22372
rect 26460 22318 26462 22370
rect 26462 22318 26514 22370
rect 26514 22318 26516 22370
rect 26460 22316 26516 22318
rect 25004 22092 25060 22148
rect 24668 21756 24724 21812
rect 24556 21586 24612 21588
rect 24556 21534 24558 21586
rect 24558 21534 24610 21586
rect 24610 21534 24612 21586
rect 24556 21532 24612 21534
rect 24108 21196 24164 21252
rect 25116 21644 25172 21700
rect 25004 21196 25060 21252
rect 24892 20972 24948 21028
rect 26460 21698 26516 21700
rect 26460 21646 26462 21698
rect 26462 21646 26514 21698
rect 26514 21646 26516 21698
rect 26460 21644 26516 21646
rect 25340 21586 25396 21588
rect 25340 21534 25342 21586
rect 25342 21534 25394 21586
rect 25394 21534 25396 21586
rect 25340 21532 25396 21534
rect 25228 21084 25284 21140
rect 24332 20188 24388 20244
rect 24108 20076 24164 20132
rect 24108 19852 24164 19908
rect 24220 19740 24276 19796
rect 24220 18956 24276 19012
rect 24332 19068 24388 19124
rect 23772 18284 23828 18340
rect 23884 18060 23940 18116
rect 23772 17164 23828 17220
rect 24668 20076 24724 20132
rect 25452 20018 25508 20020
rect 25452 19966 25454 20018
rect 25454 19966 25506 20018
rect 25506 19966 25508 20018
rect 25452 19964 25508 19966
rect 25228 19628 25284 19684
rect 24668 19122 24724 19124
rect 24668 19070 24670 19122
rect 24670 19070 24722 19122
rect 24722 19070 24724 19122
rect 24668 19068 24724 19070
rect 24556 18844 24612 18900
rect 24668 18620 24724 18676
rect 24668 17388 24724 17444
rect 24556 17106 24612 17108
rect 24556 17054 24558 17106
rect 24558 17054 24610 17106
rect 24610 17054 24612 17106
rect 24556 17052 24612 17054
rect 23884 16994 23940 16996
rect 23884 16942 23886 16994
rect 23886 16942 23938 16994
rect 23938 16942 23940 16994
rect 23884 16940 23940 16942
rect 23548 16882 23604 16884
rect 23548 16830 23550 16882
rect 23550 16830 23602 16882
rect 23602 16830 23604 16882
rect 23548 16828 23604 16830
rect 23996 16770 24052 16772
rect 23996 16718 23998 16770
rect 23998 16718 24050 16770
rect 24050 16718 24052 16770
rect 23996 16716 24052 16718
rect 23436 15986 23492 15988
rect 23436 15934 23438 15986
rect 23438 15934 23490 15986
rect 23490 15934 23492 15986
rect 23436 15932 23492 15934
rect 24108 15874 24164 15876
rect 24108 15822 24110 15874
rect 24110 15822 24162 15874
rect 24162 15822 24164 15874
rect 24108 15820 24164 15822
rect 23324 15596 23380 15652
rect 23212 15202 23268 15204
rect 23212 15150 23214 15202
rect 23214 15150 23266 15202
rect 23266 15150 23268 15202
rect 23212 15148 23268 15150
rect 22204 13468 22260 13524
rect 21980 13356 22036 13412
rect 22652 13244 22708 13300
rect 22092 12738 22148 12740
rect 22092 12686 22094 12738
rect 22094 12686 22146 12738
rect 22146 12686 22148 12738
rect 22092 12684 22148 12686
rect 22876 14364 22932 14420
rect 23100 13468 23156 13524
rect 23436 15314 23492 15316
rect 23436 15262 23438 15314
rect 23438 15262 23490 15314
rect 23490 15262 23492 15314
rect 23436 15260 23492 15262
rect 24108 15202 24164 15204
rect 24108 15150 24110 15202
rect 24110 15150 24162 15202
rect 24162 15150 24164 15202
rect 24108 15148 24164 15150
rect 24556 16044 24612 16100
rect 24332 15820 24388 15876
rect 24332 15314 24388 15316
rect 24332 15262 24334 15314
rect 24334 15262 24386 15314
rect 24386 15262 24388 15314
rect 24332 15260 24388 15262
rect 23772 14476 23828 14532
rect 23996 14364 24052 14420
rect 24444 14924 24500 14980
rect 23660 13634 23716 13636
rect 23660 13582 23662 13634
rect 23662 13582 23714 13634
rect 23714 13582 23716 13634
rect 23660 13580 23716 13582
rect 22876 13132 22932 13188
rect 22988 13244 23044 13300
rect 22876 12962 22932 12964
rect 22876 12910 22878 12962
rect 22878 12910 22930 12962
rect 22930 12910 22932 12962
rect 22876 12908 22932 12910
rect 21980 12236 22036 12292
rect 22092 12460 22148 12516
rect 22428 12348 22484 12404
rect 22316 12290 22372 12292
rect 22316 12238 22318 12290
rect 22318 12238 22370 12290
rect 22370 12238 22372 12290
rect 22316 12236 22372 12238
rect 22764 12348 22820 12404
rect 22316 11900 22372 11956
rect 21868 11394 21924 11396
rect 21868 11342 21870 11394
rect 21870 11342 21922 11394
rect 21922 11342 21924 11394
rect 21868 11340 21924 11342
rect 21868 10834 21924 10836
rect 21868 10782 21870 10834
rect 21870 10782 21922 10834
rect 21922 10782 21924 10834
rect 21868 10780 21924 10782
rect 22092 10834 22148 10836
rect 22092 10782 22094 10834
rect 22094 10782 22146 10834
rect 22146 10782 22148 10834
rect 22092 10780 22148 10782
rect 21420 9714 21476 9716
rect 21420 9662 21422 9714
rect 21422 9662 21474 9714
rect 21474 9662 21476 9714
rect 21420 9660 21476 9662
rect 21644 9660 21700 9716
rect 20188 8540 20244 8596
rect 20748 8876 20804 8932
rect 19068 5852 19124 5908
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20636 8428 20692 8484
rect 20412 8316 20468 8372
rect 20300 7586 20356 7588
rect 20300 7534 20302 7586
rect 20302 7534 20354 7586
rect 20354 7534 20356 7586
rect 20300 7532 20356 7534
rect 20076 6748 20132 6804
rect 20188 7084 20244 7140
rect 21084 9042 21140 9044
rect 21084 8990 21086 9042
rect 21086 8990 21138 9042
rect 21138 8990 21140 9042
rect 21084 8988 21140 8990
rect 21196 7644 21252 7700
rect 21084 7532 21140 7588
rect 21420 8540 21476 8596
rect 20860 6748 20916 6804
rect 19628 6578 19684 6580
rect 19628 6526 19630 6578
rect 19630 6526 19682 6578
rect 19682 6526 19684 6578
rect 19628 6524 19684 6526
rect 20412 6524 20468 6580
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20860 6300 20916 6356
rect 19852 5906 19908 5908
rect 19852 5854 19854 5906
rect 19854 5854 19906 5906
rect 19906 5854 19908 5906
rect 19852 5852 19908 5854
rect 21980 9714 22036 9716
rect 21980 9662 21982 9714
rect 21982 9662 22034 9714
rect 22034 9662 22036 9714
rect 21980 9660 22036 9662
rect 21756 8930 21812 8932
rect 21756 8878 21758 8930
rect 21758 8878 21810 8930
rect 21810 8878 21812 8930
rect 21756 8876 21812 8878
rect 21644 8428 21700 8484
rect 21644 6690 21700 6692
rect 21644 6638 21646 6690
rect 21646 6638 21698 6690
rect 21698 6638 21700 6690
rect 21644 6636 21700 6638
rect 21980 6578 22036 6580
rect 21980 6526 21982 6578
rect 21982 6526 22034 6578
rect 22034 6526 22036 6578
rect 21980 6524 22036 6526
rect 21084 6300 21140 6356
rect 20972 6130 21028 6132
rect 20972 6078 20974 6130
rect 20974 6078 21026 6130
rect 21026 6078 21028 6130
rect 20972 6076 21028 6078
rect 20860 5852 20916 5908
rect 20300 5292 20356 5348
rect 19964 5234 20020 5236
rect 19964 5182 19966 5234
rect 19966 5182 20018 5234
rect 20018 5182 20020 5234
rect 19964 5180 20020 5182
rect 21084 5292 21140 5348
rect 15484 5122 15540 5124
rect 15484 5070 15486 5122
rect 15486 5070 15538 5122
rect 15538 5070 15540 5122
rect 15484 5068 15540 5070
rect 16940 5122 16996 5124
rect 16940 5070 16942 5122
rect 16942 5070 16994 5122
rect 16994 5070 16996 5122
rect 16940 5068 16996 5070
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 22204 6802 22260 6804
rect 22204 6750 22206 6802
rect 22206 6750 22258 6802
rect 22258 6750 22260 6802
rect 22204 6748 22260 6750
rect 22540 10556 22596 10612
rect 22652 11676 22708 11732
rect 22652 11004 22708 11060
rect 22540 8876 22596 8932
rect 22428 8540 22484 8596
rect 22428 7474 22484 7476
rect 22428 7422 22430 7474
rect 22430 7422 22482 7474
rect 22482 7422 22484 7474
rect 22428 7420 22484 7422
rect 22316 6524 22372 6580
rect 22092 6300 22148 6356
rect 22204 6412 22260 6468
rect 21868 6188 21924 6244
rect 21420 6130 21476 6132
rect 21420 6078 21422 6130
rect 21422 6078 21474 6130
rect 21474 6078 21476 6130
rect 21420 6076 21476 6078
rect 21644 6076 21700 6132
rect 21644 5180 21700 5236
rect 21980 6130 22036 6132
rect 21980 6078 21982 6130
rect 21982 6078 22034 6130
rect 22034 6078 22036 6130
rect 21980 6076 22036 6078
rect 22204 6076 22260 6132
rect 22764 11340 22820 11396
rect 23212 12908 23268 12964
rect 23436 13132 23492 13188
rect 23436 12572 23492 12628
rect 23436 12178 23492 12180
rect 23436 12126 23438 12178
rect 23438 12126 23490 12178
rect 23490 12126 23492 12178
rect 23436 12124 23492 12126
rect 23996 13356 24052 13412
rect 24332 13132 24388 13188
rect 23100 11452 23156 11508
rect 23660 11900 23716 11956
rect 22876 10780 22932 10836
rect 22876 10050 22932 10052
rect 22876 9998 22878 10050
rect 22878 9998 22930 10050
rect 22930 9998 22932 10050
rect 22876 9996 22932 9998
rect 23548 11676 23604 11732
rect 23548 11116 23604 11172
rect 23660 11564 23716 11620
rect 22988 8316 23044 8372
rect 22876 7532 22932 7588
rect 23212 9826 23268 9828
rect 23212 9774 23214 9826
rect 23214 9774 23266 9826
rect 23266 9774 23268 9826
rect 23212 9772 23268 9774
rect 23548 10610 23604 10612
rect 23548 10558 23550 10610
rect 23550 10558 23602 10610
rect 23602 10558 23604 10610
rect 23548 10556 23604 10558
rect 23548 10220 23604 10276
rect 23436 9714 23492 9716
rect 23436 9662 23438 9714
rect 23438 9662 23490 9714
rect 23490 9662 23492 9714
rect 23436 9660 23492 9662
rect 23324 9436 23380 9492
rect 23324 8930 23380 8932
rect 23324 8878 23326 8930
rect 23326 8878 23378 8930
rect 23378 8878 23380 8930
rect 23324 8876 23380 8878
rect 23436 7532 23492 7588
rect 22988 6636 23044 6692
rect 23212 6412 23268 6468
rect 22428 5906 22484 5908
rect 22428 5854 22430 5906
rect 22430 5854 22482 5906
rect 22482 5854 22484 5906
rect 22428 5852 22484 5854
rect 24108 12348 24164 12404
rect 23660 7420 23716 7476
rect 23548 6636 23604 6692
rect 23548 6412 23604 6468
rect 23324 5682 23380 5684
rect 23324 5630 23326 5682
rect 23326 5630 23378 5682
rect 23378 5630 23380 5682
rect 23324 5628 23380 5630
rect 23436 6300 23492 6356
rect 22988 5234 23044 5236
rect 22988 5182 22990 5234
rect 22990 5182 23042 5234
rect 23042 5182 23044 5234
rect 22988 5180 23044 5182
rect 23212 4956 23268 5012
rect 21980 4844 22036 4900
rect 22764 4732 22820 4788
rect 16940 4284 16996 4340
rect 23772 6300 23828 6356
rect 23660 6076 23716 6132
rect 23660 5852 23716 5908
rect 23660 4732 23716 4788
rect 23772 5516 23828 5572
rect 23996 12012 24052 12068
rect 23996 11564 24052 11620
rect 23996 11228 24052 11284
rect 24332 12348 24388 12404
rect 24668 15820 24724 15876
rect 24892 19010 24948 19012
rect 24892 18958 24894 19010
rect 24894 18958 24946 19010
rect 24946 18958 24948 19010
rect 24892 18956 24948 18958
rect 24892 18396 24948 18452
rect 24892 17500 24948 17556
rect 25564 19516 25620 19572
rect 25564 18172 25620 18228
rect 25004 17052 25060 17108
rect 26236 19906 26292 19908
rect 26236 19854 26238 19906
rect 26238 19854 26290 19906
rect 26290 19854 26292 19906
rect 26236 19852 26292 19854
rect 26348 19740 26404 19796
rect 27580 26796 27636 26852
rect 27804 26908 27860 26964
rect 26684 20076 26740 20132
rect 26796 23996 26852 24052
rect 26684 19458 26740 19460
rect 26684 19406 26686 19458
rect 26686 19406 26738 19458
rect 26738 19406 26740 19458
rect 26684 19404 26740 19406
rect 26348 19180 26404 19236
rect 26236 19068 26292 19124
rect 26684 18844 26740 18900
rect 25900 18620 25956 18676
rect 25788 18562 25844 18564
rect 25788 18510 25790 18562
rect 25790 18510 25842 18562
rect 25842 18510 25844 18562
rect 25788 18508 25844 18510
rect 27132 24498 27188 24500
rect 27132 24446 27134 24498
rect 27134 24446 27186 24498
rect 27186 24446 27188 24498
rect 27132 24444 27188 24446
rect 27356 23772 27412 23828
rect 27916 26290 27972 26292
rect 27916 26238 27918 26290
rect 27918 26238 27970 26290
rect 27970 26238 27972 26290
rect 27916 26236 27972 26238
rect 28140 25228 28196 25284
rect 28140 25004 28196 25060
rect 29372 32562 29428 32564
rect 29372 32510 29374 32562
rect 29374 32510 29426 32562
rect 29426 32510 29428 32562
rect 29372 32508 29428 32510
rect 30380 43762 30436 43764
rect 30380 43710 30382 43762
rect 30382 43710 30434 43762
rect 30434 43710 30436 43762
rect 30380 43708 30436 43710
rect 30604 43596 30660 43652
rect 30604 43036 30660 43092
rect 30492 42924 30548 42980
rect 31052 43538 31108 43540
rect 31052 43486 31054 43538
rect 31054 43486 31106 43538
rect 31106 43486 31108 43538
rect 31052 43484 31108 43486
rect 31500 43372 31556 43428
rect 31164 43260 31220 43316
rect 30716 42476 30772 42532
rect 29820 41186 29876 41188
rect 29820 41134 29822 41186
rect 29822 41134 29874 41186
rect 29874 41134 29876 41186
rect 29820 41132 29876 41134
rect 29820 39788 29876 39844
rect 30156 41858 30212 41860
rect 30156 41806 30158 41858
rect 30158 41806 30210 41858
rect 30210 41806 30212 41858
rect 30156 41804 30212 41806
rect 30044 40796 30100 40852
rect 31164 42588 31220 42644
rect 31052 42476 31108 42532
rect 31388 42924 31444 42980
rect 31836 42812 31892 42868
rect 33180 49922 33236 49924
rect 33180 49870 33182 49922
rect 33182 49870 33234 49922
rect 33234 49870 33236 49922
rect 33180 49868 33236 49870
rect 33516 52332 33572 52388
rect 33404 51324 33460 51380
rect 33516 52108 33572 52164
rect 33628 51996 33684 52052
rect 36316 55244 36372 55300
rect 36428 54908 36484 54964
rect 37100 57932 37156 57988
rect 40012 58156 40068 58212
rect 39564 57820 39620 57876
rect 37324 57538 37380 57540
rect 37324 57486 37326 57538
rect 37326 57486 37378 57538
rect 37378 57486 37380 57538
rect 37324 57484 37380 57486
rect 37100 56754 37156 56756
rect 37100 56702 37102 56754
rect 37102 56702 37154 56754
rect 37154 56702 37156 56754
rect 37100 56700 37156 56702
rect 37100 56082 37156 56084
rect 37100 56030 37102 56082
rect 37102 56030 37154 56082
rect 37154 56030 37156 56082
rect 37100 56028 37156 56030
rect 36876 55468 36932 55524
rect 36540 54684 36596 54740
rect 36652 55244 36708 55300
rect 36764 54908 36820 54964
rect 35420 53506 35476 53508
rect 35420 53454 35422 53506
rect 35422 53454 35474 53506
rect 35474 53454 35476 53506
rect 35420 53452 35476 53454
rect 36204 53452 36260 53508
rect 35084 52946 35140 52948
rect 35084 52894 35086 52946
rect 35086 52894 35138 52946
rect 35138 52894 35140 52946
rect 35084 52892 35140 52894
rect 33964 51490 34020 51492
rect 33964 51438 33966 51490
rect 33966 51438 34018 51490
rect 34018 51438 34020 51490
rect 33964 51436 34020 51438
rect 33516 50706 33572 50708
rect 33516 50654 33518 50706
rect 33518 50654 33570 50706
rect 33570 50654 33572 50706
rect 33516 50652 33572 50654
rect 33180 48636 33236 48692
rect 33068 48300 33124 48356
rect 33068 47740 33124 47796
rect 33068 47516 33124 47572
rect 32508 46786 32564 46788
rect 32508 46734 32510 46786
rect 32510 46734 32562 46786
rect 32562 46734 32564 46786
rect 32508 46732 32564 46734
rect 32172 45724 32228 45780
rect 32060 43484 32116 43540
rect 32060 42812 32116 42868
rect 32172 42588 32228 42644
rect 31948 42476 32004 42532
rect 30044 40236 30100 40292
rect 30828 40908 30884 40964
rect 30492 40402 30548 40404
rect 30492 40350 30494 40402
rect 30494 40350 30546 40402
rect 30546 40350 30548 40402
rect 30492 40348 30548 40350
rect 29932 38332 29988 38388
rect 29932 37996 29988 38052
rect 30716 39004 30772 39060
rect 30268 37996 30324 38052
rect 30380 38946 30436 38948
rect 30380 38894 30382 38946
rect 30382 38894 30434 38946
rect 30434 38894 30436 38946
rect 30380 38892 30436 38894
rect 32396 45666 32452 45668
rect 32396 45614 32398 45666
rect 32398 45614 32450 45666
rect 32450 45614 32452 45666
rect 32396 45612 32452 45614
rect 34636 52668 34692 52724
rect 34300 52220 34356 52276
rect 33740 49420 33796 49476
rect 34188 49420 34244 49476
rect 33628 48860 33684 48916
rect 33740 48636 33796 48692
rect 33852 48130 33908 48132
rect 33852 48078 33854 48130
rect 33854 48078 33906 48130
rect 33906 48078 33908 48130
rect 33852 48076 33908 48078
rect 33292 45836 33348 45892
rect 33068 45724 33124 45780
rect 32844 45500 32900 45556
rect 32844 45052 32900 45108
rect 33068 43650 33124 43652
rect 33068 43598 33070 43650
rect 33070 43598 33122 43650
rect 33122 43598 33124 43650
rect 33068 43596 33124 43598
rect 32508 42866 32564 42868
rect 32508 42814 32510 42866
rect 32510 42814 32562 42866
rect 32562 42814 32564 42866
rect 32508 42812 32564 42814
rect 34076 46956 34132 47012
rect 33516 46060 33572 46116
rect 33404 45276 33460 45332
rect 33404 44940 33460 44996
rect 33292 44268 33348 44324
rect 33740 46060 33796 46116
rect 33964 45778 34020 45780
rect 33964 45726 33966 45778
rect 33966 45726 34018 45778
rect 34018 45726 34020 45778
rect 33964 45724 34020 45726
rect 33740 45106 33796 45108
rect 33740 45054 33742 45106
rect 33742 45054 33794 45106
rect 33794 45054 33796 45106
rect 33740 45052 33796 45054
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34860 52162 34916 52164
rect 34860 52110 34862 52162
rect 34862 52110 34914 52162
rect 34914 52110 34916 52162
rect 34860 52108 34916 52110
rect 34748 51996 34804 52052
rect 34636 51548 34692 51604
rect 34524 50988 34580 51044
rect 34412 48076 34468 48132
rect 34524 50540 34580 50596
rect 34300 47628 34356 47684
rect 34300 47458 34356 47460
rect 34300 47406 34302 47458
rect 34302 47406 34354 47458
rect 34354 47406 34356 47458
rect 34300 47404 34356 47406
rect 34300 45666 34356 45668
rect 34300 45614 34302 45666
rect 34302 45614 34354 45666
rect 34354 45614 34356 45666
rect 34300 45612 34356 45614
rect 33964 44994 34020 44996
rect 33964 44942 33966 44994
rect 33966 44942 34018 44994
rect 34018 44942 34020 44994
rect 33964 44940 34020 44942
rect 33628 44268 33684 44324
rect 34412 44434 34468 44436
rect 34412 44382 34414 44434
rect 34414 44382 34466 44434
rect 34466 44382 34468 44434
rect 34412 44380 34468 44382
rect 34300 44322 34356 44324
rect 34300 44270 34302 44322
rect 34302 44270 34354 44322
rect 34354 44270 34356 44322
rect 34300 44268 34356 44270
rect 34412 43708 34468 43764
rect 34300 43484 34356 43540
rect 34076 43036 34132 43092
rect 32620 42642 32676 42644
rect 32620 42590 32622 42642
rect 32622 42590 32674 42642
rect 32674 42590 32676 42642
rect 32620 42588 32676 42590
rect 32396 41916 32452 41972
rect 31836 41858 31892 41860
rect 31836 41806 31838 41858
rect 31838 41806 31890 41858
rect 31890 41806 31892 41858
rect 31836 41804 31892 41806
rect 31164 40796 31220 40852
rect 31500 40684 31556 40740
rect 31276 40236 31332 40292
rect 31164 40012 31220 40068
rect 31052 39900 31108 39956
rect 30604 38556 30660 38612
rect 30604 36988 30660 37044
rect 30380 36092 30436 36148
rect 29820 35196 29876 35252
rect 29932 34860 29988 34916
rect 29932 33346 29988 33348
rect 29932 33294 29934 33346
rect 29934 33294 29986 33346
rect 29986 33294 29988 33346
rect 29932 33292 29988 33294
rect 29932 32732 29988 32788
rect 29708 31836 29764 31892
rect 28700 30604 28756 30660
rect 28476 30380 28532 30436
rect 28700 29260 28756 29316
rect 28476 29148 28532 29204
rect 28364 28700 28420 28756
rect 28812 28364 28868 28420
rect 28588 27970 28644 27972
rect 28588 27918 28590 27970
rect 28590 27918 28642 27970
rect 28642 27918 28644 27970
rect 28588 27916 28644 27918
rect 28364 26348 28420 26404
rect 29596 30994 29652 30996
rect 29596 30942 29598 30994
rect 29598 30942 29650 30994
rect 29650 30942 29652 30994
rect 29596 30940 29652 30942
rect 29148 30380 29204 30436
rect 29036 29426 29092 29428
rect 29036 29374 29038 29426
rect 29038 29374 29090 29426
rect 29090 29374 29092 29426
rect 29036 29372 29092 29374
rect 30156 33292 30212 33348
rect 30492 32956 30548 33012
rect 30380 32508 30436 32564
rect 30268 31554 30324 31556
rect 30268 31502 30270 31554
rect 30270 31502 30322 31554
rect 30322 31502 30324 31554
rect 30268 31500 30324 31502
rect 30044 31164 30100 31220
rect 29708 29036 29764 29092
rect 29148 28754 29204 28756
rect 29148 28702 29150 28754
rect 29150 28702 29202 28754
rect 29202 28702 29204 28754
rect 29148 28700 29204 28702
rect 30492 30268 30548 30324
rect 30156 29314 30212 29316
rect 30156 29262 30158 29314
rect 30158 29262 30210 29314
rect 30210 29262 30212 29314
rect 30156 29260 30212 29262
rect 29932 28812 29988 28868
rect 28476 25676 28532 25732
rect 29036 26572 29092 26628
rect 29148 26460 29204 26516
rect 29148 26066 29204 26068
rect 29148 26014 29150 26066
rect 29150 26014 29202 26066
rect 29202 26014 29204 26066
rect 29148 26012 29204 26014
rect 28476 24220 28532 24276
rect 27916 23826 27972 23828
rect 27916 23774 27918 23826
rect 27918 23774 27970 23826
rect 27970 23774 27972 23826
rect 27916 23772 27972 23774
rect 27580 23212 27636 23268
rect 27356 21308 27412 21364
rect 27468 22428 27524 22484
rect 27916 23212 27972 23268
rect 27804 23154 27860 23156
rect 27804 23102 27806 23154
rect 27806 23102 27858 23154
rect 27858 23102 27860 23154
rect 27804 23100 27860 23102
rect 28028 22876 28084 22932
rect 28028 21196 28084 21252
rect 27244 20076 27300 20132
rect 27132 19964 27188 20020
rect 27020 18956 27076 19012
rect 27244 18508 27300 18564
rect 27020 18338 27076 18340
rect 27020 18286 27022 18338
rect 27022 18286 27074 18338
rect 27074 18286 27076 18338
rect 27020 18284 27076 18286
rect 26796 18060 26852 18116
rect 25676 17890 25732 17892
rect 25676 17838 25678 17890
rect 25678 17838 25730 17890
rect 25730 17838 25732 17890
rect 25676 17836 25732 17838
rect 26460 17948 26516 18004
rect 25116 17388 25172 17444
rect 25900 17724 25956 17780
rect 25788 16994 25844 16996
rect 25788 16942 25790 16994
rect 25790 16942 25842 16994
rect 25842 16942 25844 16994
rect 25788 16940 25844 16942
rect 25564 16716 25620 16772
rect 25564 16268 25620 16324
rect 25116 15596 25172 15652
rect 24892 15148 24948 15204
rect 24668 13468 24724 13524
rect 24556 12066 24612 12068
rect 24556 12014 24558 12066
rect 24558 12014 24610 12066
rect 24610 12014 24612 12066
rect 24556 12012 24612 12014
rect 24332 11452 24388 11508
rect 24108 10892 24164 10948
rect 24220 11116 24276 11172
rect 23996 10780 24052 10836
rect 24780 10668 24836 10724
rect 24220 10220 24276 10276
rect 25228 14530 25284 14532
rect 25228 14478 25230 14530
rect 25230 14478 25282 14530
rect 25282 14478 25284 14530
rect 25228 14476 25284 14478
rect 25340 14140 25396 14196
rect 25676 16044 25732 16100
rect 25452 14252 25508 14308
rect 25788 14476 25844 14532
rect 25564 13692 25620 13748
rect 25452 13468 25508 13524
rect 25004 12962 25060 12964
rect 25004 12910 25006 12962
rect 25006 12910 25058 12962
rect 25058 12910 25060 12962
rect 25004 12908 25060 12910
rect 25340 12178 25396 12180
rect 25340 12126 25342 12178
rect 25342 12126 25394 12178
rect 25394 12126 25396 12178
rect 25340 12124 25396 12126
rect 25228 11340 25284 11396
rect 24332 9436 24388 9492
rect 24108 9266 24164 9268
rect 24108 9214 24110 9266
rect 24110 9214 24162 9266
rect 24162 9214 24164 9266
rect 24108 9212 24164 9214
rect 24220 8370 24276 8372
rect 24220 8318 24222 8370
rect 24222 8318 24274 8370
rect 24274 8318 24276 8370
rect 24220 8316 24276 8318
rect 23884 5180 23940 5236
rect 24108 7532 24164 7588
rect 24444 8204 24500 8260
rect 25004 9100 25060 9156
rect 25228 10834 25284 10836
rect 25228 10782 25230 10834
rect 25230 10782 25282 10834
rect 25282 10782 25284 10834
rect 25228 10780 25284 10782
rect 24780 8258 24836 8260
rect 24780 8206 24782 8258
rect 24782 8206 24834 8258
rect 24834 8206 24836 8258
rect 24780 8204 24836 8206
rect 24668 8092 24724 8148
rect 24108 5516 24164 5572
rect 24556 7420 24612 7476
rect 24108 4956 24164 5012
rect 24332 6690 24388 6692
rect 24332 6638 24334 6690
rect 24334 6638 24386 6690
rect 24386 6638 24388 6690
rect 24332 6636 24388 6638
rect 24332 6130 24388 6132
rect 24332 6078 24334 6130
rect 24334 6078 24386 6130
rect 24386 6078 24388 6130
rect 24332 6076 24388 6078
rect 24220 4508 24276 4564
rect 24668 6972 24724 7028
rect 24668 6412 24724 6468
rect 25228 9996 25284 10052
rect 25452 11116 25508 11172
rect 25452 10332 25508 10388
rect 25788 13468 25844 13524
rect 26348 17164 26404 17220
rect 26012 17106 26068 17108
rect 26012 17054 26014 17106
rect 26014 17054 26066 17106
rect 26066 17054 26068 17106
rect 26012 17052 26068 17054
rect 26124 15820 26180 15876
rect 26012 15372 26068 15428
rect 26012 15148 26068 15204
rect 27244 17612 27300 17668
rect 27356 17388 27412 17444
rect 27244 17052 27300 17108
rect 27020 16828 27076 16884
rect 26796 16716 26852 16772
rect 27692 19906 27748 19908
rect 27692 19854 27694 19906
rect 27694 19854 27746 19906
rect 27746 19854 27748 19906
rect 27692 19852 27748 19854
rect 30380 28700 30436 28756
rect 29708 28642 29764 28644
rect 29708 28590 29710 28642
rect 29710 28590 29762 28642
rect 29762 28590 29764 28642
rect 29708 28588 29764 28590
rect 30492 28588 30548 28644
rect 29484 25340 29540 25396
rect 29372 23884 29428 23940
rect 29820 25228 29876 25284
rect 28588 23660 28644 23716
rect 28476 22316 28532 22372
rect 28252 22092 28308 22148
rect 28252 20018 28308 20020
rect 28252 19966 28254 20018
rect 28254 19966 28306 20018
rect 28306 19966 28308 20018
rect 28252 19964 28308 19966
rect 27580 16604 27636 16660
rect 26460 15148 26516 15204
rect 26012 14812 26068 14868
rect 26124 15036 26180 15092
rect 26124 14364 26180 14420
rect 26236 14924 26292 14980
rect 26796 15036 26852 15092
rect 26572 14364 26628 14420
rect 28140 16994 28196 16996
rect 28140 16942 28142 16994
rect 28142 16942 28194 16994
rect 28194 16942 28196 16994
rect 28140 16940 28196 16942
rect 28364 18172 28420 18228
rect 29372 23212 29428 23268
rect 31276 38722 31332 38724
rect 31276 38670 31278 38722
rect 31278 38670 31330 38722
rect 31330 38670 31332 38722
rect 31276 38668 31332 38670
rect 31724 40236 31780 40292
rect 31612 39340 31668 39396
rect 32172 41468 32228 41524
rect 32732 41580 32788 41636
rect 33740 41692 33796 41748
rect 33516 41356 33572 41412
rect 31948 38892 32004 38948
rect 32060 38668 32116 38724
rect 32172 38556 32228 38612
rect 31500 38220 31556 38276
rect 31164 38108 31220 38164
rect 32060 38162 32116 38164
rect 32060 38110 32062 38162
rect 32062 38110 32114 38162
rect 32114 38110 32116 38162
rect 32060 38108 32116 38110
rect 31948 38050 32004 38052
rect 31948 37998 31950 38050
rect 31950 37998 32002 38050
rect 32002 37998 32004 38050
rect 31948 37996 32004 37998
rect 31164 37884 31220 37940
rect 31500 37266 31556 37268
rect 31500 37214 31502 37266
rect 31502 37214 31554 37266
rect 31554 37214 31556 37266
rect 31500 37212 31556 37214
rect 32172 37100 32228 37156
rect 31612 36482 31668 36484
rect 31612 36430 31614 36482
rect 31614 36430 31666 36482
rect 31666 36430 31668 36482
rect 31612 36428 31668 36430
rect 31052 36204 31108 36260
rect 31948 36092 32004 36148
rect 33404 41074 33460 41076
rect 33404 41022 33406 41074
rect 33406 41022 33458 41074
rect 33458 41022 33460 41074
rect 33404 41020 33460 41022
rect 32732 40796 32788 40852
rect 32620 39788 32676 39844
rect 33516 40236 33572 40292
rect 34300 41186 34356 41188
rect 34300 41134 34302 41186
rect 34302 41134 34354 41186
rect 34354 41134 34356 41186
rect 34300 41132 34356 41134
rect 34972 51884 35028 51940
rect 34860 51772 34916 51828
rect 34972 51378 35028 51380
rect 34972 51326 34974 51378
rect 34974 51326 35026 51378
rect 35026 51326 35028 51378
rect 34972 51324 35028 51326
rect 35420 52220 35476 52276
rect 35532 52108 35588 52164
rect 36428 52444 36484 52500
rect 35868 52108 35924 52164
rect 36204 52162 36260 52164
rect 36204 52110 36206 52162
rect 36206 52110 36258 52162
rect 36258 52110 36260 52162
rect 36204 52108 36260 52110
rect 35420 51938 35476 51940
rect 35420 51886 35422 51938
rect 35422 51886 35474 51938
rect 35474 51886 35476 51938
rect 35420 51884 35476 51886
rect 35756 51436 35812 51492
rect 35420 51324 35476 51380
rect 35308 51212 35364 51268
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35084 50594 35140 50596
rect 35084 50542 35086 50594
rect 35086 50542 35138 50594
rect 35138 50542 35140 50594
rect 35084 50540 35140 50542
rect 34972 49250 35028 49252
rect 34972 49198 34974 49250
rect 34974 49198 35026 49250
rect 35026 49198 35028 49250
rect 34972 49196 35028 49198
rect 36316 52220 36372 52276
rect 36540 51884 36596 51940
rect 36428 51772 36484 51828
rect 35868 50540 35924 50596
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35308 48802 35364 48804
rect 35308 48750 35310 48802
rect 35310 48750 35362 48802
rect 35362 48750 35364 48802
rect 35308 48748 35364 48750
rect 35084 48636 35140 48692
rect 35308 48412 35364 48468
rect 34860 48242 34916 48244
rect 34860 48190 34862 48242
rect 34862 48190 34914 48242
rect 34914 48190 34916 48242
rect 34860 48188 34916 48190
rect 35084 48076 35140 48132
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35756 49532 35812 49588
rect 35644 48860 35700 48916
rect 35308 47628 35364 47684
rect 35644 48636 35700 48692
rect 35980 49308 36036 49364
rect 36988 55298 37044 55300
rect 36988 55246 36990 55298
rect 36990 55246 37042 55298
rect 37042 55246 37044 55298
rect 36988 55244 37044 55246
rect 36876 54572 36932 54628
rect 37212 55356 37268 55412
rect 37324 55186 37380 55188
rect 37324 55134 37326 55186
rect 37326 55134 37378 55186
rect 37378 55134 37380 55186
rect 37324 55132 37380 55134
rect 37212 54626 37268 54628
rect 37212 54574 37214 54626
rect 37214 54574 37266 54626
rect 37266 54574 37268 54626
rect 37212 54572 37268 54574
rect 36988 53676 37044 53732
rect 37212 53452 37268 53508
rect 37100 52386 37156 52388
rect 37100 52334 37102 52386
rect 37102 52334 37154 52386
rect 37154 52334 37156 52386
rect 37100 52332 37156 52334
rect 36988 52162 37044 52164
rect 36988 52110 36990 52162
rect 36990 52110 37042 52162
rect 37042 52110 37044 52162
rect 36988 52108 37044 52110
rect 36316 51212 36372 51268
rect 36316 50764 36372 50820
rect 36316 50428 36372 50484
rect 37212 51548 37268 51604
rect 37436 52780 37492 52836
rect 36092 48914 36148 48916
rect 36092 48862 36094 48914
rect 36094 48862 36146 48914
rect 36146 48862 36148 48914
rect 36092 48860 36148 48862
rect 37436 50652 37492 50708
rect 36652 50092 36708 50148
rect 37772 56476 37828 56532
rect 37996 57484 38052 57540
rect 37660 55970 37716 55972
rect 37660 55918 37662 55970
rect 37662 55918 37714 55970
rect 37714 55918 37716 55970
rect 37660 55916 37716 55918
rect 37772 55244 37828 55300
rect 38444 57148 38500 57204
rect 40684 58156 40740 58212
rect 40236 58044 40292 58100
rect 39564 56978 39620 56980
rect 39564 56926 39566 56978
rect 39566 56926 39618 56978
rect 39618 56926 39620 56978
rect 39564 56924 39620 56926
rect 39340 56700 39396 56756
rect 38556 56364 38612 56420
rect 38332 55916 38388 55972
rect 39004 56588 39060 56644
rect 39004 55970 39060 55972
rect 39004 55918 39006 55970
rect 39006 55918 39058 55970
rect 39058 55918 39060 55970
rect 39004 55916 39060 55918
rect 38892 55580 38948 55636
rect 39004 55692 39060 55748
rect 37996 55020 38052 55076
rect 38892 54908 38948 54964
rect 38444 54626 38500 54628
rect 38444 54574 38446 54626
rect 38446 54574 38498 54626
rect 38498 54574 38500 54626
rect 38444 54572 38500 54574
rect 37660 53618 37716 53620
rect 37660 53566 37662 53618
rect 37662 53566 37714 53618
rect 37714 53566 37716 53618
rect 37660 53564 37716 53566
rect 40572 57820 40628 57876
rect 40236 56700 40292 56756
rect 40460 56754 40516 56756
rect 40460 56702 40462 56754
rect 40462 56702 40514 56754
rect 40514 56702 40516 56754
rect 40460 56700 40516 56702
rect 39452 55970 39508 55972
rect 39452 55918 39454 55970
rect 39454 55918 39506 55970
rect 39506 55918 39508 55970
rect 39452 55916 39508 55918
rect 40460 56140 40516 56196
rect 39676 55298 39732 55300
rect 39676 55246 39678 55298
rect 39678 55246 39730 55298
rect 39730 55246 39732 55298
rect 39676 55244 39732 55246
rect 40124 54572 40180 54628
rect 40460 55916 40516 55972
rect 38892 54124 38948 54180
rect 38444 53340 38500 53396
rect 38108 52668 38164 52724
rect 38556 52780 38612 52836
rect 38668 53676 38724 53732
rect 38668 53004 38724 53060
rect 38444 52444 38500 52500
rect 38556 52556 38612 52612
rect 38332 51996 38388 52052
rect 37548 49868 37604 49924
rect 37436 49308 37492 49364
rect 36876 49026 36932 49028
rect 36876 48974 36878 49026
rect 36878 48974 36930 49026
rect 36930 48974 36932 49026
rect 36876 48972 36932 48974
rect 37212 48972 37268 49028
rect 36652 48748 36708 48804
rect 36316 46956 36372 47012
rect 34972 46562 35028 46564
rect 34972 46510 34974 46562
rect 34974 46510 35026 46562
rect 35026 46510 35028 46562
rect 34972 46508 35028 46510
rect 35756 46396 35812 46452
rect 34636 46172 34692 46228
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 45836 35252 45892
rect 34860 45612 34916 45668
rect 34636 45500 34692 45556
rect 35532 45388 35588 45444
rect 35196 45330 35252 45332
rect 35196 45278 35198 45330
rect 35198 45278 35250 45330
rect 35250 45278 35252 45330
rect 35196 45276 35252 45278
rect 34636 45052 34692 45108
rect 34860 44994 34916 44996
rect 34860 44942 34862 44994
rect 34862 44942 34914 44994
rect 34914 44942 34916 44994
rect 34860 44940 34916 44942
rect 34860 44380 34916 44436
rect 35420 45276 35476 45332
rect 35644 45218 35700 45220
rect 35644 45166 35646 45218
rect 35646 45166 35698 45218
rect 35698 45166 35700 45218
rect 35644 45164 35700 45166
rect 35420 45052 35476 45108
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35308 43708 35364 43764
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34748 41804 34804 41860
rect 35308 42642 35364 42644
rect 35308 42590 35310 42642
rect 35310 42590 35362 42642
rect 35362 42590 35364 42642
rect 35308 42588 35364 42590
rect 34860 41132 34916 41188
rect 35532 41916 35588 41972
rect 35084 41692 35140 41748
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35644 41858 35700 41860
rect 35644 41806 35646 41858
rect 35646 41806 35698 41858
rect 35698 41806 35700 41858
rect 35644 41804 35700 41806
rect 35532 41410 35588 41412
rect 35532 41358 35534 41410
rect 35534 41358 35586 41410
rect 35586 41358 35588 41410
rect 35532 41356 35588 41358
rect 35084 41020 35140 41076
rect 34524 40908 34580 40964
rect 34972 40796 35028 40852
rect 34188 40348 34244 40404
rect 34860 40402 34916 40404
rect 34860 40350 34862 40402
rect 34862 40350 34914 40402
rect 34914 40350 34916 40402
rect 34860 40348 34916 40350
rect 34636 40236 34692 40292
rect 34524 39788 34580 39844
rect 33964 39506 34020 39508
rect 33964 39454 33966 39506
rect 33966 39454 34018 39506
rect 34018 39454 34020 39506
rect 33964 39452 34020 39454
rect 32508 38834 32564 38836
rect 32508 38782 32510 38834
rect 32510 38782 32562 38834
rect 32562 38782 32564 38834
rect 32508 38780 32564 38782
rect 32956 38444 33012 38500
rect 32956 38220 33012 38276
rect 32508 37490 32564 37492
rect 32508 37438 32510 37490
rect 32510 37438 32562 37490
rect 32562 37438 32564 37490
rect 32508 37436 32564 37438
rect 31836 34748 31892 34804
rect 30828 33292 30884 33348
rect 31164 32956 31220 33012
rect 30716 31612 30772 31668
rect 30492 26796 30548 26852
rect 30492 26012 30548 26068
rect 30044 25282 30100 25284
rect 30044 25230 30046 25282
rect 30046 25230 30098 25282
rect 30098 25230 30100 25282
rect 30044 25228 30100 25230
rect 30492 25676 30548 25732
rect 30604 24946 30660 24948
rect 30604 24894 30606 24946
rect 30606 24894 30658 24946
rect 30658 24894 30660 24946
rect 30604 24892 30660 24894
rect 30380 24220 30436 24276
rect 30940 31836 30996 31892
rect 31724 33404 31780 33460
rect 31836 33292 31892 33348
rect 31836 32562 31892 32564
rect 31836 32510 31838 32562
rect 31838 32510 31890 32562
rect 31890 32510 31892 32562
rect 31836 32508 31892 32510
rect 32396 34354 32452 34356
rect 32396 34302 32398 34354
rect 32398 34302 32450 34354
rect 32450 34302 32452 34354
rect 32396 34300 32452 34302
rect 32060 33180 32116 33236
rect 32172 33068 32228 33124
rect 32508 33628 32564 33684
rect 32732 33458 32788 33460
rect 32732 33406 32734 33458
rect 32734 33406 32786 33458
rect 32786 33406 32788 33458
rect 32732 33404 32788 33406
rect 32172 32844 32228 32900
rect 31948 31948 32004 32004
rect 31164 31218 31220 31220
rect 31164 31166 31166 31218
rect 31166 31166 31218 31218
rect 31218 31166 31220 31218
rect 31164 31164 31220 31166
rect 31948 31388 32004 31444
rect 30940 30322 30996 30324
rect 30940 30270 30942 30322
rect 30942 30270 30994 30322
rect 30994 30270 30996 30322
rect 30940 30268 30996 30270
rect 31836 30268 31892 30324
rect 32396 31612 32452 31668
rect 32508 32450 32564 32452
rect 32508 32398 32510 32450
rect 32510 32398 32562 32450
rect 32562 32398 32564 32450
rect 32508 32396 32564 32398
rect 32732 31500 32788 31556
rect 34188 38892 34244 38948
rect 33404 38834 33460 38836
rect 33404 38782 33406 38834
rect 33406 38782 33458 38834
rect 33458 38782 33460 38834
rect 33404 38780 33460 38782
rect 33292 37996 33348 38052
rect 33404 38108 33460 38164
rect 33068 36204 33124 36260
rect 34300 38444 34356 38500
rect 36652 48188 36708 48244
rect 36652 47404 36708 47460
rect 36428 46844 36484 46900
rect 36988 47292 37044 47348
rect 36316 45836 36372 45892
rect 35868 45164 35924 45220
rect 36316 45052 36372 45108
rect 36540 44492 36596 44548
rect 36876 45052 36932 45108
rect 36204 44322 36260 44324
rect 36204 44270 36206 44322
rect 36206 44270 36258 44322
rect 36258 44270 36260 44322
rect 36204 44268 36260 44270
rect 37324 48748 37380 48804
rect 38780 52722 38836 52724
rect 38780 52670 38782 52722
rect 38782 52670 38834 52722
rect 38834 52670 38836 52722
rect 38780 52668 38836 52670
rect 38892 52108 38948 52164
rect 39340 53058 39396 53060
rect 39340 53006 39342 53058
rect 39342 53006 39394 53058
rect 39394 53006 39396 53058
rect 39340 53004 39396 53006
rect 39228 52108 39284 52164
rect 40012 53730 40068 53732
rect 40012 53678 40014 53730
rect 40014 53678 40066 53730
rect 40066 53678 40068 53730
rect 40012 53676 40068 53678
rect 39004 50540 39060 50596
rect 39116 50764 39172 50820
rect 39228 50652 39284 50708
rect 37884 49756 37940 49812
rect 37436 48412 37492 48468
rect 37660 49196 37716 49252
rect 37884 49196 37940 49252
rect 38108 49026 38164 49028
rect 38108 48974 38110 49026
rect 38110 48974 38162 49026
rect 38162 48974 38164 49026
rect 38108 48972 38164 48974
rect 37212 48242 37268 48244
rect 37212 48190 37214 48242
rect 37214 48190 37266 48242
rect 37266 48190 37268 48242
rect 37212 48188 37268 48190
rect 37772 48524 37828 48580
rect 38108 48524 38164 48580
rect 38108 47964 38164 48020
rect 37884 47852 37940 47908
rect 37212 47628 37268 47684
rect 37212 47346 37268 47348
rect 37212 47294 37214 47346
rect 37214 47294 37266 47346
rect 37266 47294 37268 47346
rect 37212 47292 37268 47294
rect 37548 45500 37604 45556
rect 37212 45106 37268 45108
rect 37212 45054 37214 45106
rect 37214 45054 37266 45106
rect 37266 45054 37268 45106
rect 37212 45052 37268 45054
rect 37100 44940 37156 44996
rect 36988 44156 37044 44212
rect 36876 43596 36932 43652
rect 36652 43538 36708 43540
rect 36652 43486 36654 43538
rect 36654 43486 36706 43538
rect 36706 43486 36708 43538
rect 36652 43484 36708 43486
rect 35756 40684 35812 40740
rect 35868 40962 35924 40964
rect 35868 40910 35870 40962
rect 35870 40910 35922 40962
rect 35922 40910 35924 40962
rect 35868 40908 35924 40910
rect 35420 40290 35476 40292
rect 35420 40238 35422 40290
rect 35422 40238 35474 40290
rect 35474 40238 35476 40290
rect 35420 40236 35476 40238
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34076 38050 34132 38052
rect 34076 37998 34078 38050
rect 34078 37998 34130 38050
rect 34130 37998 34132 38050
rect 34076 37996 34132 37998
rect 34076 37660 34132 37716
rect 33852 37154 33908 37156
rect 33852 37102 33854 37154
rect 33854 37102 33906 37154
rect 33906 37102 33908 37154
rect 33852 37100 33908 37102
rect 33628 36988 33684 37044
rect 32956 35196 33012 35252
rect 33180 34300 33236 34356
rect 33068 33346 33124 33348
rect 33068 33294 33070 33346
rect 33070 33294 33122 33346
rect 33122 33294 33124 33346
rect 33068 33292 33124 33294
rect 33292 33234 33348 33236
rect 33292 33182 33294 33234
rect 33294 33182 33346 33234
rect 33346 33182 33348 33234
rect 33292 33180 33348 33182
rect 33516 32786 33572 32788
rect 33516 32734 33518 32786
rect 33518 32734 33570 32786
rect 33570 32734 33572 32786
rect 33516 32732 33572 32734
rect 33068 32396 33124 32452
rect 34188 37212 34244 37268
rect 36092 40514 36148 40516
rect 36092 40462 36094 40514
rect 36094 40462 36146 40514
rect 36146 40462 36148 40514
rect 36092 40460 36148 40462
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34636 37884 34692 37940
rect 34412 36988 34468 37044
rect 34524 37436 34580 37492
rect 34076 35084 34132 35140
rect 33740 33292 33796 33348
rect 32956 31666 33012 31668
rect 32956 31614 32958 31666
rect 32958 31614 33010 31666
rect 33010 31614 33012 31666
rect 32956 31612 33012 31614
rect 33852 32562 33908 32564
rect 33852 32510 33854 32562
rect 33854 32510 33906 32562
rect 33906 32510 33908 32562
rect 33852 32508 33908 32510
rect 34412 35698 34468 35700
rect 34412 35646 34414 35698
rect 34414 35646 34466 35698
rect 34466 35646 34468 35698
rect 34412 35644 34468 35646
rect 34412 33346 34468 33348
rect 34412 33294 34414 33346
rect 34414 33294 34466 33346
rect 34466 33294 34468 33346
rect 34412 33292 34468 33294
rect 34524 33180 34580 33236
rect 34412 32956 34468 33012
rect 34188 32002 34244 32004
rect 34188 31950 34190 32002
rect 34190 31950 34242 32002
rect 34242 31950 34244 32002
rect 34188 31948 34244 31950
rect 34300 32396 34356 32452
rect 33740 31724 33796 31780
rect 32844 31388 32900 31444
rect 34524 32396 34580 32452
rect 34524 31666 34580 31668
rect 34524 31614 34526 31666
rect 34526 31614 34578 31666
rect 34578 31614 34580 31666
rect 34524 31612 34580 31614
rect 33852 31500 33908 31556
rect 35084 37772 35140 37828
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 34972 36428 35028 36484
rect 34860 36370 34916 36372
rect 34860 36318 34862 36370
rect 34862 36318 34914 36370
rect 34914 36318 34916 36370
rect 34860 36316 34916 36318
rect 35084 36092 35140 36148
rect 35420 36258 35476 36260
rect 35420 36206 35422 36258
rect 35422 36206 35474 36258
rect 35474 36206 35476 36258
rect 35420 36204 35476 36206
rect 35420 35922 35476 35924
rect 35420 35870 35422 35922
rect 35422 35870 35474 35922
rect 35474 35870 35476 35922
rect 35420 35868 35476 35870
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 36764 41916 36820 41972
rect 37436 44492 37492 44548
rect 37324 44268 37380 44324
rect 38780 49586 38836 49588
rect 38780 49534 38782 49586
rect 38782 49534 38834 49586
rect 38834 49534 38836 49586
rect 38780 49532 38836 49534
rect 38556 49026 38612 49028
rect 38556 48974 38558 49026
rect 38558 48974 38610 49026
rect 38610 48974 38612 49026
rect 38556 48972 38612 48974
rect 38444 47852 38500 47908
rect 38220 45778 38276 45780
rect 38220 45726 38222 45778
rect 38222 45726 38274 45778
rect 38274 45726 38276 45778
rect 38220 45724 38276 45726
rect 39564 50428 39620 50484
rect 39452 48914 39508 48916
rect 39452 48862 39454 48914
rect 39454 48862 39506 48914
rect 39506 48862 39508 48914
rect 39452 48860 39508 48862
rect 39228 48412 39284 48468
rect 39900 51548 39956 51604
rect 41132 58210 41188 58212
rect 41132 58158 41134 58210
rect 41134 58158 41186 58210
rect 41186 58158 41188 58210
rect 41132 58156 41188 58158
rect 41244 57538 41300 57540
rect 41244 57486 41246 57538
rect 41246 57486 41298 57538
rect 41298 57486 41300 57538
rect 41244 57484 41300 57486
rect 40908 56924 40964 56980
rect 41356 56978 41412 56980
rect 41356 56926 41358 56978
rect 41358 56926 41410 56978
rect 41410 56926 41412 56978
rect 41356 56924 41412 56926
rect 42252 57874 42308 57876
rect 42252 57822 42254 57874
rect 42254 57822 42306 57874
rect 42306 57822 42308 57874
rect 42252 57820 42308 57822
rect 47516 58268 47572 58324
rect 44492 58156 44548 58212
rect 41468 55970 41524 55972
rect 41468 55918 41470 55970
rect 41470 55918 41522 55970
rect 41522 55918 41524 55970
rect 41468 55916 41524 55918
rect 41020 55692 41076 55748
rect 41020 55522 41076 55524
rect 41020 55470 41022 55522
rect 41022 55470 41074 55522
rect 41074 55470 41076 55522
rect 41020 55468 41076 55470
rect 40796 55244 40852 55300
rect 40460 53900 40516 53956
rect 39788 50764 39844 50820
rect 40124 50764 40180 50820
rect 39676 48636 39732 48692
rect 40348 50316 40404 50372
rect 40348 49922 40404 49924
rect 40348 49870 40350 49922
rect 40350 49870 40402 49922
rect 40402 49870 40404 49922
rect 40348 49868 40404 49870
rect 40236 48524 40292 48580
rect 40124 48466 40180 48468
rect 40124 48414 40126 48466
rect 40126 48414 40178 48466
rect 40178 48414 40180 48466
rect 40124 48412 40180 48414
rect 40012 48354 40068 48356
rect 40012 48302 40014 48354
rect 40014 48302 40066 48354
rect 40066 48302 40068 48354
rect 40012 48300 40068 48302
rect 39564 48242 39620 48244
rect 39564 48190 39566 48242
rect 39566 48190 39618 48242
rect 39618 48190 39620 48242
rect 39564 48188 39620 48190
rect 40348 48242 40404 48244
rect 40348 48190 40350 48242
rect 40350 48190 40402 48242
rect 40402 48190 40404 48242
rect 40348 48188 40404 48190
rect 40012 48130 40068 48132
rect 40012 48078 40014 48130
rect 40014 48078 40066 48130
rect 40066 48078 40068 48130
rect 40012 48076 40068 48078
rect 39228 47516 39284 47572
rect 40236 47852 40292 47908
rect 40012 47404 40068 47460
rect 39116 47346 39172 47348
rect 39116 47294 39118 47346
rect 39118 47294 39170 47346
rect 39170 47294 39172 47346
rect 39116 47292 39172 47294
rect 38780 46732 38836 46788
rect 37996 44828 38052 44884
rect 37884 44492 37940 44548
rect 37548 44044 37604 44100
rect 37884 44156 37940 44212
rect 37660 43484 37716 43540
rect 37772 43650 37828 43652
rect 37772 43598 37774 43650
rect 37774 43598 37826 43650
rect 37826 43598 37828 43650
rect 37772 43596 37828 43598
rect 38108 44716 38164 44772
rect 38108 44268 38164 44324
rect 38108 43148 38164 43204
rect 37884 42700 37940 42756
rect 36988 41356 37044 41412
rect 37772 41970 37828 41972
rect 37772 41918 37774 41970
rect 37774 41918 37826 41970
rect 37826 41918 37828 41970
rect 37772 41916 37828 41918
rect 38108 41410 38164 41412
rect 38108 41358 38110 41410
rect 38110 41358 38162 41410
rect 38162 41358 38164 41410
rect 38108 41356 38164 41358
rect 37772 41244 37828 41300
rect 37884 41186 37940 41188
rect 37884 41134 37886 41186
rect 37886 41134 37938 41186
rect 37938 41134 37940 41186
rect 37884 41132 37940 41134
rect 36428 39788 36484 39844
rect 36092 38050 36148 38052
rect 36092 37998 36094 38050
rect 36094 37998 36146 38050
rect 36146 37998 36148 38050
rect 36092 37996 36148 37998
rect 35308 34972 35364 35028
rect 35644 36428 35700 36484
rect 35532 34188 35588 34244
rect 36540 37324 36596 37380
rect 37212 41074 37268 41076
rect 37212 41022 37214 41074
rect 37214 41022 37266 41074
rect 37266 41022 37268 41074
rect 37212 41020 37268 41022
rect 36988 40962 37044 40964
rect 36988 40910 36990 40962
rect 36990 40910 37042 40962
rect 37042 40910 37044 40962
rect 36988 40908 37044 40910
rect 36876 40796 36932 40852
rect 36652 39340 36708 39396
rect 36316 37212 36372 37268
rect 35756 36316 35812 36372
rect 36204 36876 36260 36932
rect 36204 36092 36260 36148
rect 36428 36370 36484 36372
rect 36428 36318 36430 36370
rect 36430 36318 36482 36370
rect 36482 36318 36484 36370
rect 36428 36316 36484 36318
rect 36540 36988 36596 37044
rect 36876 40348 36932 40404
rect 37436 40962 37492 40964
rect 37436 40910 37438 40962
rect 37438 40910 37490 40962
rect 37490 40910 37492 40962
rect 37436 40908 37492 40910
rect 37212 40514 37268 40516
rect 37212 40462 37214 40514
rect 37214 40462 37266 40514
rect 37266 40462 37268 40514
rect 37212 40460 37268 40462
rect 37436 40348 37492 40404
rect 37324 38556 37380 38612
rect 37100 37826 37156 37828
rect 37100 37774 37102 37826
rect 37102 37774 37154 37826
rect 37154 37774 37156 37826
rect 37100 37772 37156 37774
rect 36988 37436 37044 37492
rect 36876 37212 36932 37268
rect 36652 36876 36708 36932
rect 36876 36988 36932 37044
rect 36652 36204 36708 36260
rect 36204 35084 36260 35140
rect 36092 34636 36148 34692
rect 35868 34188 35924 34244
rect 36092 34242 36148 34244
rect 36092 34190 36094 34242
rect 36094 34190 36146 34242
rect 36146 34190 36148 34242
rect 36092 34188 36148 34190
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35084 32844 35140 32900
rect 35420 33346 35476 33348
rect 35420 33294 35422 33346
rect 35422 33294 35474 33346
rect 35474 33294 35476 33346
rect 35420 33292 35476 33294
rect 36316 34130 36372 34132
rect 36316 34078 36318 34130
rect 36318 34078 36370 34130
rect 36370 34078 36372 34130
rect 36316 34076 36372 34078
rect 36540 34412 36596 34468
rect 35532 32844 35588 32900
rect 34972 31890 35028 31892
rect 34972 31838 34974 31890
rect 34974 31838 35026 31890
rect 35026 31838 35028 31890
rect 34972 31836 35028 31838
rect 34748 31500 34804 31556
rect 33516 30156 33572 30212
rect 32060 30044 32116 30100
rect 33852 30044 33908 30100
rect 31948 29932 32004 29988
rect 32396 29650 32452 29652
rect 32396 29598 32398 29650
rect 32398 29598 32450 29650
rect 32450 29598 32452 29650
rect 32396 29596 32452 29598
rect 33180 29596 33236 29652
rect 31276 29538 31332 29540
rect 31276 29486 31278 29538
rect 31278 29486 31330 29538
rect 31330 29486 31332 29538
rect 31276 29484 31332 29486
rect 33068 29484 33124 29540
rect 31052 28866 31108 28868
rect 31052 28814 31054 28866
rect 31054 28814 31106 28866
rect 31106 28814 31108 28866
rect 31052 28812 31108 28814
rect 33180 29148 33236 29204
rect 32508 28700 32564 28756
rect 32620 28812 32676 28868
rect 31164 28642 31220 28644
rect 31164 28590 31166 28642
rect 31166 28590 31218 28642
rect 31218 28590 31220 28642
rect 31164 28588 31220 28590
rect 31388 28588 31444 28644
rect 31164 28364 31220 28420
rect 31276 27746 31332 27748
rect 31276 27694 31278 27746
rect 31278 27694 31330 27746
rect 31330 27694 31332 27746
rect 31276 27692 31332 27694
rect 30828 26796 30884 26852
rect 30828 25340 30884 25396
rect 30828 25116 30884 25172
rect 31500 28252 31556 28308
rect 31500 27580 31556 27636
rect 31612 27356 31668 27412
rect 32396 28364 32452 28420
rect 31724 27804 31780 27860
rect 31164 26290 31220 26292
rect 31164 26238 31166 26290
rect 31166 26238 31218 26290
rect 31218 26238 31220 26290
rect 31164 26236 31220 26238
rect 30044 23660 30100 23716
rect 29596 22988 29652 23044
rect 29708 23100 29764 23156
rect 29260 22930 29316 22932
rect 29260 22878 29262 22930
rect 29262 22878 29314 22930
rect 29314 22878 29316 22930
rect 29260 22876 29316 22878
rect 29148 22428 29204 22484
rect 29372 22316 29428 22372
rect 29932 23378 29988 23380
rect 29932 23326 29934 23378
rect 29934 23326 29986 23378
rect 29986 23326 29988 23378
rect 29932 23324 29988 23326
rect 29932 22540 29988 22596
rect 29260 21474 29316 21476
rect 29260 21422 29262 21474
rect 29262 21422 29314 21474
rect 29314 21422 29316 21474
rect 29260 21420 29316 21422
rect 30044 21474 30100 21476
rect 30044 21422 30046 21474
rect 30046 21422 30098 21474
rect 30098 21422 30100 21474
rect 30044 21420 30100 21422
rect 29932 21308 29988 21364
rect 30268 23324 30324 23380
rect 30604 23714 30660 23716
rect 30604 23662 30606 23714
rect 30606 23662 30658 23714
rect 30658 23662 30660 23714
rect 30604 23660 30660 23662
rect 30380 23100 30436 23156
rect 30492 23548 30548 23604
rect 30492 22988 30548 23044
rect 30828 23714 30884 23716
rect 30828 23662 30830 23714
rect 30830 23662 30882 23714
rect 30882 23662 30884 23714
rect 30828 23660 30884 23662
rect 30716 22092 30772 22148
rect 31388 26178 31444 26180
rect 31388 26126 31390 26178
rect 31390 26126 31442 26178
rect 31442 26126 31444 26178
rect 31388 26124 31444 26126
rect 31276 25116 31332 25172
rect 31164 25004 31220 25060
rect 31948 28252 32004 28308
rect 32956 28252 33012 28308
rect 31948 27132 32004 27188
rect 31052 23324 31108 23380
rect 31836 24780 31892 24836
rect 31388 24722 31444 24724
rect 31388 24670 31390 24722
rect 31390 24670 31442 24722
rect 31442 24670 31444 24722
rect 31388 24668 31444 24670
rect 31388 23548 31444 23604
rect 31052 22764 31108 22820
rect 30268 21698 30324 21700
rect 30268 21646 30270 21698
rect 30270 21646 30322 21698
rect 30322 21646 30324 21698
rect 30268 21644 30324 21646
rect 29372 19852 29428 19908
rect 29820 20188 29876 20244
rect 29036 18956 29092 19012
rect 29820 20018 29876 20020
rect 29820 19966 29822 20018
rect 29822 19966 29874 20018
rect 29874 19966 29876 20018
rect 29820 19964 29876 19966
rect 29708 18732 29764 18788
rect 29820 19404 29876 19460
rect 28476 17666 28532 17668
rect 28476 17614 28478 17666
rect 28478 17614 28530 17666
rect 28530 17614 28532 17666
rect 28476 17612 28532 17614
rect 28252 16658 28308 16660
rect 28252 16606 28254 16658
rect 28254 16606 28306 16658
rect 28306 16606 28308 16658
rect 28252 16604 28308 16606
rect 28924 17052 28980 17108
rect 28924 16828 28980 16884
rect 28028 16380 28084 16436
rect 28028 15820 28084 15876
rect 27356 14700 27412 14756
rect 27356 14364 27412 14420
rect 27244 13916 27300 13972
rect 27916 15260 27972 15316
rect 27692 15036 27748 15092
rect 27804 14588 27860 14644
rect 25900 13244 25956 13300
rect 25676 12908 25732 12964
rect 25676 12178 25732 12180
rect 25676 12126 25678 12178
rect 25678 12126 25730 12178
rect 25730 12126 25732 12178
rect 25676 12124 25732 12126
rect 25900 12348 25956 12404
rect 25788 11788 25844 11844
rect 25676 11394 25732 11396
rect 25676 11342 25678 11394
rect 25678 11342 25730 11394
rect 25730 11342 25732 11394
rect 25676 11340 25732 11342
rect 25676 10444 25732 10500
rect 25116 8204 25172 8260
rect 25900 10780 25956 10836
rect 26124 12348 26180 12404
rect 26236 11900 26292 11956
rect 26908 12684 26964 12740
rect 26348 11170 26404 11172
rect 26348 11118 26350 11170
rect 26350 11118 26402 11170
rect 26402 11118 26404 11170
rect 26348 11116 26404 11118
rect 26460 12572 26516 12628
rect 27356 12572 27412 12628
rect 26796 11900 26852 11956
rect 26572 11394 26628 11396
rect 26572 11342 26574 11394
rect 26574 11342 26626 11394
rect 26626 11342 26628 11394
rect 26572 11340 26628 11342
rect 27020 11788 27076 11844
rect 27468 12460 27524 12516
rect 26572 10668 26628 10724
rect 25900 10332 25956 10388
rect 25788 9660 25844 9716
rect 25900 9212 25956 9268
rect 26236 9938 26292 9940
rect 26236 9886 26238 9938
rect 26238 9886 26290 9938
rect 26290 9886 26292 9938
rect 26236 9884 26292 9886
rect 26684 10556 26740 10612
rect 27020 10668 27076 10724
rect 27356 11676 27412 11732
rect 26796 9996 26852 10052
rect 25900 8764 25956 8820
rect 26124 8034 26180 8036
rect 26124 7982 26126 8034
rect 26126 7982 26178 8034
rect 26178 7982 26180 8034
rect 26124 7980 26180 7982
rect 26348 8540 26404 8596
rect 26796 9660 26852 9716
rect 25564 7308 25620 7364
rect 25004 6578 25060 6580
rect 25004 6526 25006 6578
rect 25006 6526 25058 6578
rect 25058 6526 25060 6578
rect 25004 6524 25060 6526
rect 24892 6412 24948 6468
rect 24780 6130 24836 6132
rect 24780 6078 24782 6130
rect 24782 6078 24834 6130
rect 24834 6078 24836 6130
rect 24780 6076 24836 6078
rect 24668 5234 24724 5236
rect 24668 5182 24670 5234
rect 24670 5182 24722 5234
rect 24722 5182 24724 5234
rect 24668 5180 24724 5182
rect 25228 5964 25284 6020
rect 25340 6188 25396 6244
rect 24668 4562 24724 4564
rect 24668 4510 24670 4562
rect 24670 4510 24722 4562
rect 24722 4510 24724 4562
rect 24668 4508 24724 4510
rect 25452 6412 25508 6468
rect 26796 9212 26852 9268
rect 26572 9042 26628 9044
rect 26572 8990 26574 9042
rect 26574 8990 26626 9042
rect 26626 8990 26628 9042
rect 26572 8988 26628 8990
rect 27356 10780 27412 10836
rect 27356 10220 27412 10276
rect 26572 7980 26628 8036
rect 26572 7756 26628 7812
rect 25676 6578 25732 6580
rect 25676 6526 25678 6578
rect 25678 6526 25730 6578
rect 25730 6526 25732 6578
rect 25676 6524 25732 6526
rect 25564 6188 25620 6244
rect 25900 5628 25956 5684
rect 25900 5292 25956 5348
rect 25452 4562 25508 4564
rect 25452 4510 25454 4562
rect 25454 4510 25506 4562
rect 25506 4510 25508 4562
rect 25452 4508 25508 4510
rect 26348 6524 26404 6580
rect 26796 6524 26852 6580
rect 26012 5068 26068 5124
rect 26124 4898 26180 4900
rect 26124 4846 26126 4898
rect 26126 4846 26178 4898
rect 26178 4846 26180 4898
rect 26124 4844 26180 4846
rect 26684 6188 26740 6244
rect 26796 5964 26852 6020
rect 27356 8258 27412 8260
rect 27356 8206 27358 8258
rect 27358 8206 27410 8258
rect 27410 8206 27412 8258
rect 27356 8204 27412 8206
rect 27132 8092 27188 8148
rect 28140 13916 28196 13972
rect 28028 12012 28084 12068
rect 27692 8876 27748 8932
rect 27692 8034 27748 8036
rect 27692 7982 27694 8034
rect 27694 7982 27746 8034
rect 27746 7982 27748 8034
rect 27692 7980 27748 7982
rect 27020 6860 27076 6916
rect 26684 5180 26740 5236
rect 26460 4844 26516 4900
rect 26684 4844 26740 4900
rect 26908 4508 26964 4564
rect 27020 5180 27076 5236
rect 28364 16098 28420 16100
rect 28364 16046 28366 16098
rect 28366 16046 28418 16098
rect 28418 16046 28420 16098
rect 28364 16044 28420 16046
rect 28364 14530 28420 14532
rect 28364 14478 28366 14530
rect 28366 14478 28418 14530
rect 28418 14478 28420 14530
rect 28364 14476 28420 14478
rect 28812 16044 28868 16100
rect 28700 15426 28756 15428
rect 28700 15374 28702 15426
rect 28702 15374 28754 15426
rect 28754 15374 28756 15426
rect 28700 15372 28756 15374
rect 28588 14252 28644 14308
rect 28252 12402 28308 12404
rect 28252 12350 28254 12402
rect 28254 12350 28306 12402
rect 28306 12350 28308 12402
rect 28252 12348 28308 12350
rect 28700 12572 28756 12628
rect 28140 11228 28196 11284
rect 28252 12124 28308 12180
rect 27916 10668 27972 10724
rect 27804 7644 27860 7700
rect 27244 6690 27300 6692
rect 27244 6638 27246 6690
rect 27246 6638 27298 6690
rect 27298 6638 27300 6690
rect 27244 6636 27300 6638
rect 27916 10220 27972 10276
rect 28700 11900 28756 11956
rect 28364 11618 28420 11620
rect 28364 11566 28366 11618
rect 28366 11566 28418 11618
rect 28418 11566 28420 11618
rect 28364 11564 28420 11566
rect 28588 10892 28644 10948
rect 28588 9996 28644 10052
rect 28252 9772 28308 9828
rect 28028 9100 28084 9156
rect 28140 8930 28196 8932
rect 28140 8878 28142 8930
rect 28142 8878 28194 8930
rect 28194 8878 28196 8930
rect 28140 8876 28196 8878
rect 28028 8540 28084 8596
rect 28364 9660 28420 9716
rect 29148 18172 29204 18228
rect 29260 18060 29316 18116
rect 29148 17388 29204 17444
rect 29148 15820 29204 15876
rect 29484 18396 29540 18452
rect 29596 18060 29652 18116
rect 29708 17836 29764 17892
rect 29708 16658 29764 16660
rect 29708 16606 29710 16658
rect 29710 16606 29762 16658
rect 29762 16606 29764 16658
rect 29708 16604 29764 16606
rect 29708 16380 29764 16436
rect 29932 16882 29988 16884
rect 29932 16830 29934 16882
rect 29934 16830 29986 16882
rect 29986 16830 29988 16882
rect 29932 16828 29988 16830
rect 29708 15484 29764 15540
rect 29260 14642 29316 14644
rect 29260 14590 29262 14642
rect 29262 14590 29314 14642
rect 29314 14590 29316 14642
rect 29260 14588 29316 14590
rect 29372 14476 29428 14532
rect 28924 12684 28980 12740
rect 29148 12572 29204 12628
rect 29372 12738 29428 12740
rect 29372 12686 29374 12738
rect 29374 12686 29426 12738
rect 29426 12686 29428 12738
rect 29372 12684 29428 12686
rect 29036 12460 29092 12516
rect 29036 11788 29092 11844
rect 29148 12348 29204 12404
rect 29260 11676 29316 11732
rect 29372 11340 29428 11396
rect 29372 9826 29428 9828
rect 29372 9774 29374 9826
rect 29374 9774 29426 9826
rect 29426 9774 29428 9826
rect 29372 9772 29428 9774
rect 28812 9266 28868 9268
rect 28812 9214 28814 9266
rect 28814 9214 28866 9266
rect 28866 9214 28868 9266
rect 28812 9212 28868 9214
rect 28700 9042 28756 9044
rect 28700 8990 28702 9042
rect 28702 8990 28754 9042
rect 28754 8990 28756 9042
rect 28700 8988 28756 8990
rect 28252 8428 28308 8484
rect 28700 8092 28756 8148
rect 28476 8034 28532 8036
rect 28476 7982 28478 8034
rect 28478 7982 28530 8034
rect 28530 7982 28532 8034
rect 28476 7980 28532 7982
rect 28364 7644 28420 7700
rect 28476 7586 28532 7588
rect 28476 7534 28478 7586
rect 28478 7534 28530 7586
rect 28530 7534 28532 7586
rect 28476 7532 28532 7534
rect 27692 6972 27748 7028
rect 28140 6636 28196 6692
rect 27580 6412 27636 6468
rect 27244 6300 27300 6356
rect 28476 7084 28532 7140
rect 28476 6524 28532 6580
rect 28140 6018 28196 6020
rect 28140 5966 28142 6018
rect 28142 5966 28194 6018
rect 28194 5966 28196 6018
rect 28140 5964 28196 5966
rect 28028 5068 28084 5124
rect 28364 5628 28420 5684
rect 28812 6412 28868 6468
rect 28476 6076 28532 6132
rect 27468 4620 27524 4676
rect 27916 4508 27972 4564
rect 27916 4338 27972 4340
rect 27916 4286 27918 4338
rect 27918 4286 27970 4338
rect 27970 4286 27972 4338
rect 27916 4284 27972 4286
rect 27468 3836 27524 3892
rect 27020 3724 27076 3780
rect 26124 3666 26180 3668
rect 26124 3614 26126 3666
rect 26126 3614 26178 3666
rect 26178 3614 26180 3666
rect 26124 3612 26180 3614
rect 25676 3554 25732 3556
rect 25676 3502 25678 3554
rect 25678 3502 25730 3554
rect 25730 3502 25732 3554
rect 25676 3500 25732 3502
rect 26572 3442 26628 3444
rect 26572 3390 26574 3442
rect 26574 3390 26626 3442
rect 26626 3390 26628 3442
rect 26572 3388 26628 3390
rect 29260 9212 29316 9268
rect 29596 14700 29652 14756
rect 29596 14306 29652 14308
rect 29596 14254 29598 14306
rect 29598 14254 29650 14306
rect 29650 14254 29652 14306
rect 29596 14252 29652 14254
rect 29708 12796 29764 12852
rect 29596 12236 29652 12292
rect 29596 11228 29652 11284
rect 29260 8540 29316 8596
rect 29148 7756 29204 7812
rect 29372 7474 29428 7476
rect 29372 7422 29374 7474
rect 29374 7422 29426 7474
rect 29426 7422 29428 7474
rect 29372 7420 29428 7422
rect 30380 20690 30436 20692
rect 30380 20638 30382 20690
rect 30382 20638 30434 20690
rect 30434 20638 30436 20690
rect 30380 20636 30436 20638
rect 30156 20300 30212 20356
rect 30940 21756 30996 21812
rect 30604 20524 30660 20580
rect 30492 20130 30548 20132
rect 30492 20078 30494 20130
rect 30494 20078 30546 20130
rect 30546 20078 30548 20130
rect 30492 20076 30548 20078
rect 30380 19628 30436 19684
rect 30156 19346 30212 19348
rect 30156 19294 30158 19346
rect 30158 19294 30210 19346
rect 30210 19294 30212 19346
rect 30156 19292 30212 19294
rect 30492 19068 30548 19124
rect 30492 18620 30548 18676
rect 30380 17778 30436 17780
rect 30380 17726 30382 17778
rect 30382 17726 30434 17778
rect 30434 17726 30436 17778
rect 30380 17724 30436 17726
rect 30156 16716 30212 16772
rect 30380 17106 30436 17108
rect 30380 17054 30382 17106
rect 30382 17054 30434 17106
rect 30434 17054 30436 17106
rect 30380 17052 30436 17054
rect 30044 15820 30100 15876
rect 30716 20412 30772 20468
rect 32508 27356 32564 27412
rect 32172 26124 32228 26180
rect 32396 25900 32452 25956
rect 33292 28588 33348 28644
rect 33404 27356 33460 27412
rect 33516 28028 33572 28084
rect 33404 27186 33460 27188
rect 33404 27134 33406 27186
rect 33406 27134 33458 27186
rect 33458 27134 33460 27186
rect 33404 27132 33460 27134
rect 33740 29820 33796 29876
rect 33628 27858 33684 27860
rect 33628 27806 33630 27858
rect 33630 27806 33682 27858
rect 33682 27806 33684 27858
rect 33628 27804 33684 27806
rect 33852 28700 33908 28756
rect 34188 30828 34244 30884
rect 34188 30604 34244 30660
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35532 31778 35588 31780
rect 35532 31726 35534 31778
rect 35534 31726 35586 31778
rect 35586 31726 35588 31778
rect 35532 31724 35588 31726
rect 35756 31500 35812 31556
rect 36092 32732 36148 32788
rect 35980 32284 36036 32340
rect 35980 31836 36036 31892
rect 36428 31724 36484 31780
rect 36316 31666 36372 31668
rect 36316 31614 36318 31666
rect 36318 31614 36370 31666
rect 36370 31614 36372 31666
rect 36316 31612 36372 31614
rect 36652 32956 36708 33012
rect 36540 30940 36596 30996
rect 35644 30716 35700 30772
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34412 30210 34468 30212
rect 34412 30158 34414 30210
rect 34414 30158 34466 30210
rect 34466 30158 34468 30210
rect 34412 30156 34468 30158
rect 34972 29932 35028 29988
rect 34300 28252 34356 28308
rect 34076 28082 34132 28084
rect 34076 28030 34078 28082
rect 34078 28030 34130 28082
rect 34130 28030 34132 28082
rect 34076 28028 34132 28030
rect 33740 27692 33796 27748
rect 32956 25900 33012 25956
rect 33068 26796 33124 26852
rect 32732 25116 32788 25172
rect 32060 24834 32116 24836
rect 32060 24782 32062 24834
rect 32062 24782 32114 24834
rect 32114 24782 32116 24834
rect 32060 24780 32116 24782
rect 31948 24556 32004 24612
rect 32172 24108 32228 24164
rect 31612 23938 31668 23940
rect 31612 23886 31614 23938
rect 31614 23886 31666 23938
rect 31666 23886 31668 23938
rect 31612 23884 31668 23886
rect 31500 22764 31556 22820
rect 31164 21532 31220 21588
rect 31276 22652 31332 22708
rect 31500 22370 31556 22372
rect 31500 22318 31502 22370
rect 31502 22318 31554 22370
rect 31554 22318 31556 22370
rect 31500 22316 31556 22318
rect 31388 21362 31444 21364
rect 31388 21310 31390 21362
rect 31390 21310 31442 21362
rect 31442 21310 31444 21362
rect 31388 21308 31444 21310
rect 31612 21084 31668 21140
rect 32172 22652 32228 22708
rect 32284 23884 32340 23940
rect 32060 22540 32116 22596
rect 32060 21980 32116 22036
rect 31836 21756 31892 21812
rect 32172 21868 32228 21924
rect 33180 23266 33236 23268
rect 33180 23214 33182 23266
rect 33182 23214 33234 23266
rect 33234 23214 33236 23266
rect 33180 23212 33236 23214
rect 33068 22652 33124 22708
rect 32732 22428 32788 22484
rect 33404 24834 33460 24836
rect 33404 24782 33406 24834
rect 33406 24782 33458 24834
rect 33458 24782 33460 24834
rect 33404 24780 33460 24782
rect 33516 24444 33572 24500
rect 33516 23938 33572 23940
rect 33516 23886 33518 23938
rect 33518 23886 33570 23938
rect 33570 23886 33572 23938
rect 33516 23884 33572 23886
rect 33292 22428 33348 22484
rect 33404 23548 33460 23604
rect 32284 22204 32340 22260
rect 33068 22258 33124 22260
rect 33068 22206 33070 22258
rect 33070 22206 33122 22258
rect 33122 22206 33124 22258
rect 33068 22204 33124 22206
rect 32396 21756 32452 21812
rect 32732 21868 32788 21924
rect 30940 20578 30996 20580
rect 30940 20526 30942 20578
rect 30942 20526 30994 20578
rect 30994 20526 30996 20578
rect 30940 20524 30996 20526
rect 31500 20524 31556 20580
rect 31052 20300 31108 20356
rect 30940 20188 30996 20244
rect 30716 18450 30772 18452
rect 30716 18398 30718 18450
rect 30718 18398 30770 18450
rect 30770 18398 30772 18450
rect 30716 18396 30772 18398
rect 30940 18396 30996 18452
rect 30828 17666 30884 17668
rect 30828 17614 30830 17666
rect 30830 17614 30882 17666
rect 30882 17614 30884 17666
rect 30828 17612 30884 17614
rect 31164 20076 31220 20132
rect 32620 21308 32676 21364
rect 32060 21084 32116 21140
rect 31948 20914 32004 20916
rect 31948 20862 31950 20914
rect 31950 20862 32002 20914
rect 32002 20862 32004 20914
rect 31948 20860 32004 20862
rect 32396 20802 32452 20804
rect 32396 20750 32398 20802
rect 32398 20750 32450 20802
rect 32450 20750 32452 20802
rect 32396 20748 32452 20750
rect 32508 20636 32564 20692
rect 33068 21308 33124 21364
rect 33292 21810 33348 21812
rect 33292 21758 33294 21810
rect 33294 21758 33346 21810
rect 33346 21758 33348 21810
rect 33292 21756 33348 21758
rect 33292 21586 33348 21588
rect 33292 21534 33294 21586
rect 33294 21534 33346 21586
rect 33346 21534 33348 21586
rect 33292 21532 33348 21534
rect 33068 21084 33124 21140
rect 34188 27692 34244 27748
rect 34076 27244 34132 27300
rect 33964 26962 34020 26964
rect 33964 26910 33966 26962
rect 33966 26910 34018 26962
rect 34018 26910 34020 26962
rect 33964 26908 34020 26910
rect 34076 25788 34132 25844
rect 34524 29538 34580 29540
rect 34524 29486 34526 29538
rect 34526 29486 34578 29538
rect 34578 29486 34580 29538
rect 34524 29484 34580 29486
rect 34636 28418 34692 28420
rect 34636 28366 34638 28418
rect 34638 28366 34690 28418
rect 34690 28366 34692 28418
rect 34636 28364 34692 28366
rect 35084 29484 35140 29540
rect 35308 29484 35364 29540
rect 35532 29596 35588 29652
rect 34748 28252 34804 28308
rect 35084 29260 35140 29316
rect 35756 29986 35812 29988
rect 35756 29934 35758 29986
rect 35758 29934 35810 29986
rect 35810 29934 35812 29986
rect 35756 29932 35812 29934
rect 35868 29820 35924 29876
rect 35980 29596 36036 29652
rect 35644 29260 35700 29316
rect 35196 29148 35252 29204
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 28812 35252 28868
rect 35196 28588 35252 28644
rect 35868 28812 35924 28868
rect 34972 28364 35028 28420
rect 35532 28252 35588 28308
rect 35532 27858 35588 27860
rect 35532 27806 35534 27858
rect 35534 27806 35586 27858
rect 35586 27806 35588 27858
rect 35532 27804 35588 27806
rect 35980 28642 36036 28644
rect 35980 28590 35982 28642
rect 35982 28590 36034 28642
rect 36034 28590 36036 28642
rect 35980 28588 36036 28590
rect 36204 29036 36260 29092
rect 36092 28252 36148 28308
rect 36204 28364 36260 28420
rect 34860 27132 34916 27188
rect 34524 26962 34580 26964
rect 34524 26910 34526 26962
rect 34526 26910 34578 26962
rect 34578 26910 34580 26962
rect 34524 26908 34580 26910
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35868 27468 35924 27524
rect 35756 27074 35812 27076
rect 35756 27022 35758 27074
rect 35758 27022 35810 27074
rect 35810 27022 35812 27074
rect 35756 27020 35812 27022
rect 35196 26962 35252 26964
rect 35196 26910 35198 26962
rect 35198 26910 35250 26962
rect 35250 26910 35252 26962
rect 35196 26908 35252 26910
rect 34524 26290 34580 26292
rect 34524 26238 34526 26290
rect 34526 26238 34578 26290
rect 34578 26238 34580 26290
rect 34524 26236 34580 26238
rect 34748 26178 34804 26180
rect 34748 26126 34750 26178
rect 34750 26126 34802 26178
rect 34802 26126 34804 26178
rect 34748 26124 34804 26126
rect 34300 25564 34356 25620
rect 34412 25228 34468 25284
rect 34300 24108 34356 24164
rect 33852 23212 33908 23268
rect 33516 21980 33572 22036
rect 33964 22316 34020 22372
rect 34188 23212 34244 23268
rect 34524 22764 34580 22820
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35084 25564 35140 25620
rect 35420 25506 35476 25508
rect 35420 25454 35422 25506
rect 35422 25454 35474 25506
rect 35474 25454 35476 25506
rect 35420 25452 35476 25454
rect 35084 25394 35140 25396
rect 35084 25342 35086 25394
rect 35086 25342 35138 25394
rect 35138 25342 35140 25394
rect 35084 25340 35140 25342
rect 34748 24892 34804 24948
rect 34524 22540 34580 22596
rect 34300 21474 34356 21476
rect 34300 21422 34302 21474
rect 34302 21422 34354 21474
rect 34354 21422 34356 21474
rect 34300 21420 34356 21422
rect 33852 20860 33908 20916
rect 32620 20412 32676 20468
rect 32508 20188 32564 20244
rect 31948 19292 32004 19348
rect 32732 19852 32788 19908
rect 32732 18508 32788 18564
rect 32396 18450 32452 18452
rect 32396 18398 32398 18450
rect 32398 18398 32450 18450
rect 32450 18398 32452 18450
rect 32396 18396 32452 18398
rect 31052 17612 31108 17668
rect 31948 17612 32004 17668
rect 32396 17554 32452 17556
rect 32396 17502 32398 17554
rect 32398 17502 32450 17554
rect 32450 17502 32452 17554
rect 32396 17500 32452 17502
rect 32172 17388 32228 17444
rect 30828 16716 30884 16772
rect 30716 16604 30772 16660
rect 30716 15538 30772 15540
rect 30716 15486 30718 15538
rect 30718 15486 30770 15538
rect 30770 15486 30772 15538
rect 30716 15484 30772 15486
rect 30492 15260 30548 15316
rect 31500 15372 31556 15428
rect 30604 14700 30660 14756
rect 29932 13746 29988 13748
rect 29932 13694 29934 13746
rect 29934 13694 29986 13746
rect 29986 13694 29988 13746
rect 29932 13692 29988 13694
rect 30156 14418 30212 14420
rect 30156 14366 30158 14418
rect 30158 14366 30210 14418
rect 30210 14366 30212 14418
rect 30156 14364 30212 14366
rect 30380 14252 30436 14308
rect 30044 13468 30100 13524
rect 30268 13020 30324 13076
rect 29932 12572 29988 12628
rect 29932 12402 29988 12404
rect 29932 12350 29934 12402
rect 29934 12350 29986 12402
rect 29986 12350 29988 12402
rect 29932 12348 29988 12350
rect 30268 12012 30324 12068
rect 29932 11676 29988 11732
rect 31164 14754 31220 14756
rect 31164 14702 31166 14754
rect 31166 14702 31218 14754
rect 31218 14702 31220 14754
rect 31164 14700 31220 14702
rect 30716 13468 30772 13524
rect 30828 13244 30884 13300
rect 30940 13692 30996 13748
rect 30604 13020 30660 13076
rect 30604 12850 30660 12852
rect 30604 12798 30606 12850
rect 30606 12798 30658 12850
rect 30658 12798 30660 12850
rect 30604 12796 30660 12798
rect 30604 12178 30660 12180
rect 30604 12126 30606 12178
rect 30606 12126 30658 12178
rect 30658 12126 30660 12178
rect 30604 12124 30660 12126
rect 30604 11618 30660 11620
rect 30604 11566 30606 11618
rect 30606 11566 30658 11618
rect 30658 11566 30660 11618
rect 30604 11564 30660 11566
rect 30828 11564 30884 11620
rect 29708 9436 29764 9492
rect 29932 9714 29988 9716
rect 29932 9662 29934 9714
rect 29934 9662 29986 9714
rect 29986 9662 29988 9714
rect 29932 9660 29988 9662
rect 29820 9212 29876 9268
rect 29708 8092 29764 8148
rect 29932 7644 29988 7700
rect 29148 5794 29204 5796
rect 29148 5742 29150 5794
rect 29150 5742 29202 5794
rect 29202 5742 29204 5794
rect 29148 5740 29204 5742
rect 29260 4562 29316 4564
rect 29260 4510 29262 4562
rect 29262 4510 29314 4562
rect 29314 4510 29316 4562
rect 29260 4508 29316 4510
rect 29596 6578 29652 6580
rect 29596 6526 29598 6578
rect 29598 6526 29650 6578
rect 29650 6526 29652 6578
rect 29596 6524 29652 6526
rect 30716 10610 30772 10612
rect 30716 10558 30718 10610
rect 30718 10558 30770 10610
rect 30770 10558 30772 10610
rect 30716 10556 30772 10558
rect 30492 9996 30548 10052
rect 30268 9324 30324 9380
rect 30268 8930 30324 8932
rect 30268 8878 30270 8930
rect 30270 8878 30322 8930
rect 30322 8878 30324 8930
rect 30268 8876 30324 8878
rect 31164 13468 31220 13524
rect 31388 13244 31444 13300
rect 31276 12962 31332 12964
rect 31276 12910 31278 12962
rect 31278 12910 31330 12962
rect 31330 12910 31332 12962
rect 31276 12908 31332 12910
rect 31164 12684 31220 12740
rect 31052 12348 31108 12404
rect 31276 12236 31332 12292
rect 31388 11116 31444 11172
rect 32060 16994 32116 16996
rect 32060 16942 32062 16994
rect 32062 16942 32114 16994
rect 32114 16942 32116 16994
rect 32060 16940 32116 16942
rect 31948 16828 32004 16884
rect 31612 15932 31668 15988
rect 31612 14588 31668 14644
rect 32284 14530 32340 14532
rect 32284 14478 32286 14530
rect 32286 14478 32338 14530
rect 32338 14478 32340 14530
rect 32284 14476 32340 14478
rect 31836 14252 31892 14308
rect 32284 13970 32340 13972
rect 32284 13918 32286 13970
rect 32286 13918 32338 13970
rect 32338 13918 32340 13970
rect 32284 13916 32340 13918
rect 31724 13692 31780 13748
rect 31836 12908 31892 12964
rect 31836 12012 31892 12068
rect 32620 12796 32676 12852
rect 32956 20188 33012 20244
rect 33516 19964 33572 20020
rect 33292 19404 33348 19460
rect 34188 20018 34244 20020
rect 34188 19966 34190 20018
rect 34190 19966 34242 20018
rect 34242 19966 34244 20018
rect 34188 19964 34244 19966
rect 33852 19292 33908 19348
rect 34188 19234 34244 19236
rect 34188 19182 34190 19234
rect 34190 19182 34242 19234
rect 34242 19182 34244 19234
rect 34188 19180 34244 19182
rect 33068 18450 33124 18452
rect 33068 18398 33070 18450
rect 33070 18398 33122 18450
rect 33122 18398 33124 18450
rect 33068 18396 33124 18398
rect 33516 17836 33572 17892
rect 33740 18284 33796 18340
rect 33292 17052 33348 17108
rect 32956 16380 33012 16436
rect 33068 15986 33124 15988
rect 33068 15934 33070 15986
rect 33070 15934 33122 15986
rect 33122 15934 33124 15986
rect 33068 15932 33124 15934
rect 33516 16156 33572 16212
rect 33628 16604 33684 16660
rect 33180 15426 33236 15428
rect 33180 15374 33182 15426
rect 33182 15374 33234 15426
rect 33234 15374 33236 15426
rect 33180 15372 33236 15374
rect 33628 15708 33684 15764
rect 32956 14924 33012 14980
rect 33068 14700 33124 14756
rect 33404 14754 33460 14756
rect 33404 14702 33406 14754
rect 33406 14702 33458 14754
rect 33458 14702 33460 14754
rect 33404 14700 33460 14702
rect 33068 14364 33124 14420
rect 33404 14364 33460 14420
rect 33404 13858 33460 13860
rect 33404 13806 33406 13858
rect 33406 13806 33458 13858
rect 33458 13806 33460 13858
rect 33404 13804 33460 13806
rect 33292 13746 33348 13748
rect 33292 13694 33294 13746
rect 33294 13694 33346 13746
rect 33346 13694 33348 13746
rect 33292 13692 33348 13694
rect 33292 12460 33348 12516
rect 33852 18172 33908 18228
rect 34076 19068 34132 19124
rect 34300 18956 34356 19012
rect 34076 18396 34132 18452
rect 34524 21644 34580 21700
rect 35868 26908 35924 26964
rect 35756 25452 35812 25508
rect 35756 25282 35812 25284
rect 35756 25230 35758 25282
rect 35758 25230 35810 25282
rect 35810 25230 35812 25282
rect 35756 25228 35812 25230
rect 35532 24668 35588 24724
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35084 24108 35140 24164
rect 34860 23714 34916 23716
rect 34860 23662 34862 23714
rect 34862 23662 34914 23714
rect 34914 23662 34916 23714
rect 34860 23660 34916 23662
rect 35084 23660 35140 23716
rect 34748 21532 34804 21588
rect 35420 23100 35476 23156
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 22540 35252 22596
rect 35756 23884 35812 23940
rect 36092 23660 36148 23716
rect 35868 23266 35924 23268
rect 35868 23214 35870 23266
rect 35870 23214 35922 23266
rect 35922 23214 35924 23266
rect 35868 23212 35924 23214
rect 36092 23154 36148 23156
rect 36092 23102 36094 23154
rect 36094 23102 36146 23154
rect 36146 23102 36148 23154
rect 36092 23100 36148 23102
rect 35868 22876 35924 22932
rect 35532 21644 35588 21700
rect 35756 21586 35812 21588
rect 35756 21534 35758 21586
rect 35758 21534 35810 21586
rect 35810 21534 35812 21586
rect 35756 21532 35812 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34972 20748 35028 20804
rect 35084 20636 35140 20692
rect 35308 20188 35364 20244
rect 34748 20076 34804 20132
rect 34972 20076 35028 20132
rect 35756 20076 35812 20132
rect 35196 19852 35252 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34972 19292 35028 19348
rect 35420 19292 35476 19348
rect 34748 18620 34804 18676
rect 35084 18450 35140 18452
rect 35084 18398 35086 18450
rect 35086 18398 35138 18450
rect 35138 18398 35140 18450
rect 35084 18396 35140 18398
rect 35196 18284 35252 18340
rect 34412 17052 34468 17108
rect 34524 17724 34580 17780
rect 35420 18172 35476 18228
rect 35532 18732 35588 18788
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 36652 29650 36708 29652
rect 36652 29598 36654 29650
rect 36654 29598 36706 29650
rect 36706 29598 36708 29650
rect 36652 29596 36708 29598
rect 36540 29538 36596 29540
rect 36540 29486 36542 29538
rect 36542 29486 36594 29538
rect 36594 29486 36596 29538
rect 36540 29484 36596 29486
rect 36428 29372 36484 29428
rect 37212 36876 37268 36932
rect 37100 35644 37156 35700
rect 36876 34636 36932 34692
rect 37212 34524 37268 34580
rect 37436 36988 37492 37044
rect 40572 51548 40628 51604
rect 40572 49868 40628 49924
rect 40908 53058 40964 53060
rect 40908 53006 40910 53058
rect 40910 53006 40962 53058
rect 40962 53006 40964 53058
rect 40908 53004 40964 53006
rect 41356 53788 41412 53844
rect 44044 57260 44100 57316
rect 42252 56754 42308 56756
rect 42252 56702 42254 56754
rect 42254 56702 42306 56754
rect 42306 56702 42308 56754
rect 42252 56700 42308 56702
rect 42588 56252 42644 56308
rect 42252 55692 42308 55748
rect 41132 53228 41188 53284
rect 40796 50316 40852 50372
rect 40796 49756 40852 49812
rect 40684 47628 40740 47684
rect 41020 52050 41076 52052
rect 41020 51998 41022 52050
rect 41022 51998 41074 52050
rect 41074 51998 41076 52050
rect 41020 51996 41076 51998
rect 41244 50594 41300 50596
rect 41244 50542 41246 50594
rect 41246 50542 41298 50594
rect 41298 50542 41300 50594
rect 41244 50540 41300 50542
rect 41020 50482 41076 50484
rect 41020 50430 41022 50482
rect 41022 50430 41074 50482
rect 41074 50430 41076 50482
rect 41020 50428 41076 50430
rect 41132 49196 41188 49252
rect 41692 51436 41748 51492
rect 41692 50706 41748 50708
rect 41692 50654 41694 50706
rect 41694 50654 41746 50706
rect 41746 50654 41748 50706
rect 41692 50652 41748 50654
rect 41916 53228 41972 53284
rect 42588 55298 42644 55300
rect 42588 55246 42590 55298
rect 42590 55246 42642 55298
rect 42642 55246 42644 55298
rect 42588 55244 42644 55246
rect 42252 54684 42308 54740
rect 42140 54402 42196 54404
rect 42140 54350 42142 54402
rect 42142 54350 42194 54402
rect 42194 54350 42196 54402
rect 42140 54348 42196 54350
rect 42252 53676 42308 53732
rect 42812 56252 42868 56308
rect 43596 55916 43652 55972
rect 42924 55186 42980 55188
rect 42924 55134 42926 55186
rect 42926 55134 42978 55186
rect 42978 55134 42980 55186
rect 42924 55132 42980 55134
rect 43372 54012 43428 54068
rect 42700 53676 42756 53732
rect 42364 53340 42420 53396
rect 42812 53340 42868 53396
rect 42028 52332 42084 52388
rect 42700 52332 42756 52388
rect 41356 49644 41412 49700
rect 41468 48748 41524 48804
rect 41132 48636 41188 48692
rect 41580 48354 41636 48356
rect 41580 48302 41582 48354
rect 41582 48302 41634 48354
rect 41634 48302 41636 48354
rect 41580 48300 41636 48302
rect 41580 47682 41636 47684
rect 41580 47630 41582 47682
rect 41582 47630 41634 47682
rect 41634 47630 41636 47682
rect 41580 47628 41636 47630
rect 40236 46844 40292 46900
rect 38780 45052 38836 45108
rect 39004 46396 39060 46452
rect 39676 46114 39732 46116
rect 39676 46062 39678 46114
rect 39678 46062 39730 46114
rect 39730 46062 39732 46114
rect 39676 46060 39732 46062
rect 39004 45724 39060 45780
rect 38444 43596 38500 43652
rect 38556 43538 38612 43540
rect 38556 43486 38558 43538
rect 38558 43486 38610 43538
rect 38610 43486 38612 43538
rect 38556 43484 38612 43486
rect 38556 42588 38612 42644
rect 38444 41916 38500 41972
rect 38892 42754 38948 42756
rect 38892 42702 38894 42754
rect 38894 42702 38946 42754
rect 38946 42702 38948 42754
rect 38892 42700 38948 42702
rect 39228 45106 39284 45108
rect 39228 45054 39230 45106
rect 39230 45054 39282 45106
rect 39282 45054 39284 45106
rect 39228 45052 39284 45054
rect 39900 44882 39956 44884
rect 39900 44830 39902 44882
rect 39902 44830 39954 44882
rect 39954 44830 39956 44882
rect 39900 44828 39956 44830
rect 39676 44492 39732 44548
rect 39116 43484 39172 43540
rect 39564 44380 39620 44436
rect 40460 46732 40516 46788
rect 40236 45388 40292 45444
rect 40348 45052 40404 45108
rect 40124 44604 40180 44660
rect 40236 44940 40292 44996
rect 40124 44434 40180 44436
rect 40124 44382 40126 44434
rect 40126 44382 40178 44434
rect 40178 44382 40180 44434
rect 40124 44380 40180 44382
rect 40124 43820 40180 43876
rect 39900 43036 39956 43092
rect 39340 42588 39396 42644
rect 38444 40962 38500 40964
rect 38444 40910 38446 40962
rect 38446 40910 38498 40962
rect 38498 40910 38500 40962
rect 38444 40908 38500 40910
rect 38332 40460 38388 40516
rect 38220 39452 38276 39508
rect 38668 39788 38724 39844
rect 39676 40908 39732 40964
rect 39788 40796 39844 40852
rect 40348 44492 40404 44548
rect 40908 46786 40964 46788
rect 40908 46734 40910 46786
rect 40910 46734 40962 46786
rect 40962 46734 40964 46786
rect 40908 46732 40964 46734
rect 40796 46508 40852 46564
rect 41804 47458 41860 47460
rect 41804 47406 41806 47458
rect 41806 47406 41858 47458
rect 41858 47406 41860 47458
rect 41804 47404 41860 47406
rect 41916 46956 41972 47012
rect 43036 52332 43092 52388
rect 43148 52274 43204 52276
rect 43148 52222 43150 52274
rect 43150 52222 43202 52274
rect 43202 52222 43204 52274
rect 43148 52220 43204 52222
rect 42812 50540 42868 50596
rect 43036 51996 43092 52052
rect 43148 51602 43204 51604
rect 43148 51550 43150 51602
rect 43150 51550 43202 51602
rect 43202 51550 43204 51602
rect 43148 51548 43204 51550
rect 42140 49868 42196 49924
rect 42364 49026 42420 49028
rect 42364 48974 42366 49026
rect 42366 48974 42418 49026
rect 42418 48974 42420 49026
rect 42364 48972 42420 48974
rect 42028 48412 42084 48468
rect 41132 46450 41188 46452
rect 41132 46398 41134 46450
rect 41134 46398 41186 46450
rect 41186 46398 41188 46450
rect 41132 46396 41188 46398
rect 41132 45164 41188 45220
rect 41020 44434 41076 44436
rect 41020 44382 41022 44434
rect 41022 44382 41074 44434
rect 41074 44382 41076 44434
rect 41020 44380 41076 44382
rect 40908 43650 40964 43652
rect 40908 43598 40910 43650
rect 40910 43598 40962 43650
rect 40962 43598 40964 43650
rect 40908 43596 40964 43598
rect 40796 43484 40852 43540
rect 40236 43148 40292 43204
rect 40236 42754 40292 42756
rect 40236 42702 40238 42754
rect 40238 42702 40290 42754
rect 40290 42702 40292 42754
rect 40236 42700 40292 42702
rect 41132 43036 41188 43092
rect 41020 42978 41076 42980
rect 41020 42926 41022 42978
rect 41022 42926 41074 42978
rect 41074 42926 41076 42978
rect 41020 42924 41076 42926
rect 40908 42028 40964 42084
rect 40572 41074 40628 41076
rect 40572 41022 40574 41074
rect 40574 41022 40626 41074
rect 40626 41022 40628 41074
rect 40572 41020 40628 41022
rect 39564 40012 39620 40068
rect 39228 39788 39284 39844
rect 40908 40962 40964 40964
rect 40908 40910 40910 40962
rect 40910 40910 40962 40962
rect 40962 40910 40964 40962
rect 40908 40908 40964 40910
rect 40460 40572 40516 40628
rect 40796 40796 40852 40852
rect 40348 40236 40404 40292
rect 37884 37212 37940 37268
rect 37996 36876 38052 36932
rect 37772 36482 37828 36484
rect 37772 36430 37774 36482
rect 37774 36430 37826 36482
rect 37826 36430 37828 36482
rect 37772 36428 37828 36430
rect 37884 36204 37940 36260
rect 37996 35756 38052 35812
rect 38108 35980 38164 36036
rect 37436 35644 37492 35700
rect 37548 34914 37604 34916
rect 37548 34862 37550 34914
rect 37550 34862 37602 34914
rect 37602 34862 37604 34914
rect 37548 34860 37604 34862
rect 38220 34860 38276 34916
rect 38332 36204 38388 36260
rect 37324 34412 37380 34468
rect 37212 34076 37268 34132
rect 37100 33852 37156 33908
rect 36988 33122 37044 33124
rect 36988 33070 36990 33122
rect 36990 33070 37042 33122
rect 37042 33070 37044 33122
rect 36988 33068 37044 33070
rect 37100 32284 37156 32340
rect 37100 30940 37156 30996
rect 37548 33740 37604 33796
rect 38556 35756 38612 35812
rect 39452 37660 39508 37716
rect 38780 37154 38836 37156
rect 38780 37102 38782 37154
rect 38782 37102 38834 37154
rect 38834 37102 38836 37154
rect 38780 37100 38836 37102
rect 38780 35698 38836 35700
rect 38780 35646 38782 35698
rect 38782 35646 38834 35698
rect 38834 35646 38836 35698
rect 38780 35644 38836 35646
rect 39340 35084 39396 35140
rect 37884 33964 37940 34020
rect 37996 34076 38052 34132
rect 38220 33740 38276 33796
rect 37660 32508 37716 32564
rect 37436 31836 37492 31892
rect 37324 31666 37380 31668
rect 37324 31614 37326 31666
rect 37326 31614 37378 31666
rect 37378 31614 37380 31666
rect 37324 31612 37380 31614
rect 37772 33068 37828 33124
rect 37996 32620 38052 32676
rect 37884 32396 37940 32452
rect 38220 33346 38276 33348
rect 38220 33294 38222 33346
rect 38222 33294 38274 33346
rect 38274 33294 38276 33346
rect 38220 33292 38276 33294
rect 38668 34412 38724 34468
rect 38892 34412 38948 34468
rect 39340 34188 39396 34244
rect 38892 33964 38948 34020
rect 39340 33906 39396 33908
rect 39340 33854 39342 33906
rect 39342 33854 39394 33906
rect 39394 33854 39396 33906
rect 39340 33852 39396 33854
rect 39788 37436 39844 37492
rect 39676 37378 39732 37380
rect 39676 37326 39678 37378
rect 39678 37326 39730 37378
rect 39730 37326 39732 37378
rect 39676 37324 39732 37326
rect 39676 36988 39732 37044
rect 40012 39788 40068 39844
rect 40460 39394 40516 39396
rect 40460 39342 40462 39394
rect 40462 39342 40514 39394
rect 40514 39342 40516 39394
rect 40460 39340 40516 39342
rect 40348 38946 40404 38948
rect 40348 38894 40350 38946
rect 40350 38894 40402 38946
rect 40402 38894 40404 38946
rect 40348 38892 40404 38894
rect 40908 40460 40964 40516
rect 40348 37772 40404 37828
rect 41468 44940 41524 44996
rect 41692 46620 41748 46676
rect 42364 48524 42420 48580
rect 42028 46284 42084 46340
rect 42140 48076 42196 48132
rect 41692 45724 41748 45780
rect 41356 43932 41412 43988
rect 41580 43820 41636 43876
rect 41692 43538 41748 43540
rect 41692 43486 41694 43538
rect 41694 43486 41746 43538
rect 41746 43486 41748 43538
rect 41692 43484 41748 43486
rect 42140 45948 42196 46004
rect 42140 45500 42196 45556
rect 42812 49810 42868 49812
rect 42812 49758 42814 49810
rect 42814 49758 42866 49810
rect 42866 49758 42868 49810
rect 42812 49756 42868 49758
rect 42700 49250 42756 49252
rect 42700 49198 42702 49250
rect 42702 49198 42754 49250
rect 42754 49198 42756 49250
rect 42700 49196 42756 49198
rect 44268 56588 44324 56644
rect 43708 53730 43764 53732
rect 43708 53678 43710 53730
rect 43710 53678 43762 53730
rect 43762 53678 43764 53730
rect 43708 53676 43764 53678
rect 43932 55074 43988 55076
rect 43932 55022 43934 55074
rect 43934 55022 43986 55074
rect 43986 55022 43988 55074
rect 43932 55020 43988 55022
rect 43932 53788 43988 53844
rect 44268 53730 44324 53732
rect 44268 53678 44270 53730
rect 44270 53678 44322 53730
rect 44322 53678 44324 53730
rect 44268 53676 44324 53678
rect 44044 52892 44100 52948
rect 43708 52444 43764 52500
rect 43708 51548 43764 51604
rect 44940 57260 44996 57316
rect 44716 56476 44772 56532
rect 45612 58210 45668 58212
rect 45612 58158 45614 58210
rect 45614 58158 45666 58210
rect 45666 58158 45668 58210
rect 45612 58156 45668 58158
rect 46060 58210 46116 58212
rect 46060 58158 46062 58210
rect 46062 58158 46114 58210
rect 46114 58158 46116 58210
rect 46060 58156 46116 58158
rect 45164 56700 45220 56756
rect 45500 56476 45556 56532
rect 44492 54572 44548 54628
rect 45052 55580 45108 55636
rect 44716 55132 44772 55188
rect 45388 55356 45444 55412
rect 45836 56754 45892 56756
rect 45836 56702 45838 56754
rect 45838 56702 45890 56754
rect 45890 56702 45892 56754
rect 45836 56700 45892 56702
rect 46172 56642 46228 56644
rect 46172 56590 46174 56642
rect 46174 56590 46226 56642
rect 46226 56590 46228 56642
rect 46172 56588 46228 56590
rect 45948 56476 46004 56532
rect 46172 55410 46228 55412
rect 46172 55358 46174 55410
rect 46174 55358 46226 55410
rect 46226 55358 46228 55410
rect 46172 55356 46228 55358
rect 45612 54626 45668 54628
rect 45612 54574 45614 54626
rect 45614 54574 45666 54626
rect 45666 54574 45668 54626
rect 45612 54572 45668 54574
rect 45388 54460 45444 54516
rect 44940 54348 44996 54404
rect 44716 53340 44772 53396
rect 44604 52834 44660 52836
rect 44604 52782 44606 52834
rect 44606 52782 44658 52834
rect 44658 52782 44660 52834
rect 44604 52780 44660 52782
rect 44604 52556 44660 52612
rect 43820 51100 43876 51156
rect 43484 49980 43540 50036
rect 42588 48242 42644 48244
rect 42588 48190 42590 48242
rect 42590 48190 42642 48242
rect 42642 48190 42644 48242
rect 42588 48188 42644 48190
rect 42700 47516 42756 47572
rect 43372 49532 43428 49588
rect 43260 48914 43316 48916
rect 43260 48862 43262 48914
rect 43262 48862 43314 48914
rect 43314 48862 43316 48914
rect 43260 48860 43316 48862
rect 43148 48524 43204 48580
rect 43260 48636 43316 48692
rect 43036 48130 43092 48132
rect 43036 48078 43038 48130
rect 43038 48078 43090 48130
rect 43090 48078 43092 48130
rect 43036 48076 43092 48078
rect 42588 47346 42644 47348
rect 42588 47294 42590 47346
rect 42590 47294 42642 47346
rect 42642 47294 42644 47346
rect 42588 47292 42644 47294
rect 43148 47068 43204 47124
rect 42812 46956 42868 47012
rect 43484 48860 43540 48916
rect 43372 48188 43428 48244
rect 43596 48076 43652 48132
rect 43484 47404 43540 47460
rect 43372 47346 43428 47348
rect 43372 47294 43374 47346
rect 43374 47294 43426 47346
rect 43426 47294 43428 47346
rect 43372 47292 43428 47294
rect 43820 48748 43876 48804
rect 43708 47740 43764 47796
rect 43260 46844 43316 46900
rect 43372 46508 43428 46564
rect 43260 45500 43316 45556
rect 43260 45276 43316 45332
rect 43372 45164 43428 45220
rect 41356 41916 41412 41972
rect 41468 42028 41524 42084
rect 41468 41020 41524 41076
rect 42812 44210 42868 44212
rect 42812 44158 42814 44210
rect 42814 44158 42866 44210
rect 42866 44158 42868 44210
rect 42812 44156 42868 44158
rect 42252 43762 42308 43764
rect 42252 43710 42254 43762
rect 42254 43710 42306 43762
rect 42306 43710 42308 43762
rect 42252 43708 42308 43710
rect 42140 42700 42196 42756
rect 41916 42194 41972 42196
rect 41916 42142 41918 42194
rect 41918 42142 41970 42194
rect 41970 42142 41972 42194
rect 41916 42140 41972 42142
rect 42028 42028 42084 42084
rect 42252 43484 42308 43540
rect 41244 40572 41300 40628
rect 41132 39506 41188 39508
rect 41132 39454 41134 39506
rect 41134 39454 41186 39506
rect 41186 39454 41188 39506
rect 41132 39452 41188 39454
rect 41132 39058 41188 39060
rect 41132 39006 41134 39058
rect 41134 39006 41186 39058
rect 41186 39006 41188 39058
rect 41132 39004 41188 39006
rect 41356 38946 41412 38948
rect 41356 38894 41358 38946
rect 41358 38894 41410 38946
rect 41410 38894 41412 38946
rect 41356 38892 41412 38894
rect 41244 38722 41300 38724
rect 41244 38670 41246 38722
rect 41246 38670 41298 38722
rect 41298 38670 41300 38722
rect 41244 38668 41300 38670
rect 41580 38780 41636 38836
rect 41468 38220 41524 38276
rect 42028 40460 42084 40516
rect 42028 39116 42084 39172
rect 42140 38556 42196 38612
rect 41804 38444 41860 38500
rect 42028 38332 42084 38388
rect 41020 37266 41076 37268
rect 41020 37214 41022 37266
rect 41022 37214 41074 37266
rect 41074 37214 41076 37266
rect 41020 37212 41076 37214
rect 40348 37100 40404 37156
rect 41132 37100 41188 37156
rect 39788 36540 39844 36596
rect 39564 35308 39620 35364
rect 39564 34914 39620 34916
rect 39564 34862 39566 34914
rect 39566 34862 39618 34914
rect 39618 34862 39620 34914
rect 39564 34860 39620 34862
rect 39788 36316 39844 36372
rect 39900 35868 39956 35924
rect 40124 36092 40180 36148
rect 39788 35810 39844 35812
rect 39788 35758 39790 35810
rect 39790 35758 39842 35810
rect 39842 35758 39844 35810
rect 39788 35756 39844 35758
rect 39900 35308 39956 35364
rect 41020 36764 41076 36820
rect 40684 35868 40740 35924
rect 40348 35810 40404 35812
rect 40348 35758 40350 35810
rect 40350 35758 40402 35810
rect 40402 35758 40404 35810
rect 40348 35756 40404 35758
rect 40124 35308 40180 35364
rect 40012 34860 40068 34916
rect 39900 34412 39956 34468
rect 39788 34188 39844 34244
rect 40572 35138 40628 35140
rect 40572 35086 40574 35138
rect 40574 35086 40626 35138
rect 40626 35086 40628 35138
rect 40572 35084 40628 35086
rect 40348 34354 40404 34356
rect 40348 34302 40350 34354
rect 40350 34302 40402 34354
rect 40402 34302 40404 34354
rect 40348 34300 40404 34302
rect 40012 33964 40068 34020
rect 40348 33852 40404 33908
rect 38668 33628 38724 33684
rect 39452 33516 39508 33572
rect 38780 32786 38836 32788
rect 38780 32734 38782 32786
rect 38782 32734 38834 32786
rect 38834 32734 38836 32786
rect 38780 32732 38836 32734
rect 38556 32674 38612 32676
rect 38556 32622 38558 32674
rect 38558 32622 38610 32674
rect 38610 32622 38612 32674
rect 38556 32620 38612 32622
rect 39452 32562 39508 32564
rect 39452 32510 39454 32562
rect 39454 32510 39506 32562
rect 39506 32510 39508 32562
rect 39452 32508 39508 32510
rect 39228 32450 39284 32452
rect 39228 32398 39230 32450
rect 39230 32398 39282 32450
rect 39282 32398 39284 32450
rect 39228 32396 39284 32398
rect 38556 31778 38612 31780
rect 38556 31726 38558 31778
rect 38558 31726 38610 31778
rect 38610 31726 38612 31778
rect 38556 31724 38612 31726
rect 38332 31500 38388 31556
rect 38780 31164 38836 31220
rect 37660 31052 37716 31108
rect 37324 30604 37380 30660
rect 36876 29260 36932 29316
rect 36428 28252 36484 28308
rect 36988 29036 37044 29092
rect 36652 28924 36708 28980
rect 36988 28642 37044 28644
rect 36988 28590 36990 28642
rect 36990 28590 37042 28642
rect 37042 28590 37044 28642
rect 36988 28588 37044 28590
rect 37212 29932 37268 29988
rect 37212 29426 37268 29428
rect 37212 29374 37214 29426
rect 37214 29374 37266 29426
rect 37266 29374 37268 29426
rect 37212 29372 37268 29374
rect 37212 28812 37268 28868
rect 38108 30940 38164 30996
rect 37772 30828 37828 30884
rect 37436 29932 37492 29988
rect 36316 26796 36372 26852
rect 36764 27804 36820 27860
rect 36316 22370 36372 22372
rect 36316 22318 36318 22370
rect 36318 22318 36370 22370
rect 36370 22318 36372 22370
rect 36316 22316 36372 22318
rect 37100 27692 37156 27748
rect 37212 27580 37268 27636
rect 37212 27020 37268 27076
rect 36988 25506 37044 25508
rect 36988 25454 36990 25506
rect 36990 25454 37042 25506
rect 37042 25454 37044 25506
rect 36988 25452 37044 25454
rect 36540 24332 36596 24388
rect 36652 24668 36708 24724
rect 36988 23714 37044 23716
rect 36988 23662 36990 23714
rect 36990 23662 37042 23714
rect 37042 23662 37044 23714
rect 36988 23660 37044 23662
rect 37324 26796 37380 26852
rect 37996 30156 38052 30212
rect 37996 29596 38052 29652
rect 41020 36428 41076 36484
rect 40908 36370 40964 36372
rect 40908 36318 40910 36370
rect 40910 36318 40962 36370
rect 40962 36318 40964 36370
rect 40908 36316 40964 36318
rect 41020 35980 41076 36036
rect 41468 37436 41524 37492
rect 41356 36764 41412 36820
rect 41132 34636 41188 34692
rect 41244 34412 41300 34468
rect 40908 34188 40964 34244
rect 40796 34130 40852 34132
rect 40796 34078 40798 34130
rect 40798 34078 40850 34130
rect 40850 34078 40852 34130
rect 40796 34076 40852 34078
rect 41132 33852 41188 33908
rect 41020 33516 41076 33572
rect 40348 33180 40404 33236
rect 39788 32786 39844 32788
rect 39788 32734 39790 32786
rect 39790 32734 39842 32786
rect 39842 32734 39844 32786
rect 39788 32732 39844 32734
rect 39676 32620 39732 32676
rect 39676 31836 39732 31892
rect 41132 33068 41188 33124
rect 40012 31164 40068 31220
rect 40124 32562 40180 32564
rect 40124 32510 40126 32562
rect 40126 32510 40178 32562
rect 40178 32510 40180 32562
rect 40124 32508 40180 32510
rect 40684 31778 40740 31780
rect 40684 31726 40686 31778
rect 40686 31726 40738 31778
rect 40738 31726 40740 31778
rect 40684 31724 40740 31726
rect 40124 31052 40180 31108
rect 40908 30882 40964 30884
rect 40908 30830 40910 30882
rect 40910 30830 40962 30882
rect 40962 30830 40964 30882
rect 40908 30828 40964 30830
rect 41692 37100 41748 37156
rect 41692 36876 41748 36932
rect 41468 35586 41524 35588
rect 41468 35534 41470 35586
rect 41470 35534 41522 35586
rect 41522 35534 41524 35586
rect 41468 35532 41524 35534
rect 41580 34860 41636 34916
rect 41356 33964 41412 34020
rect 41580 33852 41636 33908
rect 42140 37996 42196 38052
rect 42028 36482 42084 36484
rect 42028 36430 42030 36482
rect 42030 36430 42082 36482
rect 42082 36430 42084 36482
rect 42028 36428 42084 36430
rect 42924 43538 42980 43540
rect 42924 43486 42926 43538
rect 42926 43486 42978 43538
rect 42978 43486 42980 43538
rect 42924 43484 42980 43486
rect 42924 42140 42980 42196
rect 42700 41970 42756 41972
rect 42700 41918 42702 41970
rect 42702 41918 42754 41970
rect 42754 41918 42756 41970
rect 42700 41916 42756 41918
rect 42476 40796 42532 40852
rect 43148 44994 43204 44996
rect 43148 44942 43150 44994
rect 43150 44942 43202 44994
rect 43202 44942 43204 44994
rect 43148 44940 43204 44942
rect 43820 47628 43876 47684
rect 44604 51996 44660 52052
rect 44268 50316 44324 50372
rect 44380 50428 44436 50484
rect 44044 49138 44100 49140
rect 44044 49086 44046 49138
rect 44046 49086 44098 49138
rect 44098 49086 44100 49138
rect 44044 49084 44100 49086
rect 44492 50876 44548 50932
rect 45052 53618 45108 53620
rect 45052 53566 45054 53618
rect 45054 53566 45106 53618
rect 45106 53566 45108 53618
rect 45052 53564 45108 53566
rect 45724 54514 45780 54516
rect 45724 54462 45726 54514
rect 45726 54462 45778 54514
rect 45778 54462 45780 54514
rect 45724 54460 45780 54462
rect 45612 54348 45668 54404
rect 45388 53842 45444 53844
rect 45388 53790 45390 53842
rect 45390 53790 45442 53842
rect 45442 53790 45444 53842
rect 45388 53788 45444 53790
rect 46620 57372 46676 57428
rect 46508 56754 46564 56756
rect 46508 56702 46510 56754
rect 46510 56702 46562 56754
rect 46562 56702 46564 56754
rect 46508 56700 46564 56702
rect 47068 57260 47124 57316
rect 47628 57484 47684 57540
rect 46620 55580 46676 55636
rect 46844 55916 46900 55972
rect 46508 55186 46564 55188
rect 46508 55134 46510 55186
rect 46510 55134 46562 55186
rect 46562 55134 46564 55186
rect 46508 55132 46564 55134
rect 46396 54908 46452 54964
rect 46284 54796 46340 54852
rect 46620 54514 46676 54516
rect 46620 54462 46622 54514
rect 46622 54462 46674 54514
rect 46674 54462 46676 54514
rect 46620 54460 46676 54462
rect 47180 55074 47236 55076
rect 47180 55022 47182 55074
rect 47182 55022 47234 55074
rect 47234 55022 47236 55074
rect 47180 55020 47236 55022
rect 47404 55074 47460 55076
rect 47404 55022 47406 55074
rect 47406 55022 47458 55074
rect 47458 55022 47460 55074
rect 47404 55020 47460 55022
rect 48972 60226 49028 60228
rect 48972 60174 48974 60226
rect 48974 60174 49026 60226
rect 49026 60174 49028 60226
rect 48972 60172 49028 60174
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 48412 59388 48468 59444
rect 49756 59442 49812 59444
rect 49756 59390 49758 59442
rect 49758 59390 49810 59442
rect 49810 59390 49812 59442
rect 49756 59388 49812 59390
rect 48076 58492 48132 58548
rect 52108 58546 52164 58548
rect 52108 58494 52110 58546
rect 52110 58494 52162 58546
rect 52162 58494 52164 58546
rect 52108 58492 52164 58494
rect 51324 58434 51380 58436
rect 51324 58382 51326 58434
rect 51326 58382 51378 58434
rect 51378 58382 51380 58434
rect 51324 58380 51380 58382
rect 50764 58322 50820 58324
rect 50764 58270 50766 58322
rect 50766 58270 50818 58322
rect 50818 58270 50820 58322
rect 50764 58268 50820 58270
rect 51548 58268 51604 58324
rect 48524 58210 48580 58212
rect 48524 58158 48526 58210
rect 48526 58158 48578 58210
rect 48578 58158 48580 58210
rect 48524 58156 48580 58158
rect 48972 58044 49028 58100
rect 49196 58156 49252 58212
rect 48412 57932 48468 57988
rect 48076 57708 48132 57764
rect 47964 57650 48020 57652
rect 47964 57598 47966 57650
rect 47966 57598 48018 57650
rect 48018 57598 48020 57650
rect 47964 57596 48020 57598
rect 47628 56754 47684 56756
rect 47628 56702 47630 56754
rect 47630 56702 47682 56754
rect 47682 56702 47684 56754
rect 47628 56700 47684 56702
rect 48076 56140 48132 56196
rect 48188 56082 48244 56084
rect 48188 56030 48190 56082
rect 48190 56030 48242 56082
rect 48242 56030 48244 56082
rect 48188 56028 48244 56030
rect 47628 55692 47684 55748
rect 47740 55410 47796 55412
rect 47740 55358 47742 55410
rect 47742 55358 47794 55410
rect 47794 55358 47796 55410
rect 47740 55356 47796 55358
rect 47964 55298 48020 55300
rect 47964 55246 47966 55298
rect 47966 55246 48018 55298
rect 48018 55246 48020 55298
rect 47964 55244 48020 55246
rect 46284 54348 46340 54404
rect 46620 54124 46676 54180
rect 45836 53676 45892 53732
rect 46508 53676 46564 53732
rect 45724 53564 45780 53620
rect 45052 52556 45108 52612
rect 45388 52780 45444 52836
rect 46060 53452 46116 53508
rect 45836 53004 45892 53060
rect 46508 53340 46564 53396
rect 46396 53170 46452 53172
rect 46396 53118 46398 53170
rect 46398 53118 46450 53170
rect 46450 53118 46452 53170
rect 46396 53116 46452 53118
rect 46508 52892 46564 52948
rect 45164 52162 45220 52164
rect 45164 52110 45166 52162
rect 45166 52110 45218 52162
rect 45218 52110 45220 52162
rect 45164 52108 45220 52110
rect 45052 50316 45108 50372
rect 45052 48860 45108 48916
rect 44604 48242 44660 48244
rect 44604 48190 44606 48242
rect 44606 48190 44658 48242
rect 44658 48190 44660 48242
rect 44604 48188 44660 48190
rect 44156 47404 44212 47460
rect 44828 47516 44884 47572
rect 44268 47234 44324 47236
rect 44268 47182 44270 47234
rect 44270 47182 44322 47234
rect 44322 47182 44324 47234
rect 44268 47180 44324 47182
rect 44044 46898 44100 46900
rect 44044 46846 44046 46898
rect 44046 46846 44098 46898
rect 44098 46846 44100 46898
rect 44044 46844 44100 46846
rect 43820 45724 43876 45780
rect 44268 45612 44324 45668
rect 44380 45500 44436 45556
rect 43932 45388 43988 45444
rect 44828 46674 44884 46676
rect 44828 46622 44830 46674
rect 44830 46622 44882 46674
rect 44882 46622 44884 46674
rect 44828 46620 44884 46622
rect 45164 48300 45220 48356
rect 44940 46508 44996 46564
rect 44940 46284 44996 46340
rect 45164 46060 45220 46116
rect 44940 46002 44996 46004
rect 44940 45950 44942 46002
rect 44942 45950 44994 46002
rect 44994 45950 44996 46002
rect 44940 45948 44996 45950
rect 45948 52332 46004 52388
rect 45836 52108 45892 52164
rect 45724 50428 45780 50484
rect 45500 49980 45556 50036
rect 45500 49084 45556 49140
rect 45836 49308 45892 49364
rect 46060 49532 46116 49588
rect 45948 48972 46004 49028
rect 45388 48188 45444 48244
rect 45500 48076 45556 48132
rect 45612 47628 45668 47684
rect 45724 47404 45780 47460
rect 45388 45778 45444 45780
rect 45388 45726 45390 45778
rect 45390 45726 45442 45778
rect 45442 45726 45444 45778
rect 45388 45724 45444 45726
rect 44828 45612 44884 45668
rect 43820 45218 43876 45220
rect 43820 45166 43822 45218
rect 43822 45166 43874 45218
rect 43874 45166 43876 45218
rect 43820 45164 43876 45166
rect 43708 44492 43764 44548
rect 43148 44322 43204 44324
rect 43148 44270 43150 44322
rect 43150 44270 43202 44322
rect 43202 44270 43204 44322
rect 43148 44268 43204 44270
rect 43932 44546 43988 44548
rect 43932 44494 43934 44546
rect 43934 44494 43986 44546
rect 43986 44494 43988 44546
rect 43932 44492 43988 44494
rect 43484 43596 43540 43652
rect 43820 43650 43876 43652
rect 43820 43598 43822 43650
rect 43822 43598 43874 43650
rect 43874 43598 43876 43650
rect 43820 43596 43876 43598
rect 43596 43484 43652 43540
rect 44492 45106 44548 45108
rect 44492 45054 44494 45106
rect 44494 45054 44546 45106
rect 44546 45054 44548 45106
rect 44492 45052 44548 45054
rect 44156 43538 44212 43540
rect 44156 43486 44158 43538
rect 44158 43486 44210 43538
rect 44210 43486 44212 43538
rect 44156 43484 44212 43486
rect 44268 43708 44324 43764
rect 44380 44156 44436 44212
rect 44716 44940 44772 44996
rect 45164 45164 45220 45220
rect 44940 44322 44996 44324
rect 44940 44270 44942 44322
rect 44942 44270 44994 44322
rect 44994 44270 44996 44322
rect 44940 44268 44996 44270
rect 44828 43820 44884 43876
rect 45388 44210 45444 44212
rect 45388 44158 45390 44210
rect 45390 44158 45442 44210
rect 45442 44158 45444 44210
rect 45388 44156 45444 44158
rect 43708 42140 43764 42196
rect 43260 41970 43316 41972
rect 43260 41918 43262 41970
rect 43262 41918 43314 41970
rect 43314 41918 43316 41970
rect 43260 41916 43316 41918
rect 44380 42588 44436 42644
rect 45052 42476 45108 42532
rect 44380 42194 44436 42196
rect 44380 42142 44382 42194
rect 44382 42142 44434 42194
rect 44434 42142 44436 42194
rect 44380 42140 44436 42142
rect 44940 42028 44996 42084
rect 42700 39506 42756 39508
rect 42700 39454 42702 39506
rect 42702 39454 42754 39506
rect 42754 39454 42756 39506
rect 42700 39452 42756 39454
rect 43036 40626 43092 40628
rect 43036 40574 43038 40626
rect 43038 40574 43090 40626
rect 43090 40574 43092 40626
rect 43036 40572 43092 40574
rect 42924 40236 42980 40292
rect 43932 39730 43988 39732
rect 43932 39678 43934 39730
rect 43934 39678 43986 39730
rect 43986 39678 43988 39730
rect 43932 39676 43988 39678
rect 42812 39228 42868 39284
rect 43036 39116 43092 39172
rect 42364 36540 42420 36596
rect 42364 35698 42420 35700
rect 42364 35646 42366 35698
rect 42366 35646 42418 35698
rect 42418 35646 42420 35698
rect 42364 35644 42420 35646
rect 42028 35308 42084 35364
rect 42476 35532 42532 35588
rect 41692 32396 41748 32452
rect 41916 35084 41972 35140
rect 41692 32060 41748 32116
rect 41244 30716 41300 30772
rect 41468 31500 41524 31556
rect 40012 30268 40068 30324
rect 38556 30044 38612 30100
rect 37772 28082 37828 28084
rect 37772 28030 37774 28082
rect 37774 28030 37826 28082
rect 37826 28030 37828 28082
rect 37772 28028 37828 28030
rect 37548 27858 37604 27860
rect 37548 27806 37550 27858
rect 37550 27806 37602 27858
rect 37602 27806 37604 27858
rect 37548 27804 37604 27806
rect 37772 27244 37828 27300
rect 37660 27074 37716 27076
rect 37660 27022 37662 27074
rect 37662 27022 37714 27074
rect 37714 27022 37716 27074
rect 37660 27020 37716 27022
rect 38892 29986 38948 29988
rect 38892 29934 38894 29986
rect 38894 29934 38946 29986
rect 38946 29934 38948 29986
rect 38892 29932 38948 29934
rect 39228 29932 39284 29988
rect 38780 29202 38836 29204
rect 38780 29150 38782 29202
rect 38782 29150 38834 29202
rect 38834 29150 38836 29202
rect 38780 29148 38836 29150
rect 39004 28812 39060 28868
rect 38556 28588 38612 28644
rect 39788 29986 39844 29988
rect 39788 29934 39790 29986
rect 39790 29934 39842 29986
rect 39842 29934 39844 29986
rect 39788 29932 39844 29934
rect 39340 29596 39396 29652
rect 39116 28418 39172 28420
rect 39116 28366 39118 28418
rect 39118 28366 39170 28418
rect 39170 28366 39172 28418
rect 39116 28364 39172 28366
rect 38444 28252 38500 28308
rect 38556 28140 38612 28196
rect 39900 28812 39956 28868
rect 39676 28588 39732 28644
rect 38332 27804 38388 27860
rect 38668 27804 38724 27860
rect 38332 27244 38388 27300
rect 38444 27692 38500 27748
rect 39228 28028 39284 28084
rect 39788 28364 39844 28420
rect 39788 27692 39844 27748
rect 41356 30156 41412 30212
rect 40460 29986 40516 29988
rect 40460 29934 40462 29986
rect 40462 29934 40514 29986
rect 40514 29934 40516 29986
rect 40460 29932 40516 29934
rect 40124 29596 40180 29652
rect 40348 29426 40404 29428
rect 40348 29374 40350 29426
rect 40350 29374 40402 29426
rect 40402 29374 40404 29426
rect 40348 29372 40404 29374
rect 40236 29314 40292 29316
rect 40236 29262 40238 29314
rect 40238 29262 40290 29314
rect 40290 29262 40292 29314
rect 40236 29260 40292 29262
rect 40124 29036 40180 29092
rect 39900 28252 39956 28308
rect 39116 27132 39172 27188
rect 38220 26796 38276 26852
rect 37772 25900 37828 25956
rect 37324 24108 37380 24164
rect 37324 23884 37380 23940
rect 36988 23436 37044 23492
rect 36652 23324 36708 23380
rect 36988 23266 37044 23268
rect 36988 23214 36990 23266
rect 36990 23214 37042 23266
rect 37042 23214 37044 23266
rect 36988 23212 37044 23214
rect 36652 23154 36708 23156
rect 36652 23102 36654 23154
rect 36654 23102 36706 23154
rect 36706 23102 36708 23154
rect 36652 23100 36708 23102
rect 36428 22146 36484 22148
rect 36428 22094 36430 22146
rect 36430 22094 36482 22146
rect 36482 22094 36484 22146
rect 36428 22092 36484 22094
rect 35980 20076 36036 20132
rect 36092 20018 36148 20020
rect 36092 19966 36094 20018
rect 36094 19966 36146 20018
rect 36146 19966 36148 20018
rect 36092 19964 36148 19966
rect 35756 19234 35812 19236
rect 35756 19182 35758 19234
rect 35758 19182 35810 19234
rect 35810 19182 35812 19234
rect 35756 19180 35812 19182
rect 35980 19852 36036 19908
rect 35868 18172 35924 18228
rect 35868 17724 35924 17780
rect 34636 15820 34692 15876
rect 33964 14700 34020 14756
rect 34636 14924 34692 14980
rect 34524 14754 34580 14756
rect 34524 14702 34526 14754
rect 34526 14702 34578 14754
rect 34578 14702 34580 14754
rect 34524 14700 34580 14702
rect 34524 14364 34580 14420
rect 34412 14252 34468 14308
rect 34076 12850 34132 12852
rect 34076 12798 34078 12850
rect 34078 12798 34130 12850
rect 34130 12798 34132 12850
rect 34076 12796 34132 12798
rect 33180 12012 33236 12068
rect 33292 11900 33348 11956
rect 31276 10386 31332 10388
rect 31276 10334 31278 10386
rect 31278 10334 31330 10386
rect 31330 10334 31332 10386
rect 31276 10332 31332 10334
rect 31276 9996 31332 10052
rect 31388 9938 31444 9940
rect 31388 9886 31390 9938
rect 31390 9886 31442 9938
rect 31442 9886 31444 9938
rect 31388 9884 31444 9886
rect 31276 9324 31332 9380
rect 31612 9266 31668 9268
rect 31612 9214 31614 9266
rect 31614 9214 31666 9266
rect 31666 9214 31668 9266
rect 31612 9212 31668 9214
rect 31164 8764 31220 8820
rect 30492 7474 30548 7476
rect 30492 7422 30494 7474
rect 30494 7422 30546 7474
rect 30546 7422 30548 7474
rect 30492 7420 30548 7422
rect 29820 6748 29876 6804
rect 30268 7308 30324 7364
rect 29596 5628 29652 5684
rect 29596 4284 29652 4340
rect 29484 3500 29540 3556
rect 30268 6860 30324 6916
rect 30492 6860 30548 6916
rect 30044 6300 30100 6356
rect 30828 7980 30884 8036
rect 31388 8204 31444 8260
rect 30940 6748 30996 6804
rect 31276 6466 31332 6468
rect 31276 6414 31278 6466
rect 31278 6414 31330 6466
rect 31330 6414 31332 6466
rect 31276 6412 31332 6414
rect 31500 7980 31556 8036
rect 31612 6914 31668 6916
rect 31612 6862 31614 6914
rect 31614 6862 31666 6914
rect 31666 6862 31668 6914
rect 31612 6860 31668 6862
rect 31724 6300 31780 6356
rect 31388 6188 31444 6244
rect 30156 5964 30212 6020
rect 30380 5516 30436 5572
rect 30156 5068 30212 5124
rect 30716 5068 30772 5124
rect 31052 6018 31108 6020
rect 31052 5966 31054 6018
rect 31054 5966 31106 6018
rect 31106 5966 31108 6018
rect 31052 5964 31108 5966
rect 31612 5964 31668 6020
rect 31724 5852 31780 5908
rect 31500 5516 31556 5572
rect 30828 4956 30884 5012
rect 30044 3554 30100 3556
rect 30044 3502 30046 3554
rect 30046 3502 30098 3554
rect 30098 3502 30100 3554
rect 30044 3500 30100 3502
rect 31052 3836 31108 3892
rect 31500 3612 31556 3668
rect 30268 3500 30324 3556
rect 23212 3164 23268 3220
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 13804 2940 13860 2996
rect 31948 9826 32004 9828
rect 31948 9774 31950 9826
rect 31950 9774 32002 9826
rect 32002 9774 32004 9826
rect 31948 9772 32004 9774
rect 32508 9602 32564 9604
rect 32508 9550 32510 9602
rect 32510 9550 32562 9602
rect 32562 9550 32564 9602
rect 32508 9548 32564 9550
rect 32396 9154 32452 9156
rect 32396 9102 32398 9154
rect 32398 9102 32450 9154
rect 32450 9102 32452 9154
rect 32396 9100 32452 9102
rect 32284 9042 32340 9044
rect 32284 8990 32286 9042
rect 32286 8990 32338 9042
rect 32338 8990 32340 9042
rect 32284 8988 32340 8990
rect 31948 8764 32004 8820
rect 32172 8428 32228 8484
rect 32508 8988 32564 9044
rect 32508 8428 32564 8484
rect 32732 8316 32788 8372
rect 31948 6748 32004 6804
rect 32172 6972 32228 7028
rect 32620 6972 32676 7028
rect 32508 6860 32564 6916
rect 32060 6636 32116 6692
rect 31948 6412 32004 6468
rect 32620 6188 32676 6244
rect 32396 5852 32452 5908
rect 32060 5404 32116 5460
rect 32060 5122 32116 5124
rect 32060 5070 32062 5122
rect 32062 5070 32114 5122
rect 32114 5070 32116 5122
rect 32060 5068 32116 5070
rect 32172 5010 32228 5012
rect 32172 4958 32174 5010
rect 32174 4958 32226 5010
rect 32226 4958 32228 5010
rect 32172 4956 32228 4958
rect 32620 5964 32676 6020
rect 32508 5628 32564 5684
rect 32284 3388 32340 3444
rect 33516 12012 33572 12068
rect 34524 12908 34580 12964
rect 34524 12684 34580 12740
rect 33068 11170 33124 11172
rect 33068 11118 33070 11170
rect 33070 11118 33122 11170
rect 33122 11118 33124 11170
rect 33068 11116 33124 11118
rect 33964 11170 34020 11172
rect 33964 11118 33966 11170
rect 33966 11118 34018 11170
rect 34018 11118 34020 11170
rect 33964 11116 34020 11118
rect 33516 10834 33572 10836
rect 33516 10782 33518 10834
rect 33518 10782 33570 10834
rect 33570 10782 33572 10834
rect 33516 10780 33572 10782
rect 33404 10668 33460 10724
rect 34188 10668 34244 10724
rect 33180 10556 33236 10612
rect 33292 9772 33348 9828
rect 32956 9100 33012 9156
rect 33404 9548 33460 9604
rect 33628 8930 33684 8932
rect 33628 8878 33630 8930
rect 33630 8878 33682 8930
rect 33682 8878 33684 8930
rect 33628 8876 33684 8878
rect 34076 10556 34132 10612
rect 35868 17442 35924 17444
rect 35868 17390 35870 17442
rect 35870 17390 35922 17442
rect 35922 17390 35924 17442
rect 35868 17388 35924 17390
rect 36316 20524 36372 20580
rect 36092 18956 36148 19012
rect 36204 18732 36260 18788
rect 36092 18284 36148 18340
rect 36092 17724 36148 17780
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34972 14924 35028 14980
rect 35084 15708 35140 15764
rect 34748 14418 34804 14420
rect 34748 14366 34750 14418
rect 34750 14366 34802 14418
rect 34802 14366 34804 14418
rect 34748 14364 34804 14366
rect 34972 14418 35028 14420
rect 34972 14366 34974 14418
rect 34974 14366 35026 14418
rect 35026 14366 35028 14418
rect 34972 14364 35028 14366
rect 34748 14140 34804 14196
rect 33964 9826 34020 9828
rect 33964 9774 33966 9826
rect 33966 9774 34018 9826
rect 34018 9774 34020 9826
rect 33964 9772 34020 9774
rect 33852 9154 33908 9156
rect 33852 9102 33854 9154
rect 33854 9102 33906 9154
rect 33906 9102 33908 9154
rect 33852 9100 33908 9102
rect 33964 9042 34020 9044
rect 33964 8990 33966 9042
rect 33966 8990 34018 9042
rect 34018 8990 34020 9042
rect 33964 8988 34020 8990
rect 32956 8146 33012 8148
rect 32956 8094 32958 8146
rect 32958 8094 33010 8146
rect 33010 8094 33012 8146
rect 32956 8092 33012 8094
rect 33628 8034 33684 8036
rect 33628 7982 33630 8034
rect 33630 7982 33682 8034
rect 33682 7982 33684 8034
rect 33628 7980 33684 7982
rect 33516 7474 33572 7476
rect 33516 7422 33518 7474
rect 33518 7422 33570 7474
rect 33570 7422 33572 7474
rect 33516 7420 33572 7422
rect 33180 7362 33236 7364
rect 33180 7310 33182 7362
rect 33182 7310 33234 7362
rect 33234 7310 33236 7362
rect 33180 7308 33236 7310
rect 33292 6914 33348 6916
rect 33292 6862 33294 6914
rect 33294 6862 33346 6914
rect 33346 6862 33348 6914
rect 33292 6860 33348 6862
rect 32956 6636 33012 6692
rect 33628 6412 33684 6468
rect 33516 6188 33572 6244
rect 32844 5628 32900 5684
rect 33292 5906 33348 5908
rect 33292 5854 33294 5906
rect 33294 5854 33346 5906
rect 33346 5854 33348 5906
rect 33292 5852 33348 5854
rect 33516 5852 33572 5908
rect 33068 5740 33124 5796
rect 33628 5740 33684 5796
rect 33404 5292 33460 5348
rect 33516 4956 33572 5012
rect 32956 3724 33012 3780
rect 33404 4338 33460 4340
rect 33404 4286 33406 4338
rect 33406 4286 33458 4338
rect 33458 4286 33460 4338
rect 33404 4284 33460 4286
rect 33852 7532 33908 7588
rect 33852 7084 33908 7140
rect 33964 6860 34020 6916
rect 34524 9826 34580 9828
rect 34524 9774 34526 9826
rect 34526 9774 34578 9826
rect 34578 9774 34580 9826
rect 34524 9772 34580 9774
rect 34860 13468 34916 13524
rect 35868 15036 35924 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35532 14754 35588 14756
rect 35532 14702 35534 14754
rect 35534 14702 35586 14754
rect 35586 14702 35588 14754
rect 35532 14700 35588 14702
rect 35868 14476 35924 14532
rect 36092 14418 36148 14420
rect 36092 14366 36094 14418
rect 36094 14366 36146 14418
rect 36146 14366 36148 14418
rect 36092 14364 36148 14366
rect 35868 14140 35924 14196
rect 35420 13858 35476 13860
rect 35420 13806 35422 13858
rect 35422 13806 35474 13858
rect 35474 13806 35476 13858
rect 35420 13804 35476 13806
rect 35196 13746 35252 13748
rect 35196 13694 35198 13746
rect 35198 13694 35250 13746
rect 35250 13694 35252 13746
rect 35196 13692 35252 13694
rect 35644 13522 35700 13524
rect 35644 13470 35646 13522
rect 35646 13470 35698 13522
rect 35698 13470 35700 13522
rect 35644 13468 35700 13470
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 12962 35252 12964
rect 35196 12910 35198 12962
rect 35198 12910 35250 12962
rect 35250 12910 35252 12962
rect 35196 12908 35252 12910
rect 35532 12796 35588 12852
rect 35308 12348 35364 12404
rect 36316 17388 36372 17444
rect 36540 19292 36596 19348
rect 37436 23436 37492 23492
rect 38108 25900 38164 25956
rect 38108 25676 38164 25732
rect 39004 26236 39060 26292
rect 38220 25564 38276 25620
rect 38892 25228 38948 25284
rect 37996 23100 38052 23156
rect 38108 24108 38164 24164
rect 37996 22930 38052 22932
rect 37996 22878 37998 22930
rect 37998 22878 38050 22930
rect 38050 22878 38052 22930
rect 37996 22876 38052 22878
rect 37548 22316 37604 22372
rect 37436 20636 37492 20692
rect 37212 19964 37268 20020
rect 37324 19852 37380 19908
rect 37100 19010 37156 19012
rect 37100 18958 37102 19010
rect 37102 18958 37154 19010
rect 37154 18958 37156 19010
rect 37100 18956 37156 18958
rect 36428 18396 36484 18452
rect 36652 17948 36708 18004
rect 36428 16044 36484 16100
rect 36540 14364 36596 14420
rect 35980 13746 36036 13748
rect 35980 13694 35982 13746
rect 35982 13694 36034 13746
rect 36034 13694 36036 13746
rect 35980 13692 36036 13694
rect 35868 12402 35924 12404
rect 35868 12350 35870 12402
rect 35870 12350 35922 12402
rect 35922 12350 35924 12402
rect 35868 12348 35924 12350
rect 35756 11900 35812 11956
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34972 10892 35028 10948
rect 35084 11452 35140 11508
rect 35868 11506 35924 11508
rect 35868 11454 35870 11506
rect 35870 11454 35922 11506
rect 35922 11454 35924 11506
rect 35868 11452 35924 11454
rect 34860 10780 34916 10836
rect 34972 10610 35028 10612
rect 34972 10558 34974 10610
rect 34974 10558 35026 10610
rect 35026 10558 35028 10610
rect 34972 10556 35028 10558
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34412 8316 34468 8372
rect 34972 9100 35028 9156
rect 34748 8988 34804 9044
rect 34860 8876 34916 8932
rect 34636 8146 34692 8148
rect 34636 8094 34638 8146
rect 34638 8094 34690 8146
rect 34690 8094 34692 8146
rect 34636 8092 34692 8094
rect 34300 6300 34356 6356
rect 34076 6018 34132 6020
rect 34076 5966 34078 6018
rect 34078 5966 34130 6018
rect 34130 5966 34132 6018
rect 34076 5964 34132 5966
rect 33964 5292 34020 5348
rect 34300 5906 34356 5908
rect 34300 5854 34302 5906
rect 34302 5854 34354 5906
rect 34354 5854 34356 5906
rect 34300 5852 34356 5854
rect 34300 5068 34356 5124
rect 33964 3724 34020 3780
rect 34524 6578 34580 6580
rect 34524 6526 34526 6578
rect 34526 6526 34578 6578
rect 34578 6526 34580 6578
rect 34524 6524 34580 6526
rect 34748 7308 34804 7364
rect 36092 9772 36148 9828
rect 35980 9714 36036 9716
rect 35980 9662 35982 9714
rect 35982 9662 36034 9714
rect 36034 9662 36036 9714
rect 35980 9660 36036 9662
rect 35532 9602 35588 9604
rect 35532 9550 35534 9602
rect 35534 9550 35586 9602
rect 35586 9550 35588 9602
rect 35532 9548 35588 9550
rect 35420 8764 35476 8820
rect 35644 9154 35700 9156
rect 35644 9102 35646 9154
rect 35646 9102 35698 9154
rect 35698 9102 35700 9154
rect 35644 9100 35700 9102
rect 35532 8988 35588 9044
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35420 8428 35476 8484
rect 35756 8988 35812 9044
rect 36092 8988 36148 9044
rect 35980 8258 36036 8260
rect 35980 8206 35982 8258
rect 35982 8206 36034 8258
rect 36034 8206 36036 8258
rect 35980 8204 36036 8206
rect 35868 7980 35924 8036
rect 36092 8092 36148 8148
rect 35420 7532 35476 7588
rect 35756 7532 35812 7588
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 6636 35252 6692
rect 35308 6578 35364 6580
rect 35308 6526 35310 6578
rect 35310 6526 35362 6578
rect 35362 6526 35364 6578
rect 35308 6524 35364 6526
rect 34972 6466 35028 6468
rect 34972 6414 34974 6466
rect 34974 6414 35026 6466
rect 35026 6414 35028 6466
rect 34972 6412 35028 6414
rect 35644 7308 35700 7364
rect 35196 6018 35252 6020
rect 35196 5966 35198 6018
rect 35198 5966 35250 6018
rect 35250 5966 35252 6018
rect 35196 5964 35252 5966
rect 35756 6412 35812 6468
rect 35980 6300 36036 6356
rect 36092 7420 36148 7476
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35980 5346 36036 5348
rect 35980 5294 35982 5346
rect 35982 5294 36034 5346
rect 36034 5294 36036 5346
rect 35980 5292 36036 5294
rect 34972 5122 35028 5124
rect 34972 5070 34974 5122
rect 34974 5070 35026 5122
rect 35026 5070 35028 5122
rect 34972 5068 35028 5070
rect 34860 5010 34916 5012
rect 34860 4958 34862 5010
rect 34862 4958 34914 5010
rect 34914 4958 34916 5010
rect 34860 4956 34916 4958
rect 35980 4844 36036 4900
rect 34972 4620 35028 4676
rect 36092 4508 36148 4564
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 37996 21084 38052 21140
rect 38668 24722 38724 24724
rect 38668 24670 38670 24722
rect 38670 24670 38722 24722
rect 38722 24670 38724 24722
rect 38668 24668 38724 24670
rect 38220 23324 38276 23380
rect 38668 23548 38724 23604
rect 38332 22988 38388 23044
rect 39452 27356 39508 27412
rect 40012 28028 40068 28084
rect 40124 27916 40180 27972
rect 42028 34748 42084 34804
rect 42028 34300 42084 34356
rect 42924 38556 42980 38612
rect 42812 38444 42868 38500
rect 42700 38274 42756 38276
rect 42700 38222 42702 38274
rect 42702 38222 42754 38274
rect 42754 38222 42756 38274
rect 42700 38220 42756 38222
rect 42700 38050 42756 38052
rect 42700 37998 42702 38050
rect 42702 37998 42754 38050
rect 42754 37998 42756 38050
rect 42700 37996 42756 37998
rect 42700 36540 42756 36596
rect 43484 38780 43540 38836
rect 42924 36204 42980 36260
rect 42812 36092 42868 36148
rect 42924 35420 42980 35476
rect 42700 34860 42756 34916
rect 42812 35308 42868 35364
rect 42476 34748 42532 34804
rect 42812 34636 42868 34692
rect 42140 34130 42196 34132
rect 42140 34078 42142 34130
rect 42142 34078 42194 34130
rect 42194 34078 42196 34130
rect 42140 34076 42196 34078
rect 42028 32508 42084 32564
rect 42140 33852 42196 33908
rect 42588 34242 42644 34244
rect 42588 34190 42590 34242
rect 42590 34190 42642 34242
rect 42642 34190 42644 34242
rect 42588 34188 42644 34190
rect 43148 37826 43204 37828
rect 43148 37774 43150 37826
rect 43150 37774 43202 37826
rect 43202 37774 43204 37826
rect 43148 37772 43204 37774
rect 43596 38444 43652 38500
rect 43596 38220 43652 38276
rect 43708 37884 43764 37940
rect 43820 37772 43876 37828
rect 43708 36988 43764 37044
rect 43596 36428 43652 36484
rect 43148 35644 43204 35700
rect 43148 33180 43204 33236
rect 43484 35868 43540 35924
rect 43932 35868 43988 35924
rect 42252 31948 42308 32004
rect 42140 31612 42196 31668
rect 42252 31724 42308 31780
rect 41916 31388 41972 31444
rect 41356 29596 41412 29652
rect 41244 29372 41300 29428
rect 40796 28812 40852 28868
rect 40460 28140 40516 28196
rect 39676 26348 39732 26404
rect 39452 26290 39508 26292
rect 39452 26238 39454 26290
rect 39454 26238 39506 26290
rect 39506 26238 39508 26290
rect 39452 26236 39508 26238
rect 40348 27356 40404 27412
rect 41244 28700 41300 28756
rect 41356 28588 41412 28644
rect 41244 28364 41300 28420
rect 40908 27244 40964 27300
rect 40460 26572 40516 26628
rect 40012 26348 40068 26404
rect 40124 26236 40180 26292
rect 39116 25340 39172 25396
rect 39676 24220 39732 24276
rect 39004 23436 39060 23492
rect 39116 22764 39172 22820
rect 39564 23154 39620 23156
rect 39564 23102 39566 23154
rect 39566 23102 39618 23154
rect 39618 23102 39620 23154
rect 39564 23100 39620 23102
rect 39340 22876 39396 22932
rect 39564 22316 39620 22372
rect 39340 22092 39396 22148
rect 37772 20076 37828 20132
rect 37660 20018 37716 20020
rect 37660 19966 37662 20018
rect 37662 19966 37714 20018
rect 37714 19966 37716 20018
rect 37660 19964 37716 19966
rect 36988 18060 37044 18116
rect 36988 17388 37044 17444
rect 37548 16380 37604 16436
rect 37548 16098 37604 16100
rect 37548 16046 37550 16098
rect 37550 16046 37602 16098
rect 37602 16046 37604 16098
rect 37548 16044 37604 16046
rect 36988 15874 37044 15876
rect 36988 15822 36990 15874
rect 36990 15822 37042 15874
rect 37042 15822 37044 15874
rect 36988 15820 37044 15822
rect 37996 17836 38052 17892
rect 38108 18956 38164 19012
rect 37884 17778 37940 17780
rect 37884 17726 37886 17778
rect 37886 17726 37938 17778
rect 37938 17726 37940 17778
rect 37884 17724 37940 17726
rect 38332 18620 38388 18676
rect 38220 18338 38276 18340
rect 38220 18286 38222 18338
rect 38222 18286 38274 18338
rect 38274 18286 38276 18338
rect 38220 18284 38276 18286
rect 37884 16882 37940 16884
rect 37884 16830 37886 16882
rect 37886 16830 37938 16882
rect 37938 16830 37940 16882
rect 37884 16828 37940 16830
rect 38556 20188 38612 20244
rect 39116 21644 39172 21700
rect 39004 20412 39060 20468
rect 39116 19852 39172 19908
rect 38444 17724 38500 17780
rect 38444 16828 38500 16884
rect 39116 19180 39172 19236
rect 38332 16380 38388 16436
rect 37772 15986 37828 15988
rect 37772 15934 37774 15986
rect 37774 15934 37826 15986
rect 37826 15934 37828 15986
rect 37772 15932 37828 15934
rect 37660 15538 37716 15540
rect 37660 15486 37662 15538
rect 37662 15486 37714 15538
rect 37714 15486 37716 15538
rect 37660 15484 37716 15486
rect 37548 15260 37604 15316
rect 37100 15036 37156 15092
rect 37100 14700 37156 14756
rect 36764 14140 36820 14196
rect 37548 14530 37604 14532
rect 37548 14478 37550 14530
rect 37550 14478 37602 14530
rect 37602 14478 37604 14530
rect 37548 14476 37604 14478
rect 36876 13746 36932 13748
rect 36876 13694 36878 13746
rect 36878 13694 36930 13746
rect 36930 13694 36932 13746
rect 36876 13692 36932 13694
rect 36652 13356 36708 13412
rect 36316 12012 36372 12068
rect 36764 10834 36820 10836
rect 36764 10782 36766 10834
rect 36766 10782 36818 10834
rect 36818 10782 36820 10834
rect 36764 10780 36820 10782
rect 36988 12236 37044 12292
rect 38108 15484 38164 15540
rect 37996 14306 38052 14308
rect 37996 14254 37998 14306
rect 37998 14254 38050 14306
rect 38050 14254 38052 14306
rect 37996 14252 38052 14254
rect 37884 13020 37940 13076
rect 38220 14476 38276 14532
rect 37436 12460 37492 12516
rect 37212 11506 37268 11508
rect 37212 11454 37214 11506
rect 37214 11454 37266 11506
rect 37266 11454 37268 11506
rect 37212 11452 37268 11454
rect 37996 12348 38052 12404
rect 38108 12460 38164 12516
rect 37660 11788 37716 11844
rect 36876 10108 36932 10164
rect 36540 9772 36596 9828
rect 38108 11788 38164 11844
rect 38556 16098 38612 16100
rect 38556 16046 38558 16098
rect 38558 16046 38610 16098
rect 38610 16046 38612 16098
rect 38556 16044 38612 16046
rect 38892 17164 38948 17220
rect 39452 21644 39508 21700
rect 40124 25452 40180 25508
rect 40684 25564 40740 25620
rect 41132 27132 41188 27188
rect 40348 24108 40404 24164
rect 40012 23884 40068 23940
rect 39788 23436 39844 23492
rect 39900 23660 39956 23716
rect 40236 23660 40292 23716
rect 40124 23378 40180 23380
rect 40124 23326 40126 23378
rect 40126 23326 40178 23378
rect 40178 23326 40180 23378
rect 40124 23324 40180 23326
rect 40012 22876 40068 22932
rect 38892 16716 38948 16772
rect 39228 16716 39284 16772
rect 38780 15932 38836 15988
rect 39452 18620 39508 18676
rect 39564 18284 39620 18340
rect 39452 17554 39508 17556
rect 39452 17502 39454 17554
rect 39454 17502 39506 17554
rect 39506 17502 39508 17554
rect 39452 17500 39508 17502
rect 40012 22092 40068 22148
rect 40124 21756 40180 21812
rect 39900 21084 39956 21140
rect 39900 19404 39956 19460
rect 40348 20300 40404 20356
rect 40124 20188 40180 20244
rect 40348 19516 40404 19572
rect 40236 19292 40292 19348
rect 40012 18284 40068 18340
rect 39900 17500 39956 17556
rect 39900 16882 39956 16884
rect 39900 16830 39902 16882
rect 39902 16830 39954 16882
rect 39954 16830 39956 16882
rect 39900 16828 39956 16830
rect 39676 16716 39732 16772
rect 39452 16604 39508 16660
rect 38444 13020 38500 13076
rect 38444 12236 38500 12292
rect 38220 10780 38276 10836
rect 37212 9826 37268 9828
rect 37212 9774 37214 9826
rect 37214 9774 37266 9826
rect 37266 9774 37268 9826
rect 37212 9772 37268 9774
rect 36988 9100 37044 9156
rect 37100 8428 37156 8484
rect 37548 9100 37604 9156
rect 37548 8764 37604 8820
rect 37772 9042 37828 9044
rect 37772 8990 37774 9042
rect 37774 8990 37826 9042
rect 37826 8990 37828 9042
rect 37772 8988 37828 8990
rect 37212 8370 37268 8372
rect 37212 8318 37214 8370
rect 37214 8318 37266 8370
rect 37266 8318 37268 8370
rect 37212 8316 37268 8318
rect 36316 7474 36372 7476
rect 36316 7422 36318 7474
rect 36318 7422 36370 7474
rect 36370 7422 36372 7474
rect 36316 7420 36372 7422
rect 36316 6300 36372 6356
rect 36316 5852 36372 5908
rect 36988 6524 37044 6580
rect 37324 5964 37380 6020
rect 36988 4844 37044 4900
rect 36876 4562 36932 4564
rect 36876 4510 36878 4562
rect 36878 4510 36930 4562
rect 36930 4510 36932 4562
rect 36876 4508 36932 4510
rect 37436 7196 37492 7252
rect 37436 4396 37492 4452
rect 37996 8204 38052 8260
rect 37884 6748 37940 6804
rect 38108 5964 38164 6020
rect 38220 7420 38276 7476
rect 38668 13074 38724 13076
rect 38668 13022 38670 13074
rect 38670 13022 38722 13074
rect 38722 13022 38724 13074
rect 38668 13020 38724 13022
rect 38892 14364 38948 14420
rect 39004 15260 39060 15316
rect 38892 14140 38948 14196
rect 39116 14924 39172 14980
rect 39228 16044 39284 16100
rect 40572 22764 40628 22820
rect 40684 22370 40740 22372
rect 40684 22318 40686 22370
rect 40686 22318 40738 22370
rect 40738 22318 40740 22370
rect 40684 22316 40740 22318
rect 41020 25228 41076 25284
rect 41020 24946 41076 24948
rect 41020 24894 41022 24946
rect 41022 24894 41074 24946
rect 41074 24894 41076 24946
rect 41020 24892 41076 24894
rect 41132 23324 41188 23380
rect 41020 22930 41076 22932
rect 41020 22878 41022 22930
rect 41022 22878 41074 22930
rect 41074 22878 41076 22930
rect 41020 22876 41076 22878
rect 41020 22316 41076 22372
rect 41020 21756 41076 21812
rect 41580 28028 41636 28084
rect 41468 27916 41524 27972
rect 41692 27746 41748 27748
rect 41692 27694 41694 27746
rect 41694 27694 41746 27746
rect 41746 27694 41748 27746
rect 41692 27692 41748 27694
rect 41580 27580 41636 27636
rect 41692 27356 41748 27412
rect 41692 26178 41748 26180
rect 41692 26126 41694 26178
rect 41694 26126 41746 26178
rect 41746 26126 41748 26178
rect 41692 26124 41748 26126
rect 41356 25564 41412 25620
rect 41692 25506 41748 25508
rect 41692 25454 41694 25506
rect 41694 25454 41746 25506
rect 41746 25454 41748 25506
rect 41692 25452 41748 25454
rect 41580 23938 41636 23940
rect 41580 23886 41582 23938
rect 41582 23886 41634 23938
rect 41634 23886 41636 23938
rect 41580 23884 41636 23886
rect 41916 30098 41972 30100
rect 41916 30046 41918 30098
rect 41918 30046 41970 30098
rect 41970 30046 41972 30098
rect 41916 30044 41972 30046
rect 43148 32396 43204 32452
rect 43148 32060 43204 32116
rect 42252 30156 42308 30212
rect 42028 29202 42084 29204
rect 42028 29150 42030 29202
rect 42030 29150 42082 29202
rect 42082 29150 42084 29202
rect 42028 29148 42084 29150
rect 41916 28252 41972 28308
rect 42028 28476 42084 28532
rect 43260 30828 43316 30884
rect 43036 30380 43092 30436
rect 43596 34636 43652 34692
rect 43484 34524 43540 34580
rect 43484 34076 43540 34132
rect 43708 33964 43764 34020
rect 44268 40626 44324 40628
rect 44268 40574 44270 40626
rect 44270 40574 44322 40626
rect 44322 40574 44324 40626
rect 44268 40572 44324 40574
rect 45164 40572 45220 40628
rect 46396 50876 46452 50932
rect 46956 53788 47012 53844
rect 47516 53676 47572 53732
rect 46844 53564 46900 53620
rect 47516 53452 47572 53508
rect 46732 53058 46788 53060
rect 46732 53006 46734 53058
rect 46734 53006 46786 53058
rect 46786 53006 46788 53058
rect 46732 53004 46788 53006
rect 48860 57596 48916 57652
rect 48972 56028 49028 56084
rect 48636 55692 48692 55748
rect 47740 53676 47796 53732
rect 47740 53228 47796 53284
rect 47852 54012 47908 54068
rect 47628 53116 47684 53172
rect 47740 52946 47796 52948
rect 47740 52894 47742 52946
rect 47742 52894 47794 52946
rect 47794 52894 47796 52946
rect 47740 52892 47796 52894
rect 48188 53788 48244 53844
rect 48300 53116 48356 53172
rect 48076 53004 48132 53060
rect 47964 52780 48020 52836
rect 47292 52444 47348 52500
rect 46732 51996 46788 52052
rect 46620 49420 46676 49476
rect 46956 49756 47012 49812
rect 47068 49644 47124 49700
rect 47180 49196 47236 49252
rect 49084 56252 49140 56308
rect 48860 54236 48916 54292
rect 48972 54796 49028 54852
rect 49756 56252 49812 56308
rect 50092 56476 50148 56532
rect 50092 56252 50148 56308
rect 49756 56082 49812 56084
rect 49756 56030 49758 56082
rect 49758 56030 49810 56082
rect 49810 56030 49812 56082
rect 49756 56028 49812 56030
rect 49420 55692 49476 55748
rect 49196 55132 49252 55188
rect 51324 58156 51380 58212
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 49868 55244 49924 55300
rect 50316 56252 50372 56308
rect 49308 54796 49364 54852
rect 49980 54572 50036 54628
rect 49084 54290 49140 54292
rect 49084 54238 49086 54290
rect 49086 54238 49138 54290
rect 49138 54238 49140 54290
rect 49084 54236 49140 54238
rect 49308 54124 49364 54180
rect 48188 52668 48244 52724
rect 48300 52220 48356 52276
rect 48076 52108 48132 52164
rect 47964 50988 48020 51044
rect 48636 50876 48692 50932
rect 47292 50316 47348 50372
rect 46284 48972 46340 49028
rect 46060 48748 46116 48804
rect 46284 48018 46340 48020
rect 46284 47966 46286 48018
rect 46286 47966 46338 48018
rect 46338 47966 46340 48018
rect 46284 47964 46340 47966
rect 45836 47292 45892 47348
rect 45836 47068 45892 47124
rect 45948 46956 46004 47012
rect 45612 46786 45668 46788
rect 45612 46734 45614 46786
rect 45614 46734 45666 46786
rect 45666 46734 45668 46786
rect 45612 46732 45668 46734
rect 47180 49026 47236 49028
rect 47180 48974 47182 49026
rect 47182 48974 47234 49026
rect 47234 48974 47236 49026
rect 47180 48972 47236 48974
rect 47068 48860 47124 48916
rect 46620 48188 46676 48244
rect 46060 46732 46116 46788
rect 45724 46508 45780 46564
rect 46732 48076 46788 48132
rect 46844 47404 46900 47460
rect 46060 44716 46116 44772
rect 46172 44434 46228 44436
rect 46172 44382 46174 44434
rect 46174 44382 46226 44434
rect 46226 44382 46228 44434
rect 46172 44380 46228 44382
rect 46732 46060 46788 46116
rect 46956 45836 47012 45892
rect 46508 42530 46564 42532
rect 46508 42478 46510 42530
rect 46510 42478 46562 42530
rect 46562 42478 46564 42530
rect 46508 42476 46564 42478
rect 45724 42028 45780 42084
rect 46060 42028 46116 42084
rect 47404 50428 47460 50484
rect 47516 49644 47572 49700
rect 47740 49810 47796 49812
rect 47740 49758 47742 49810
rect 47742 49758 47794 49810
rect 47794 49758 47796 49810
rect 47740 49756 47796 49758
rect 47964 49308 48020 49364
rect 47740 49196 47796 49252
rect 47740 48914 47796 48916
rect 47740 48862 47742 48914
rect 47742 48862 47794 48914
rect 47794 48862 47796 48914
rect 47740 48860 47796 48862
rect 47628 48748 47684 48804
rect 48188 48748 48244 48804
rect 47740 47964 47796 48020
rect 47516 47740 47572 47796
rect 48076 47628 48132 47684
rect 47516 47458 47572 47460
rect 47516 47406 47518 47458
rect 47518 47406 47570 47458
rect 47570 47406 47572 47458
rect 47516 47404 47572 47406
rect 47516 46956 47572 47012
rect 47068 45724 47124 45780
rect 47516 45948 47572 46004
rect 47180 44940 47236 44996
rect 48524 50316 48580 50372
rect 49084 53452 49140 53508
rect 48972 53228 49028 53284
rect 50092 55020 50148 55076
rect 49532 53452 49588 53508
rect 49420 53116 49476 53172
rect 49308 52892 49364 52948
rect 49196 52556 49252 52612
rect 49196 51378 49252 51380
rect 49196 51326 49198 51378
rect 49198 51326 49250 51378
rect 49250 51326 49252 51378
rect 49196 51324 49252 51326
rect 48972 51266 49028 51268
rect 48972 51214 48974 51266
rect 48974 51214 49026 51266
rect 49026 51214 49028 51266
rect 48972 51212 49028 51214
rect 49196 50316 49252 50372
rect 48860 49308 48916 49364
rect 48972 49644 49028 49700
rect 48748 48914 48804 48916
rect 48748 48862 48750 48914
rect 48750 48862 48802 48914
rect 48802 48862 48804 48914
rect 48748 48860 48804 48862
rect 48748 48412 48804 48468
rect 49532 51324 49588 51380
rect 49420 50818 49476 50820
rect 49420 50766 49422 50818
rect 49422 50766 49474 50818
rect 49474 50766 49476 50818
rect 49420 50764 49476 50766
rect 49756 53730 49812 53732
rect 49756 53678 49758 53730
rect 49758 53678 49810 53730
rect 49810 53678 49812 53730
rect 49756 53676 49812 53678
rect 49980 53340 50036 53396
rect 49868 52780 49924 52836
rect 50092 52556 50148 52612
rect 50204 52668 50260 52724
rect 49980 52162 50036 52164
rect 49980 52110 49982 52162
rect 49982 52110 50034 52162
rect 50034 52110 50036 52162
rect 49980 52108 50036 52110
rect 49756 50706 49812 50708
rect 49756 50654 49758 50706
rect 49758 50654 49810 50706
rect 49810 50654 49812 50706
rect 49756 50652 49812 50654
rect 49980 50652 50036 50708
rect 49980 50482 50036 50484
rect 49980 50430 49982 50482
rect 49982 50430 50034 50482
rect 50034 50430 50036 50482
rect 49980 50428 50036 50430
rect 49644 50204 49700 50260
rect 49980 50204 50036 50260
rect 49756 49868 49812 49924
rect 49308 49138 49364 49140
rect 49308 49086 49310 49138
rect 49310 49086 49362 49138
rect 49362 49086 49364 49138
rect 49308 49084 49364 49086
rect 49196 48748 49252 48804
rect 49196 48524 49252 48580
rect 48300 47404 48356 47460
rect 48188 46786 48244 46788
rect 48188 46734 48190 46786
rect 48190 46734 48242 46786
rect 48242 46734 48244 46786
rect 48188 46732 48244 46734
rect 48076 46620 48132 46676
rect 47852 45890 47908 45892
rect 47852 45838 47854 45890
rect 47854 45838 47906 45890
rect 47906 45838 47908 45890
rect 47852 45836 47908 45838
rect 47628 45218 47684 45220
rect 47628 45166 47630 45218
rect 47630 45166 47682 45218
rect 47682 45166 47684 45218
rect 47628 45164 47684 45166
rect 47740 45106 47796 45108
rect 47740 45054 47742 45106
rect 47742 45054 47794 45106
rect 47794 45054 47796 45106
rect 47740 45052 47796 45054
rect 47404 44716 47460 44772
rect 47964 44716 48020 44772
rect 46732 43596 46788 43652
rect 46956 43372 47012 43428
rect 47180 43426 47236 43428
rect 47180 43374 47182 43426
rect 47182 43374 47234 43426
rect 47234 43374 47236 43426
rect 47180 43372 47236 43374
rect 47068 42140 47124 42196
rect 46844 42028 46900 42084
rect 46508 41692 46564 41748
rect 45500 40236 45556 40292
rect 46060 40962 46116 40964
rect 46060 40910 46062 40962
rect 46062 40910 46114 40962
rect 46114 40910 46116 40962
rect 46060 40908 46116 40910
rect 45724 40572 45780 40628
rect 44268 40012 44324 40068
rect 44940 40012 44996 40068
rect 46060 40348 46116 40404
rect 47628 41858 47684 41860
rect 47628 41806 47630 41858
rect 47630 41806 47682 41858
rect 47682 41806 47684 41858
rect 47628 41804 47684 41806
rect 47068 40684 47124 40740
rect 46844 40012 46900 40068
rect 47292 40908 47348 40964
rect 47404 40684 47460 40740
rect 48300 45612 48356 45668
rect 48076 44268 48132 44324
rect 48188 45164 48244 45220
rect 47964 44044 48020 44100
rect 47852 43596 47908 43652
rect 48188 43708 48244 43764
rect 47852 41970 47908 41972
rect 47852 41918 47854 41970
rect 47854 41918 47906 41970
rect 47906 41918 47908 41970
rect 47852 41916 47908 41918
rect 47740 41132 47796 41188
rect 47852 40796 47908 40852
rect 47404 39676 47460 39732
rect 47292 39506 47348 39508
rect 47292 39454 47294 39506
rect 47294 39454 47346 39506
rect 47346 39454 47348 39506
rect 47292 39452 47348 39454
rect 47404 39394 47460 39396
rect 47404 39342 47406 39394
rect 47406 39342 47458 39394
rect 47458 39342 47460 39394
rect 47404 39340 47460 39342
rect 47516 39228 47572 39284
rect 46508 39058 46564 39060
rect 46508 39006 46510 39058
rect 46510 39006 46562 39058
rect 46562 39006 46564 39058
rect 46508 39004 46564 39006
rect 45052 38780 45108 38836
rect 44940 38162 44996 38164
rect 44940 38110 44942 38162
rect 44942 38110 44994 38162
rect 44994 38110 44996 38162
rect 44940 38108 44996 38110
rect 44716 37884 44772 37940
rect 44268 37436 44324 37492
rect 44380 35980 44436 36036
rect 44268 35644 44324 35700
rect 44268 35308 44324 35364
rect 44156 34130 44212 34132
rect 44156 34078 44158 34130
rect 44158 34078 44210 34130
rect 44210 34078 44212 34130
rect 44156 34076 44212 34078
rect 45836 38834 45892 38836
rect 45836 38782 45838 38834
rect 45838 38782 45890 38834
rect 45890 38782 45892 38834
rect 45836 38780 45892 38782
rect 44940 37212 44996 37268
rect 44828 36482 44884 36484
rect 44828 36430 44830 36482
rect 44830 36430 44882 36482
rect 44882 36430 44884 36482
rect 44828 36428 44884 36430
rect 45164 35868 45220 35924
rect 45276 36540 45332 36596
rect 45052 35810 45108 35812
rect 45052 35758 45054 35810
rect 45054 35758 45106 35810
rect 45106 35758 45108 35810
rect 45052 35756 45108 35758
rect 44940 35644 44996 35700
rect 45164 35532 45220 35588
rect 44492 34076 44548 34132
rect 45724 37772 45780 37828
rect 45836 37378 45892 37380
rect 45836 37326 45838 37378
rect 45838 37326 45890 37378
rect 45890 37326 45892 37378
rect 45836 37324 45892 37326
rect 45724 36764 45780 36820
rect 45612 36428 45668 36484
rect 45612 35644 45668 35700
rect 45612 34636 45668 34692
rect 46172 37212 46228 37268
rect 46172 36594 46228 36596
rect 46172 36542 46174 36594
rect 46174 36542 46226 36594
rect 46226 36542 46228 36594
rect 46172 36540 46228 36542
rect 46396 37212 46452 37268
rect 46060 36204 46116 36260
rect 46396 36204 46452 36260
rect 46732 38556 46788 38612
rect 46956 38780 47012 38836
rect 46732 38332 46788 38388
rect 46620 38108 46676 38164
rect 46844 37436 46900 37492
rect 46620 36988 46676 37044
rect 45836 35420 45892 35476
rect 46844 35810 46900 35812
rect 46844 35758 46846 35810
rect 46846 35758 46898 35810
rect 46898 35758 46900 35810
rect 46844 35756 46900 35758
rect 45836 34300 45892 34356
rect 45724 33964 45780 34020
rect 44156 33346 44212 33348
rect 44156 33294 44158 33346
rect 44158 33294 44210 33346
rect 44210 33294 44212 33346
rect 44156 33292 44212 33294
rect 45836 33740 45892 33796
rect 45836 33404 45892 33460
rect 44044 33068 44100 33124
rect 44268 33180 44324 33236
rect 43820 32172 43876 32228
rect 43596 31890 43652 31892
rect 43596 31838 43598 31890
rect 43598 31838 43650 31890
rect 43650 31838 43652 31890
rect 43596 31836 43652 31838
rect 43708 31724 43764 31780
rect 42476 29484 42532 29540
rect 43372 30156 43428 30212
rect 43932 32060 43988 32116
rect 43932 31836 43988 31892
rect 43932 30434 43988 30436
rect 43932 30382 43934 30434
rect 43934 30382 43986 30434
rect 43986 30382 43988 30434
rect 43932 30380 43988 30382
rect 43820 30044 43876 30100
rect 43372 29932 43428 29988
rect 42700 29036 42756 29092
rect 42700 28476 42756 28532
rect 43148 28082 43204 28084
rect 43148 28030 43150 28082
rect 43150 28030 43202 28082
rect 43202 28030 43204 28082
rect 43148 28028 43204 28030
rect 42252 26290 42308 26292
rect 42252 26238 42254 26290
rect 42254 26238 42306 26290
rect 42306 26238 42308 26290
rect 42252 26236 42308 26238
rect 41916 25004 41972 25060
rect 41804 23772 41860 23828
rect 41692 23714 41748 23716
rect 41692 23662 41694 23714
rect 41694 23662 41746 23714
rect 41746 23662 41748 23714
rect 41692 23660 41748 23662
rect 41580 23548 41636 23604
rect 41356 22988 41412 23044
rect 40684 20412 40740 20468
rect 40684 19740 40740 19796
rect 41804 23436 41860 23492
rect 41692 23324 41748 23380
rect 41804 22540 41860 22596
rect 43596 29260 43652 29316
rect 43932 28700 43988 28756
rect 45724 33346 45780 33348
rect 45724 33294 45726 33346
rect 45726 33294 45778 33346
rect 45778 33294 45780 33346
rect 45724 33292 45780 33294
rect 45052 33180 45108 33236
rect 44716 31836 44772 31892
rect 45388 32562 45444 32564
rect 45388 32510 45390 32562
rect 45390 32510 45442 32562
rect 45442 32510 45444 32562
rect 45388 32508 45444 32510
rect 45164 31836 45220 31892
rect 44156 31666 44212 31668
rect 44156 31614 44158 31666
rect 44158 31614 44210 31666
rect 44210 31614 44212 31666
rect 44156 31612 44212 31614
rect 45276 31500 45332 31556
rect 44828 31218 44884 31220
rect 44828 31166 44830 31218
rect 44830 31166 44882 31218
rect 44882 31166 44884 31218
rect 44828 31164 44884 31166
rect 46508 34636 46564 34692
rect 46844 34354 46900 34356
rect 46844 34302 46846 34354
rect 46846 34302 46898 34354
rect 46898 34302 46900 34354
rect 46844 34300 46900 34302
rect 47180 38050 47236 38052
rect 47180 37998 47182 38050
rect 47182 37998 47234 38050
rect 47234 37998 47236 38050
rect 47180 37996 47236 37998
rect 47292 37938 47348 37940
rect 47292 37886 47294 37938
rect 47294 37886 47346 37938
rect 47346 37886 47348 37938
rect 47292 37884 47348 37886
rect 47964 39618 48020 39620
rect 47964 39566 47966 39618
rect 47966 39566 48018 39618
rect 48018 39566 48020 39618
rect 47964 39564 48020 39566
rect 47964 39058 48020 39060
rect 47964 39006 47966 39058
rect 47966 39006 48018 39058
rect 48018 39006 48020 39058
rect 47964 39004 48020 39006
rect 47628 38946 47684 38948
rect 47628 38894 47630 38946
rect 47630 38894 47682 38946
rect 47682 38894 47684 38946
rect 47628 38892 47684 38894
rect 47740 38780 47796 38836
rect 47516 38556 47572 38612
rect 47516 37660 47572 37716
rect 47180 36876 47236 36932
rect 47180 35698 47236 35700
rect 47180 35646 47182 35698
rect 47182 35646 47234 35698
rect 47234 35646 47236 35698
rect 47180 35644 47236 35646
rect 46956 34188 47012 34244
rect 47180 34130 47236 34132
rect 47180 34078 47182 34130
rect 47182 34078 47234 34130
rect 47234 34078 47236 34130
rect 47180 34076 47236 34078
rect 46284 34018 46340 34020
rect 46284 33966 46286 34018
rect 46286 33966 46338 34018
rect 46338 33966 46340 34018
rect 46284 33964 46340 33966
rect 47068 33516 47124 33572
rect 46844 33234 46900 33236
rect 46844 33182 46846 33234
rect 46846 33182 46898 33234
rect 46898 33182 46900 33234
rect 46844 33180 46900 33182
rect 46508 31948 46564 32004
rect 46284 31836 46340 31892
rect 46060 31554 46116 31556
rect 46060 31502 46062 31554
rect 46062 31502 46114 31554
rect 46114 31502 46116 31554
rect 46060 31500 46116 31502
rect 45948 31164 46004 31220
rect 46284 31164 46340 31220
rect 44380 30828 44436 30884
rect 44156 30210 44212 30212
rect 44156 30158 44158 30210
rect 44158 30158 44210 30210
rect 44210 30158 44212 30210
rect 44156 30156 44212 30158
rect 44156 29148 44212 29204
rect 43820 27580 43876 27636
rect 42588 25676 42644 25732
rect 42700 27132 42756 27188
rect 42588 25506 42644 25508
rect 42588 25454 42590 25506
rect 42590 25454 42642 25506
rect 42642 25454 42644 25506
rect 42588 25452 42644 25454
rect 43148 27186 43204 27188
rect 43148 27134 43150 27186
rect 43150 27134 43202 27186
rect 43202 27134 43204 27186
rect 43148 27132 43204 27134
rect 42812 26908 42868 26964
rect 42476 23548 42532 23604
rect 42028 23212 42084 23268
rect 42364 23154 42420 23156
rect 42364 23102 42366 23154
rect 42366 23102 42418 23154
rect 42418 23102 42420 23154
rect 42364 23100 42420 23102
rect 42140 21810 42196 21812
rect 42140 21758 42142 21810
rect 42142 21758 42194 21810
rect 42194 21758 42196 21810
rect 42140 21756 42196 21758
rect 41468 21644 41524 21700
rect 40124 15820 40180 15876
rect 41244 19516 41300 19572
rect 39228 14530 39284 14532
rect 39228 14478 39230 14530
rect 39230 14478 39282 14530
rect 39282 14478 39284 14530
rect 39228 14476 39284 14478
rect 39452 14924 39508 14980
rect 39452 14364 39508 14420
rect 39564 14140 39620 14196
rect 39564 13468 39620 13524
rect 39228 12908 39284 12964
rect 39228 12684 39284 12740
rect 38668 11676 38724 11732
rect 39116 12460 39172 12516
rect 38892 12178 38948 12180
rect 38892 12126 38894 12178
rect 38894 12126 38946 12178
rect 38946 12126 38948 12178
rect 38892 12124 38948 12126
rect 38668 9548 38724 9604
rect 38892 9324 38948 9380
rect 38780 9100 38836 9156
rect 38444 5906 38500 5908
rect 38444 5854 38446 5906
rect 38446 5854 38498 5906
rect 38498 5854 38500 5906
rect 38444 5852 38500 5854
rect 38332 5516 38388 5572
rect 37548 4284 37604 4340
rect 38332 5068 38388 5124
rect 35532 3276 35588 3332
rect 36316 3276 36372 3332
rect 38668 8764 38724 8820
rect 39004 8652 39060 8708
rect 40012 14700 40068 14756
rect 39900 14588 39956 14644
rect 40012 13580 40068 13636
rect 40348 14812 40404 14868
rect 40348 13916 40404 13972
rect 40236 13522 40292 13524
rect 40236 13470 40238 13522
rect 40238 13470 40290 13522
rect 40290 13470 40292 13522
rect 40236 13468 40292 13470
rect 40124 13020 40180 13076
rect 39676 12348 39732 12404
rect 40460 12908 40516 12964
rect 41356 20300 41412 20356
rect 41020 19180 41076 19236
rect 40796 17948 40852 18004
rect 40796 17554 40852 17556
rect 40796 17502 40798 17554
rect 40798 17502 40850 17554
rect 40850 17502 40852 17554
rect 40796 17500 40852 17502
rect 42028 21586 42084 21588
rect 42028 21534 42030 21586
rect 42030 21534 42082 21586
rect 42082 21534 42084 21586
rect 42028 21532 42084 21534
rect 42364 21698 42420 21700
rect 42364 21646 42366 21698
rect 42366 21646 42418 21698
rect 42418 21646 42420 21698
rect 42364 21644 42420 21646
rect 43484 26962 43540 26964
rect 43484 26910 43486 26962
rect 43486 26910 43538 26962
rect 43538 26910 43540 26962
rect 43484 26908 43540 26910
rect 43372 26796 43428 26852
rect 42924 26572 42980 26628
rect 42924 24108 42980 24164
rect 43148 25004 43204 25060
rect 43036 23436 43092 23492
rect 43036 21868 43092 21924
rect 43260 23100 43316 23156
rect 43260 22316 43316 22372
rect 43148 21756 43204 21812
rect 41692 20188 41748 20244
rect 41804 20300 41860 20356
rect 41580 19628 41636 19684
rect 41132 17666 41188 17668
rect 41132 17614 41134 17666
rect 41134 17614 41186 17666
rect 41186 17614 41188 17666
rect 41132 17612 41188 17614
rect 41356 17500 41412 17556
rect 42140 20748 42196 20804
rect 43036 20802 43092 20804
rect 43036 20750 43038 20802
rect 43038 20750 43090 20802
rect 43090 20750 43092 20802
rect 43036 20748 43092 20750
rect 42252 20300 42308 20356
rect 42364 20524 42420 20580
rect 42252 19346 42308 19348
rect 42252 19294 42254 19346
rect 42254 19294 42306 19346
rect 42306 19294 42308 19346
rect 42252 19292 42308 19294
rect 42140 18450 42196 18452
rect 42140 18398 42142 18450
rect 42142 18398 42194 18450
rect 42194 18398 42196 18450
rect 42140 18396 42196 18398
rect 42252 17554 42308 17556
rect 42252 17502 42254 17554
rect 42254 17502 42306 17554
rect 42306 17502 42308 17554
rect 42252 17500 42308 17502
rect 41132 16882 41188 16884
rect 41132 16830 41134 16882
rect 41134 16830 41186 16882
rect 41186 16830 41188 16882
rect 41132 16828 41188 16830
rect 40684 16716 40740 16772
rect 41468 16210 41524 16212
rect 41468 16158 41470 16210
rect 41470 16158 41522 16210
rect 41522 16158 41524 16210
rect 41468 16156 41524 16158
rect 40796 14924 40852 14980
rect 40908 14588 40964 14644
rect 41468 15148 41524 15204
rect 42028 16044 42084 16100
rect 42924 20524 42980 20580
rect 43820 26908 43876 26964
rect 43708 26236 43764 26292
rect 43820 26572 43876 26628
rect 43596 25228 43652 25284
rect 43484 22428 43540 22484
rect 43596 23772 43652 23828
rect 43596 21980 43652 22036
rect 45052 29986 45108 29988
rect 45052 29934 45054 29986
rect 45054 29934 45106 29986
rect 45106 29934 45108 29986
rect 45052 29932 45108 29934
rect 46060 29986 46116 29988
rect 46060 29934 46062 29986
rect 46062 29934 46114 29986
rect 46114 29934 46116 29986
rect 46060 29932 46116 29934
rect 46060 29372 46116 29428
rect 48636 46956 48692 47012
rect 48748 47068 48804 47124
rect 48972 46956 49028 47012
rect 49420 47964 49476 48020
rect 49420 47180 49476 47236
rect 49420 46844 49476 46900
rect 49532 46732 49588 46788
rect 49868 49026 49924 49028
rect 49868 48974 49870 49026
rect 49870 48974 49922 49026
rect 49922 48974 49924 49026
rect 49868 48972 49924 48974
rect 49868 48300 49924 48356
rect 50540 55356 50596 55412
rect 50988 56028 51044 56084
rect 51100 57260 51156 57316
rect 50876 55020 50932 55076
rect 50988 55356 51044 55412
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50876 54684 50932 54740
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50316 52108 50372 52164
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 51212 55074 51268 55076
rect 51212 55022 51214 55074
rect 51214 55022 51266 55074
rect 51266 55022 51268 55074
rect 51212 55020 51268 55022
rect 51212 53618 51268 53620
rect 51212 53566 51214 53618
rect 51214 53566 51266 53618
rect 51266 53566 51268 53618
rect 51212 53564 51268 53566
rect 51436 55356 51492 55412
rect 51436 53452 51492 53508
rect 50988 52946 51044 52948
rect 50988 52894 50990 52946
rect 50990 52894 51042 52946
rect 51042 52894 51044 52946
rect 50988 52892 51044 52894
rect 50204 50092 50260 50148
rect 50316 51436 50372 51492
rect 50764 50764 50820 50820
rect 50988 50594 51044 50596
rect 50988 50542 50990 50594
rect 50990 50542 51042 50594
rect 51042 50542 51044 50594
rect 50988 50540 51044 50542
rect 50428 50370 50484 50372
rect 50428 50318 50430 50370
rect 50430 50318 50482 50370
rect 50482 50318 50484 50370
rect 50428 50316 50484 50318
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50204 49868 50260 49924
rect 50428 49196 50484 49252
rect 50988 50092 51044 50148
rect 51660 58210 51716 58212
rect 51660 58158 51662 58210
rect 51662 58158 51714 58210
rect 51714 58158 51716 58210
rect 51660 58156 51716 58158
rect 52108 57762 52164 57764
rect 52108 57710 52110 57762
rect 52110 57710 52162 57762
rect 52162 57710 52164 57762
rect 52108 57708 52164 57710
rect 51884 57596 51940 57652
rect 51660 56306 51716 56308
rect 51660 56254 51662 56306
rect 51662 56254 51714 56306
rect 51714 56254 51716 56306
rect 51660 56252 51716 56254
rect 51660 54908 51716 54964
rect 51660 54514 51716 54516
rect 51660 54462 51662 54514
rect 51662 54462 51714 54514
rect 51714 54462 51716 54514
rect 51660 54460 51716 54462
rect 51660 53618 51716 53620
rect 51660 53566 51662 53618
rect 51662 53566 51714 53618
rect 51714 53566 51716 53618
rect 51660 53564 51716 53566
rect 52332 57372 52388 57428
rect 52220 55580 52276 55636
rect 51996 55074 52052 55076
rect 51996 55022 51998 55074
rect 51998 55022 52050 55074
rect 52050 55022 52052 55074
rect 51996 55020 52052 55022
rect 52108 54626 52164 54628
rect 52108 54574 52110 54626
rect 52110 54574 52162 54626
rect 52162 54574 52164 54626
rect 52108 54572 52164 54574
rect 51884 53788 51940 53844
rect 52108 54348 52164 54404
rect 51548 52668 51604 52724
rect 51324 52332 51380 52388
rect 51212 50652 51268 50708
rect 51324 52108 51380 52164
rect 50876 49084 50932 49140
rect 50764 49026 50820 49028
rect 50764 48974 50766 49026
rect 50766 48974 50818 49026
rect 50818 48974 50820 49026
rect 50764 48972 50820 48974
rect 51100 48748 51156 48804
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50876 48354 50932 48356
rect 50876 48302 50878 48354
rect 50878 48302 50930 48354
rect 50930 48302 50932 48354
rect 50876 48300 50932 48302
rect 49196 45948 49252 46004
rect 48860 45218 48916 45220
rect 48860 45166 48862 45218
rect 48862 45166 48914 45218
rect 48914 45166 48916 45218
rect 48860 45164 48916 45166
rect 48972 45106 49028 45108
rect 48972 45054 48974 45106
rect 48974 45054 49026 45106
rect 49026 45054 49028 45106
rect 48972 45052 49028 45054
rect 48860 44492 48916 44548
rect 48524 43596 48580 43652
rect 48748 44098 48804 44100
rect 48748 44046 48750 44098
rect 48750 44046 48802 44098
rect 48802 44046 48804 44098
rect 48748 44044 48804 44046
rect 48412 42140 48468 42196
rect 48748 43820 48804 43876
rect 49756 45948 49812 46004
rect 49532 45164 49588 45220
rect 49868 45164 49924 45220
rect 50652 47740 50708 47796
rect 50204 47346 50260 47348
rect 50204 47294 50206 47346
rect 50206 47294 50258 47346
rect 50258 47294 50260 47346
rect 50204 47292 50260 47294
rect 50316 46956 50372 47012
rect 50092 45890 50148 45892
rect 50092 45838 50094 45890
rect 50094 45838 50146 45890
rect 50146 45838 50148 45890
rect 50092 45836 50148 45838
rect 50204 46844 50260 46900
rect 50092 45500 50148 45556
rect 48860 42252 48916 42308
rect 49084 43036 49140 43092
rect 49196 43708 49252 43764
rect 48972 41804 49028 41860
rect 48972 41020 49028 41076
rect 48860 40236 48916 40292
rect 48748 39564 48804 39620
rect 49084 40012 49140 40068
rect 48748 38946 48804 38948
rect 48748 38894 48750 38946
rect 48750 38894 48802 38946
rect 48802 38894 48804 38946
rect 48748 38892 48804 38894
rect 49308 43650 49364 43652
rect 49308 43598 49310 43650
rect 49310 43598 49362 43650
rect 49362 43598 49364 43650
rect 49308 43596 49364 43598
rect 49308 43372 49364 43428
rect 49420 42082 49476 42084
rect 49420 42030 49422 42082
rect 49422 42030 49474 42082
rect 49474 42030 49476 42082
rect 49420 42028 49476 42030
rect 49644 44210 49700 44212
rect 49644 44158 49646 44210
rect 49646 44158 49698 44210
rect 49698 44158 49700 44210
rect 49644 44156 49700 44158
rect 49756 44492 49812 44548
rect 50876 47852 50932 47908
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50428 46396 50484 46452
rect 50316 46060 50372 46116
rect 50428 45948 50484 46004
rect 50764 46060 50820 46116
rect 51548 50764 51604 50820
rect 51436 50652 51492 50708
rect 51436 50316 51492 50372
rect 51884 50482 51940 50484
rect 51884 50430 51886 50482
rect 51886 50430 51938 50482
rect 51938 50430 51940 50482
rect 51884 50428 51940 50430
rect 51660 50092 51716 50148
rect 51772 50204 51828 50260
rect 51660 49532 51716 49588
rect 62188 58492 62244 58548
rect 52892 57650 52948 57652
rect 52892 57598 52894 57650
rect 52894 57598 52946 57650
rect 52946 57598 52948 57650
rect 52892 57596 52948 57598
rect 52780 57538 52836 57540
rect 52780 57486 52782 57538
rect 52782 57486 52834 57538
rect 52834 57486 52836 57538
rect 52780 57484 52836 57486
rect 53116 57260 53172 57316
rect 53788 57708 53844 57764
rect 53228 57596 53284 57652
rect 52444 54348 52500 54404
rect 52444 54124 52500 54180
rect 52892 56642 52948 56644
rect 52892 56590 52894 56642
rect 52894 56590 52946 56642
rect 52946 56590 52948 56642
rect 52892 56588 52948 56590
rect 54012 57650 54068 57652
rect 54012 57598 54014 57650
rect 54014 57598 54066 57650
rect 54066 57598 54068 57650
rect 54012 57596 54068 57598
rect 53564 57372 53620 57428
rect 52668 54684 52724 54740
rect 52780 54626 52836 54628
rect 52780 54574 52782 54626
rect 52782 54574 52834 54626
rect 52834 54574 52836 54626
rect 52780 54572 52836 54574
rect 53676 57260 53732 57316
rect 53788 56252 53844 56308
rect 55356 57820 55412 57876
rect 55020 57538 55076 57540
rect 55020 57486 55022 57538
rect 55022 57486 55074 57538
rect 55074 57486 55076 57538
rect 55020 57484 55076 57486
rect 53228 55298 53284 55300
rect 53228 55246 53230 55298
rect 53230 55246 53282 55298
rect 53282 55246 53284 55298
rect 53228 55244 53284 55246
rect 53452 55020 53508 55076
rect 53900 55298 53956 55300
rect 53900 55246 53902 55298
rect 53902 55246 53954 55298
rect 53954 55246 53956 55298
rect 53900 55244 53956 55246
rect 53676 55020 53732 55076
rect 53564 54908 53620 54964
rect 53228 54348 53284 54404
rect 52892 54236 52948 54292
rect 53676 54572 53732 54628
rect 52892 53676 52948 53732
rect 52556 53564 52612 53620
rect 52668 53116 52724 53172
rect 52220 52220 52276 52276
rect 52892 52444 52948 52500
rect 52108 51436 52164 51492
rect 52444 51884 52500 51940
rect 52108 51100 52164 51156
rect 51996 49084 52052 49140
rect 51772 48802 51828 48804
rect 51772 48750 51774 48802
rect 51774 48750 51826 48802
rect 51826 48750 51828 48802
rect 51772 48748 51828 48750
rect 51324 48130 51380 48132
rect 51324 48078 51326 48130
rect 51326 48078 51378 48130
rect 51378 48078 51380 48130
rect 51324 48076 51380 48078
rect 51436 47740 51492 47796
rect 51212 47628 51268 47684
rect 51772 48242 51828 48244
rect 51772 48190 51774 48242
rect 51774 48190 51826 48242
rect 51826 48190 51828 48242
rect 51772 48188 51828 48190
rect 51324 47570 51380 47572
rect 51324 47518 51326 47570
rect 51326 47518 51378 47570
rect 51378 47518 51380 47570
rect 51324 47516 51380 47518
rect 52780 52162 52836 52164
rect 52780 52110 52782 52162
rect 52782 52110 52834 52162
rect 52834 52110 52836 52162
rect 52780 52108 52836 52110
rect 53228 52668 53284 52724
rect 53228 52444 53284 52500
rect 53004 51324 53060 51380
rect 52556 49644 52612 49700
rect 53788 54514 53844 54516
rect 53788 54462 53790 54514
rect 53790 54462 53842 54514
rect 53842 54462 53844 54514
rect 53788 54460 53844 54462
rect 53788 53676 53844 53732
rect 53900 53116 53956 53172
rect 53452 52892 53508 52948
rect 53676 51938 53732 51940
rect 53676 51886 53678 51938
rect 53678 51886 53730 51938
rect 53730 51886 53732 51938
rect 53676 51884 53732 51886
rect 53228 50706 53284 50708
rect 53228 50654 53230 50706
rect 53230 50654 53282 50706
rect 53282 50654 53284 50706
rect 53228 50652 53284 50654
rect 53564 50988 53620 51044
rect 53564 50540 53620 50596
rect 53116 49868 53172 49924
rect 53228 49980 53284 50036
rect 52892 49196 52948 49252
rect 52780 49138 52836 49140
rect 52780 49086 52782 49138
rect 52782 49086 52834 49138
rect 52834 49086 52836 49138
rect 52780 49084 52836 49086
rect 52556 48860 52612 48916
rect 52444 47516 52500 47572
rect 51436 46732 51492 46788
rect 51212 46172 51268 46228
rect 51436 46060 51492 46116
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50316 45106 50372 45108
rect 50316 45054 50318 45106
rect 50318 45054 50370 45106
rect 50370 45054 50372 45106
rect 50316 45052 50372 45054
rect 50428 44322 50484 44324
rect 50428 44270 50430 44322
rect 50430 44270 50482 44322
rect 50482 44270 50484 44322
rect 50428 44268 50484 44270
rect 50652 44380 50708 44436
rect 51100 45052 51156 45108
rect 51212 45836 51268 45892
rect 50204 43596 50260 43652
rect 50652 44044 50708 44100
rect 50092 41916 50148 41972
rect 50316 42028 50372 42084
rect 49868 41074 49924 41076
rect 49868 41022 49870 41074
rect 49870 41022 49922 41074
rect 49922 41022 49924 41074
rect 49868 41020 49924 41022
rect 49980 40514 50036 40516
rect 49980 40462 49982 40514
rect 49982 40462 50034 40514
rect 50034 40462 50036 40514
rect 49980 40460 50036 40462
rect 49644 40124 49700 40180
rect 49756 40348 49812 40404
rect 48076 38220 48132 38276
rect 48188 38556 48244 38612
rect 47964 38108 48020 38164
rect 47852 37772 47908 37828
rect 48076 37996 48132 38052
rect 48412 38444 48468 38500
rect 48748 38108 48804 38164
rect 47852 36652 47908 36708
rect 48188 36764 48244 36820
rect 48412 37772 48468 37828
rect 49420 38668 49476 38724
rect 49532 38780 49588 38836
rect 49308 37996 49364 38052
rect 49532 37884 49588 37940
rect 48972 37660 49028 37716
rect 48860 37490 48916 37492
rect 48860 37438 48862 37490
rect 48862 37438 48914 37490
rect 48914 37438 48916 37490
rect 48860 37436 48916 37438
rect 49420 37378 49476 37380
rect 49420 37326 49422 37378
rect 49422 37326 49474 37378
rect 49474 37326 49476 37378
rect 49420 37324 49476 37326
rect 48748 36988 48804 37044
rect 49308 36988 49364 37044
rect 49084 36652 49140 36708
rect 48076 36092 48132 36148
rect 47628 35810 47684 35812
rect 47628 35758 47630 35810
rect 47630 35758 47682 35810
rect 47682 35758 47684 35810
rect 47628 35756 47684 35758
rect 47852 35698 47908 35700
rect 47852 35646 47854 35698
rect 47854 35646 47906 35698
rect 47906 35646 47908 35698
rect 47852 35644 47908 35646
rect 47740 35586 47796 35588
rect 47740 35534 47742 35586
rect 47742 35534 47794 35586
rect 47794 35534 47796 35586
rect 47740 35532 47796 35534
rect 47404 33458 47460 33460
rect 47404 33406 47406 33458
rect 47406 33406 47458 33458
rect 47458 33406 47460 33458
rect 47404 33404 47460 33406
rect 47852 33122 47908 33124
rect 47852 33070 47854 33122
rect 47854 33070 47906 33122
rect 47906 33070 47908 33122
rect 47852 33068 47908 33070
rect 46620 30380 46676 30436
rect 46732 30492 46788 30548
rect 47404 30268 47460 30324
rect 46396 29932 46452 29988
rect 44716 29314 44772 29316
rect 44716 29262 44718 29314
rect 44718 29262 44770 29314
rect 44770 29262 44772 29314
rect 44716 29260 44772 29262
rect 45836 29260 45892 29316
rect 45276 29202 45332 29204
rect 45276 29150 45278 29202
rect 45278 29150 45330 29202
rect 45330 29150 45332 29202
rect 45276 29148 45332 29150
rect 44044 26012 44100 26068
rect 43932 23324 43988 23380
rect 44268 25506 44324 25508
rect 44268 25454 44270 25506
rect 44270 25454 44322 25506
rect 44322 25454 44324 25506
rect 44268 25452 44324 25454
rect 45164 28252 45220 28308
rect 44828 26962 44884 26964
rect 44828 26910 44830 26962
rect 44830 26910 44882 26962
rect 44882 26910 44884 26962
rect 44828 26908 44884 26910
rect 44828 26684 44884 26740
rect 45948 28588 46004 28644
rect 45948 28140 46004 28196
rect 46956 30156 47012 30212
rect 46508 29314 46564 29316
rect 46508 29262 46510 29314
rect 46510 29262 46562 29314
rect 46562 29262 46564 29314
rect 46508 29260 46564 29262
rect 46060 27804 46116 27860
rect 46732 29148 46788 29204
rect 46732 28924 46788 28980
rect 47628 31218 47684 31220
rect 47628 31166 47630 31218
rect 47630 31166 47682 31218
rect 47682 31166 47684 31218
rect 47628 31164 47684 31166
rect 48860 35474 48916 35476
rect 48860 35422 48862 35474
rect 48862 35422 48914 35474
rect 48914 35422 48916 35474
rect 48860 35420 48916 35422
rect 48748 34860 48804 34916
rect 48188 34300 48244 34356
rect 48188 33906 48244 33908
rect 48188 33854 48190 33906
rect 48190 33854 48242 33906
rect 48242 33854 48244 33906
rect 48188 33852 48244 33854
rect 49420 36652 49476 36708
rect 49308 35308 49364 35364
rect 49420 35644 49476 35700
rect 49196 35196 49252 35252
rect 49084 34242 49140 34244
rect 49084 34190 49086 34242
rect 49086 34190 49138 34242
rect 49138 34190 49140 34242
rect 49084 34188 49140 34190
rect 48972 33852 49028 33908
rect 48860 33404 48916 33460
rect 48076 33180 48132 33236
rect 48748 33234 48804 33236
rect 48748 33182 48750 33234
rect 48750 33182 48802 33234
rect 48802 33182 48804 33234
rect 48748 33180 48804 33182
rect 48300 32284 48356 32340
rect 48188 31554 48244 31556
rect 48188 31502 48190 31554
rect 48190 31502 48242 31554
rect 48242 31502 48244 31554
rect 48188 31500 48244 31502
rect 47628 30156 47684 30212
rect 47292 29426 47348 29428
rect 47292 29374 47294 29426
rect 47294 29374 47346 29426
rect 47346 29374 47348 29426
rect 47292 29372 47348 29374
rect 47852 29426 47908 29428
rect 47852 29374 47854 29426
rect 47854 29374 47906 29426
rect 47906 29374 47908 29426
rect 47852 29372 47908 29374
rect 47180 29148 47236 29204
rect 46956 28700 47012 28756
rect 46732 27858 46788 27860
rect 46732 27806 46734 27858
rect 46734 27806 46786 27858
rect 46786 27806 46788 27858
rect 46732 27804 46788 27806
rect 45612 27298 45668 27300
rect 45612 27246 45614 27298
rect 45614 27246 45666 27298
rect 45666 27246 45668 27298
rect 45612 27244 45668 27246
rect 46172 27074 46228 27076
rect 46172 27022 46174 27074
rect 46174 27022 46226 27074
rect 46226 27022 46228 27074
rect 46172 27020 46228 27022
rect 46396 27634 46452 27636
rect 46396 27582 46398 27634
rect 46398 27582 46450 27634
rect 46450 27582 46452 27634
rect 46396 27580 46452 27582
rect 46508 27468 46564 27524
rect 45164 26572 45220 26628
rect 45052 25676 45108 25732
rect 45276 26236 45332 26292
rect 45164 25618 45220 25620
rect 45164 25566 45166 25618
rect 45166 25566 45218 25618
rect 45218 25566 45220 25618
rect 45164 25564 45220 25566
rect 44604 25116 44660 25172
rect 44940 25228 44996 25284
rect 44268 24668 44324 24724
rect 44380 24162 44436 24164
rect 44380 24110 44382 24162
rect 44382 24110 44434 24162
rect 44434 24110 44436 24162
rect 44380 24108 44436 24110
rect 43820 21698 43876 21700
rect 43820 21646 43822 21698
rect 43822 21646 43874 21698
rect 43874 21646 43876 21698
rect 43820 21644 43876 21646
rect 43596 21586 43652 21588
rect 43596 21534 43598 21586
rect 43598 21534 43650 21586
rect 43650 21534 43652 21586
rect 43596 21532 43652 21534
rect 43148 20300 43204 20356
rect 43484 20748 43540 20804
rect 43036 19516 43092 19572
rect 42700 18620 42756 18676
rect 42812 18508 42868 18564
rect 42700 18450 42756 18452
rect 42700 18398 42702 18450
rect 42702 18398 42754 18450
rect 42754 18398 42756 18450
rect 42700 18396 42756 18398
rect 43036 18338 43092 18340
rect 43036 18286 43038 18338
rect 43038 18286 43090 18338
rect 43090 18286 43092 18338
rect 43036 18284 43092 18286
rect 43148 18172 43204 18228
rect 42812 18060 42868 18116
rect 42476 16716 42532 16772
rect 42476 16044 42532 16100
rect 41804 15538 41860 15540
rect 41804 15486 41806 15538
rect 41806 15486 41858 15538
rect 41858 15486 41860 15538
rect 41804 15484 41860 15486
rect 41692 15426 41748 15428
rect 41692 15374 41694 15426
rect 41694 15374 41746 15426
rect 41746 15374 41748 15426
rect 41692 15372 41748 15374
rect 42028 15314 42084 15316
rect 42028 15262 42030 15314
rect 42030 15262 42082 15314
rect 42082 15262 42084 15314
rect 42028 15260 42084 15262
rect 41916 14924 41972 14980
rect 42140 14700 42196 14756
rect 42252 15148 42308 15204
rect 42588 15484 42644 15540
rect 42812 15986 42868 15988
rect 42812 15934 42814 15986
rect 42814 15934 42866 15986
rect 42866 15934 42868 15986
rect 42812 15932 42868 15934
rect 42924 15426 42980 15428
rect 42924 15374 42926 15426
rect 42926 15374 42978 15426
rect 42978 15374 42980 15426
rect 42924 15372 42980 15374
rect 42812 15260 42868 15316
rect 41020 14364 41076 14420
rect 41132 14306 41188 14308
rect 41132 14254 41134 14306
rect 41134 14254 41186 14306
rect 41186 14254 41188 14306
rect 41132 14252 41188 14254
rect 41132 13692 41188 13748
rect 40796 13580 40852 13636
rect 40684 13074 40740 13076
rect 40684 13022 40686 13074
rect 40686 13022 40738 13074
rect 40738 13022 40740 13074
rect 40684 13020 40740 13022
rect 40684 12796 40740 12852
rect 39900 9884 39956 9940
rect 39676 9602 39732 9604
rect 39676 9550 39678 9602
rect 39678 9550 39730 9602
rect 39730 9550 39732 9602
rect 39676 9548 39732 9550
rect 39564 9100 39620 9156
rect 39340 8988 39396 9044
rect 39900 8988 39956 9044
rect 40348 9996 40404 10052
rect 40124 9212 40180 9268
rect 40124 9042 40180 9044
rect 40124 8990 40126 9042
rect 40126 8990 40178 9042
rect 40178 8990 40180 9042
rect 40124 8988 40180 8990
rect 39564 8930 39620 8932
rect 39564 8878 39566 8930
rect 39566 8878 39618 8930
rect 39618 8878 39620 8930
rect 39564 8876 39620 8878
rect 39004 8092 39060 8148
rect 39228 7980 39284 8036
rect 38780 5292 38836 5348
rect 38444 4844 38500 4900
rect 38668 4844 38724 4900
rect 38332 3500 38388 3556
rect 39340 7586 39396 7588
rect 39340 7534 39342 7586
rect 39342 7534 39394 7586
rect 39394 7534 39396 7586
rect 39340 7532 39396 7534
rect 39340 6972 39396 7028
rect 39340 6748 39396 6804
rect 39228 6578 39284 6580
rect 39228 6526 39230 6578
rect 39230 6526 39282 6578
rect 39282 6526 39284 6578
rect 39228 6524 39284 6526
rect 39900 8764 39956 8820
rect 40572 10780 40628 10836
rect 41356 14418 41412 14420
rect 41356 14366 41358 14418
rect 41358 14366 41410 14418
rect 41410 14366 41412 14418
rect 41356 14364 41412 14366
rect 41356 13580 41412 13636
rect 42588 14530 42644 14532
rect 42588 14478 42590 14530
rect 42590 14478 42642 14530
rect 42642 14478 42644 14530
rect 42588 14476 42644 14478
rect 41916 13580 41972 13636
rect 41468 12962 41524 12964
rect 41468 12910 41470 12962
rect 41470 12910 41522 12962
rect 41522 12910 41524 12962
rect 41468 12908 41524 12910
rect 41468 12402 41524 12404
rect 41468 12350 41470 12402
rect 41470 12350 41522 12402
rect 41522 12350 41524 12402
rect 41468 12348 41524 12350
rect 41244 12290 41300 12292
rect 41244 12238 41246 12290
rect 41246 12238 41298 12290
rect 41298 12238 41300 12290
rect 41244 12236 41300 12238
rect 41132 11564 41188 11620
rect 41692 12124 41748 12180
rect 41244 11394 41300 11396
rect 41244 11342 41246 11394
rect 41246 11342 41298 11394
rect 41298 11342 41300 11394
rect 41244 11340 41300 11342
rect 42028 12124 42084 12180
rect 41804 11788 41860 11844
rect 40908 11004 40964 11060
rect 40684 9884 40740 9940
rect 41356 10610 41412 10612
rect 41356 10558 41358 10610
rect 41358 10558 41410 10610
rect 41410 10558 41412 10610
rect 41356 10556 41412 10558
rect 43820 20578 43876 20580
rect 43820 20526 43822 20578
rect 43822 20526 43874 20578
rect 43874 20526 43876 20578
rect 43820 20524 43876 20526
rect 44604 23266 44660 23268
rect 44604 23214 44606 23266
rect 44606 23214 44658 23266
rect 44658 23214 44660 23266
rect 44604 23212 44660 23214
rect 45052 24722 45108 24724
rect 45052 24670 45054 24722
rect 45054 24670 45106 24722
rect 45106 24670 45108 24722
rect 45052 24668 45108 24670
rect 45612 26124 45668 26180
rect 45500 26066 45556 26068
rect 45500 26014 45502 26066
rect 45502 26014 45554 26066
rect 45554 26014 45556 26066
rect 45500 26012 45556 26014
rect 45388 25788 45444 25844
rect 45500 25228 45556 25284
rect 44716 22764 44772 22820
rect 45052 23548 45108 23604
rect 44940 23154 44996 23156
rect 44940 23102 44942 23154
rect 44942 23102 44994 23154
rect 44994 23102 44996 23154
rect 44940 23100 44996 23102
rect 44828 22540 44884 22596
rect 45388 24668 45444 24724
rect 45276 22482 45332 22484
rect 45276 22430 45278 22482
rect 45278 22430 45330 22482
rect 45330 22430 45332 22482
rect 45276 22428 45332 22430
rect 44828 22370 44884 22372
rect 44828 22318 44830 22370
rect 44830 22318 44882 22370
rect 44882 22318 44884 22370
rect 44828 22316 44884 22318
rect 44492 21810 44548 21812
rect 44492 21758 44494 21810
rect 44494 21758 44546 21810
rect 44546 21758 44548 21810
rect 44492 21756 44548 21758
rect 44380 21532 44436 21588
rect 48188 30994 48244 30996
rect 48188 30942 48190 30994
rect 48190 30942 48242 30994
rect 48242 30942 48244 30994
rect 48188 30940 48244 30942
rect 48076 30604 48132 30660
rect 48076 29538 48132 29540
rect 48076 29486 48078 29538
rect 48078 29486 48130 29538
rect 48130 29486 48132 29538
rect 48076 29484 48132 29486
rect 47180 28028 47236 28084
rect 47292 28140 47348 28196
rect 46508 26460 46564 26516
rect 46060 26348 46116 26404
rect 46060 25730 46116 25732
rect 46060 25678 46062 25730
rect 46062 25678 46114 25730
rect 46114 25678 46116 25730
rect 46060 25676 46116 25678
rect 46620 26012 46676 26068
rect 46172 25394 46228 25396
rect 46172 25342 46174 25394
rect 46174 25342 46226 25394
rect 46226 25342 46228 25394
rect 46172 25340 46228 25342
rect 46396 25788 46452 25844
rect 45612 23212 45668 23268
rect 45948 23212 46004 23268
rect 44716 21644 44772 21700
rect 45052 21586 45108 21588
rect 45052 21534 45054 21586
rect 45054 21534 45106 21586
rect 45106 21534 45108 21586
rect 45052 21532 45108 21534
rect 45836 22482 45892 22484
rect 45836 22430 45838 22482
rect 45838 22430 45890 22482
rect 45890 22430 45892 22482
rect 45836 22428 45892 22430
rect 45836 21810 45892 21812
rect 45836 21758 45838 21810
rect 45838 21758 45890 21810
rect 45890 21758 45892 21810
rect 45836 21756 45892 21758
rect 45724 21586 45780 21588
rect 45724 21534 45726 21586
rect 45726 21534 45778 21586
rect 45778 21534 45780 21586
rect 45724 21532 45780 21534
rect 44156 21084 44212 21140
rect 45948 20860 46004 20916
rect 45164 20802 45220 20804
rect 45164 20750 45166 20802
rect 45166 20750 45218 20802
rect 45218 20750 45220 20802
rect 45164 20748 45220 20750
rect 45612 20748 45668 20804
rect 44156 20242 44212 20244
rect 44156 20190 44158 20242
rect 44158 20190 44210 20242
rect 44210 20190 44212 20242
rect 44156 20188 44212 20190
rect 43596 18338 43652 18340
rect 43596 18286 43598 18338
rect 43598 18286 43650 18338
rect 43650 18286 43652 18338
rect 43596 18284 43652 18286
rect 43708 18172 43764 18228
rect 43932 19010 43988 19012
rect 43932 18958 43934 19010
rect 43934 18958 43986 19010
rect 43986 18958 43988 19010
rect 43932 18956 43988 18958
rect 45500 20018 45556 20020
rect 45500 19966 45502 20018
rect 45502 19966 45554 20018
rect 45554 19966 45556 20018
rect 45500 19964 45556 19966
rect 45612 19852 45668 19908
rect 44044 18620 44100 18676
rect 44156 18508 44212 18564
rect 44940 18844 44996 18900
rect 43708 17554 43764 17556
rect 43708 17502 43710 17554
rect 43710 17502 43762 17554
rect 43762 17502 43764 17554
rect 43708 17500 43764 17502
rect 43260 17388 43316 17444
rect 43596 17276 43652 17332
rect 43596 16604 43652 16660
rect 43036 14476 43092 14532
rect 43148 15260 43204 15316
rect 42588 13468 42644 13524
rect 42700 14252 42756 14308
rect 42700 13692 42756 13748
rect 43036 13580 43092 13636
rect 42812 13468 42868 13524
rect 42812 12236 42868 12292
rect 42700 12178 42756 12180
rect 42700 12126 42702 12178
rect 42702 12126 42754 12178
rect 42754 12126 42756 12178
rect 42700 12124 42756 12126
rect 42476 11788 42532 11844
rect 43036 12348 43092 12404
rect 42140 10556 42196 10612
rect 41580 9826 41636 9828
rect 41580 9774 41582 9826
rect 41582 9774 41634 9826
rect 41634 9774 41636 9826
rect 41580 9772 41636 9774
rect 41356 9714 41412 9716
rect 41356 9662 41358 9714
rect 41358 9662 41410 9714
rect 41410 9662 41412 9714
rect 41356 9660 41412 9662
rect 41468 9548 41524 9604
rect 41020 9042 41076 9044
rect 41020 8990 41022 9042
rect 41022 8990 41074 9042
rect 41074 8990 41076 9042
rect 41020 8988 41076 8990
rect 40012 8540 40068 8596
rect 39788 7420 39844 7476
rect 39788 7250 39844 7252
rect 39788 7198 39790 7250
rect 39790 7198 39842 7250
rect 39842 7198 39844 7250
rect 39788 7196 39844 7198
rect 40124 7250 40180 7252
rect 40124 7198 40126 7250
rect 40126 7198 40178 7250
rect 40178 7198 40180 7250
rect 40124 7196 40180 7198
rect 39676 6748 39732 6804
rect 41580 8876 41636 8932
rect 40236 6636 40292 6692
rect 39788 6130 39844 6132
rect 39788 6078 39790 6130
rect 39790 6078 39842 6130
rect 39842 6078 39844 6130
rect 39788 6076 39844 6078
rect 41356 8034 41412 8036
rect 41356 7982 41358 8034
rect 41358 7982 41410 8034
rect 41410 7982 41412 8034
rect 41356 7980 41412 7982
rect 41916 7532 41972 7588
rect 41244 7474 41300 7476
rect 41244 7422 41246 7474
rect 41246 7422 41298 7474
rect 41298 7422 41300 7474
rect 41244 7420 41300 7422
rect 41020 7196 41076 7252
rect 40460 6748 40516 6804
rect 40012 5852 40068 5908
rect 40124 5068 40180 5124
rect 40236 5516 40292 5572
rect 40236 4396 40292 4452
rect 39900 3724 39956 3780
rect 38668 3500 38724 3556
rect 40572 6636 40628 6692
rect 40572 6300 40628 6356
rect 41020 6524 41076 6580
rect 41916 7362 41972 7364
rect 41916 7310 41918 7362
rect 41918 7310 41970 7362
rect 41970 7310 41972 7362
rect 41916 7308 41972 7310
rect 41916 5906 41972 5908
rect 41916 5854 41918 5906
rect 41918 5854 41970 5906
rect 41970 5854 41972 5906
rect 41916 5852 41972 5854
rect 43260 14476 43316 14532
rect 43708 14700 43764 14756
rect 43596 14364 43652 14420
rect 43708 13746 43764 13748
rect 43708 13694 43710 13746
rect 43710 13694 43762 13746
rect 43762 13694 43764 13746
rect 43708 13692 43764 13694
rect 43260 12908 43316 12964
rect 43372 12290 43428 12292
rect 43372 12238 43374 12290
rect 43374 12238 43426 12290
rect 43426 12238 43428 12290
rect 43372 12236 43428 12238
rect 43260 12124 43316 12180
rect 43260 11394 43316 11396
rect 43260 11342 43262 11394
rect 43262 11342 43314 11394
rect 43314 11342 43316 11394
rect 43260 11340 43316 11342
rect 42252 9996 42308 10052
rect 42700 9826 42756 9828
rect 42700 9774 42702 9826
rect 42702 9774 42754 9826
rect 42754 9774 42756 9826
rect 42700 9772 42756 9774
rect 42476 9660 42532 9716
rect 42364 9266 42420 9268
rect 42364 9214 42366 9266
rect 42366 9214 42418 9266
rect 42418 9214 42420 9266
rect 42364 9212 42420 9214
rect 42364 9042 42420 9044
rect 42364 8990 42366 9042
rect 42366 8990 42418 9042
rect 42418 8990 42420 9042
rect 42364 8988 42420 8990
rect 42588 9602 42644 9604
rect 42588 9550 42590 9602
rect 42590 9550 42642 9602
rect 42642 9550 42644 9602
rect 42588 9548 42644 9550
rect 42140 7980 42196 8036
rect 42476 6860 42532 6916
rect 43484 10892 43540 10948
rect 43260 9884 43316 9940
rect 43148 9772 43204 9828
rect 43148 8540 43204 8596
rect 43596 10780 43652 10836
rect 43596 9996 43652 10052
rect 43596 9266 43652 9268
rect 43596 9214 43598 9266
rect 43598 9214 43650 9266
rect 43650 9214 43652 9266
rect 43596 9212 43652 9214
rect 43820 8988 43876 9044
rect 43708 8652 43764 8708
rect 42812 7980 42868 8036
rect 42924 7532 42980 7588
rect 42700 7308 42756 7364
rect 42700 6578 42756 6580
rect 42700 6526 42702 6578
rect 42702 6526 42754 6578
rect 42754 6526 42756 6578
rect 42700 6524 42756 6526
rect 42252 5180 42308 5236
rect 43036 5234 43092 5236
rect 43036 5182 43038 5234
rect 43038 5182 43090 5234
rect 43090 5182 43092 5234
rect 43036 5180 43092 5182
rect 42028 5010 42084 5012
rect 42028 4958 42030 5010
rect 42030 4958 42082 5010
rect 42082 4958 42084 5010
rect 42028 4956 42084 4958
rect 41356 4284 41412 4340
rect 42700 4284 42756 4340
rect 43372 7586 43428 7588
rect 43372 7534 43374 7586
rect 43374 7534 43426 7586
rect 43426 7534 43428 7586
rect 43372 7532 43428 7534
rect 43484 7420 43540 7476
rect 43260 6690 43316 6692
rect 43260 6638 43262 6690
rect 43262 6638 43314 6690
rect 43314 6638 43316 6690
rect 43260 6636 43316 6638
rect 43260 6466 43316 6468
rect 43260 6414 43262 6466
rect 43262 6414 43314 6466
rect 43314 6414 43316 6466
rect 43260 6412 43316 6414
rect 43596 6860 43652 6916
rect 43708 6076 43764 6132
rect 43372 4956 43428 5012
rect 43148 4284 43204 4340
rect 42700 3666 42756 3668
rect 42700 3614 42702 3666
rect 42702 3614 42754 3666
rect 42754 3614 42756 3666
rect 42700 3612 42756 3614
rect 44044 17442 44100 17444
rect 44044 17390 44046 17442
rect 44046 17390 44098 17442
rect 44098 17390 44100 17442
rect 44044 17388 44100 17390
rect 44268 16098 44324 16100
rect 44268 16046 44270 16098
rect 44270 16046 44322 16098
rect 44322 16046 44324 16098
rect 44268 16044 44324 16046
rect 44268 15484 44324 15540
rect 44044 15314 44100 15316
rect 44044 15262 44046 15314
rect 44046 15262 44098 15314
rect 44098 15262 44100 15314
rect 44044 15260 44100 15262
rect 44828 18396 44884 18452
rect 46396 24722 46452 24724
rect 46396 24670 46398 24722
rect 46398 24670 46450 24722
rect 46450 24670 46452 24722
rect 46396 24668 46452 24670
rect 46620 25228 46676 25284
rect 47292 27020 47348 27076
rect 47068 26460 47124 26516
rect 47068 25564 47124 25620
rect 47068 25340 47124 25396
rect 49308 33180 49364 33236
rect 49196 32786 49252 32788
rect 49196 32734 49198 32786
rect 49198 32734 49250 32786
rect 49250 32734 49252 32786
rect 49196 32732 49252 32734
rect 48748 31836 48804 31892
rect 49532 32620 49588 32676
rect 48300 28140 48356 28196
rect 48860 29372 48916 29428
rect 48748 29314 48804 29316
rect 48748 29262 48750 29314
rect 48750 29262 48802 29314
rect 48802 29262 48804 29314
rect 48748 29260 48804 29262
rect 48636 29036 48692 29092
rect 47516 27970 47572 27972
rect 47516 27918 47518 27970
rect 47518 27918 47570 27970
rect 47570 27918 47572 27970
rect 47516 27916 47572 27918
rect 47628 26178 47684 26180
rect 47628 26126 47630 26178
rect 47630 26126 47682 26178
rect 47682 26126 47684 26178
rect 47628 26124 47684 26126
rect 47740 25900 47796 25956
rect 47964 25452 48020 25508
rect 47628 24780 47684 24836
rect 46732 24108 46788 24164
rect 46732 23938 46788 23940
rect 46732 23886 46734 23938
rect 46734 23886 46786 23938
rect 46786 23886 46788 23938
rect 46732 23884 46788 23886
rect 46620 23436 46676 23492
rect 46396 23100 46452 23156
rect 45612 19292 45668 19348
rect 45500 19122 45556 19124
rect 45500 19070 45502 19122
rect 45502 19070 45554 19122
rect 45554 19070 45556 19122
rect 45500 19068 45556 19070
rect 45388 18396 45444 18452
rect 45612 18844 45668 18900
rect 45500 18284 45556 18340
rect 45276 17890 45332 17892
rect 45276 17838 45278 17890
rect 45278 17838 45330 17890
rect 45330 17838 45332 17890
rect 45276 17836 45332 17838
rect 44828 15874 44884 15876
rect 44828 15822 44830 15874
rect 44830 15822 44882 15874
rect 44882 15822 44884 15874
rect 44828 15820 44884 15822
rect 44492 13522 44548 13524
rect 44492 13470 44494 13522
rect 44494 13470 44546 13522
rect 44546 13470 44548 13522
rect 44492 13468 44548 13470
rect 44268 12850 44324 12852
rect 44268 12798 44270 12850
rect 44270 12798 44322 12850
rect 44322 12798 44324 12850
rect 44268 12796 44324 12798
rect 44268 12178 44324 12180
rect 44268 12126 44270 12178
rect 44270 12126 44322 12178
rect 44322 12126 44324 12178
rect 44268 12124 44324 12126
rect 44156 11228 44212 11284
rect 44940 14754 44996 14756
rect 44940 14702 44942 14754
rect 44942 14702 44994 14754
rect 44994 14702 44996 14754
rect 44940 14700 44996 14702
rect 44940 12850 44996 12852
rect 44940 12798 44942 12850
rect 44942 12798 44994 12850
rect 44994 12798 44996 12850
rect 44940 12796 44996 12798
rect 46060 19292 46116 19348
rect 46172 19180 46228 19236
rect 45948 18396 46004 18452
rect 45724 17724 45780 17780
rect 45724 17276 45780 17332
rect 45836 18060 45892 18116
rect 46620 22316 46676 22372
rect 46844 23660 46900 23716
rect 47404 23436 47460 23492
rect 47180 23266 47236 23268
rect 47180 23214 47182 23266
rect 47182 23214 47234 23266
rect 47234 23214 47236 23266
rect 47180 23212 47236 23214
rect 47516 23378 47572 23380
rect 47516 23326 47518 23378
rect 47518 23326 47570 23378
rect 47570 23326 47572 23378
rect 47516 23324 47572 23326
rect 46844 23154 46900 23156
rect 46844 23102 46846 23154
rect 46846 23102 46898 23154
rect 46898 23102 46900 23154
rect 46844 23100 46900 23102
rect 47068 22764 47124 22820
rect 47068 22204 47124 22260
rect 47964 24892 48020 24948
rect 48188 26460 48244 26516
rect 48860 28812 48916 28868
rect 48748 28476 48804 28532
rect 48972 29202 49028 29204
rect 48972 29150 48974 29202
rect 48974 29150 49026 29202
rect 49026 29150 49028 29202
rect 48972 29148 49028 29150
rect 48748 27020 48804 27076
rect 47852 23154 47908 23156
rect 47852 23102 47854 23154
rect 47854 23102 47906 23154
rect 47906 23102 47908 23154
rect 47852 23100 47908 23102
rect 47852 22540 47908 22596
rect 47964 23884 48020 23940
rect 47852 22204 47908 22260
rect 48748 26124 48804 26180
rect 48972 25452 49028 25508
rect 48636 25228 48692 25284
rect 48860 24610 48916 24612
rect 48860 24558 48862 24610
rect 48862 24558 48914 24610
rect 48914 24558 48916 24610
rect 48860 24556 48916 24558
rect 48860 23772 48916 23828
rect 48188 23042 48244 23044
rect 48188 22990 48190 23042
rect 48190 22990 48242 23042
rect 48242 22990 48244 23042
rect 48188 22988 48244 22990
rect 48524 22204 48580 22260
rect 47740 21868 47796 21924
rect 47964 21756 48020 21812
rect 47628 21586 47684 21588
rect 47628 21534 47630 21586
rect 47630 21534 47682 21586
rect 47682 21534 47684 21586
rect 47628 21532 47684 21534
rect 47068 20018 47124 20020
rect 47068 19966 47070 20018
rect 47070 19966 47122 20018
rect 47122 19966 47124 20018
rect 47068 19964 47124 19966
rect 46396 19292 46452 19348
rect 46284 18450 46340 18452
rect 46284 18398 46286 18450
rect 46286 18398 46338 18450
rect 46338 18398 46340 18450
rect 46284 18396 46340 18398
rect 45836 16940 45892 16996
rect 45500 15484 45556 15540
rect 45276 15090 45332 15092
rect 45276 15038 45278 15090
rect 45278 15038 45330 15090
rect 45330 15038 45332 15090
rect 45276 15036 45332 15038
rect 45276 13580 45332 13636
rect 44716 11228 44772 11284
rect 45276 12124 45332 12180
rect 46172 14418 46228 14420
rect 46172 14366 46174 14418
rect 46174 14366 46226 14418
rect 46226 14366 46228 14418
rect 46172 14364 46228 14366
rect 46060 13692 46116 13748
rect 46060 13356 46116 13412
rect 46508 18284 46564 18340
rect 46508 17836 46564 17892
rect 46844 19292 46900 19348
rect 47292 19964 47348 20020
rect 46844 19122 46900 19124
rect 46844 19070 46846 19122
rect 46846 19070 46898 19122
rect 46898 19070 46900 19122
rect 46844 19068 46900 19070
rect 47068 19010 47124 19012
rect 47068 18958 47070 19010
rect 47070 18958 47122 19010
rect 47122 18958 47124 19010
rect 47068 18956 47124 18958
rect 46956 18844 47012 18900
rect 46732 18508 46788 18564
rect 47628 20300 47684 20356
rect 47740 20076 47796 20132
rect 47852 21420 47908 21476
rect 48300 21644 48356 21700
rect 49084 22204 49140 22260
rect 48860 21644 48916 21700
rect 48972 21532 49028 21588
rect 48860 21474 48916 21476
rect 48860 21422 48862 21474
rect 48862 21422 48914 21474
rect 48914 21422 48916 21474
rect 48860 21420 48916 21422
rect 49084 21420 49140 21476
rect 48412 21308 48468 21364
rect 48748 20636 48804 20692
rect 47740 19234 47796 19236
rect 47740 19182 47742 19234
rect 47742 19182 47794 19234
rect 47794 19182 47796 19234
rect 47740 19180 47796 19182
rect 46508 16156 46564 16212
rect 47068 15372 47124 15428
rect 47180 14924 47236 14980
rect 46508 14364 46564 14420
rect 47068 14418 47124 14420
rect 47068 14366 47070 14418
rect 47070 14366 47122 14418
rect 47122 14366 47124 14418
rect 47068 14364 47124 14366
rect 46844 14252 46900 14308
rect 46732 13692 46788 13748
rect 45164 11282 45220 11284
rect 45164 11230 45166 11282
rect 45166 11230 45218 11282
rect 45218 11230 45220 11282
rect 45164 11228 45220 11230
rect 44604 10108 44660 10164
rect 44268 9826 44324 9828
rect 44268 9774 44270 9826
rect 44270 9774 44322 9826
rect 44322 9774 44324 9826
rect 44268 9772 44324 9774
rect 45948 10892 46004 10948
rect 46396 10780 46452 10836
rect 47068 13020 47124 13076
rect 46844 11506 46900 11508
rect 46844 11454 46846 11506
rect 46846 11454 46898 11506
rect 46898 11454 46900 11506
rect 46844 11452 46900 11454
rect 47404 16044 47460 16100
rect 47852 17666 47908 17668
rect 47852 17614 47854 17666
rect 47854 17614 47906 17666
rect 47906 17614 47908 17666
rect 47852 17612 47908 17614
rect 49084 20578 49140 20580
rect 49084 20526 49086 20578
rect 49086 20526 49138 20578
rect 49138 20526 49140 20578
rect 49084 20524 49140 20526
rect 48860 20130 48916 20132
rect 48860 20078 48862 20130
rect 48862 20078 48914 20130
rect 48914 20078 48916 20130
rect 48860 20076 48916 20078
rect 48748 19852 48804 19908
rect 48748 18508 48804 18564
rect 49980 39452 50036 39508
rect 49868 38834 49924 38836
rect 49868 38782 49870 38834
rect 49870 38782 49922 38834
rect 49922 38782 49924 38834
rect 49868 38780 49924 38782
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50764 43484 50820 43540
rect 51548 46002 51604 46004
rect 51548 45950 51550 46002
rect 51550 45950 51602 46002
rect 51602 45950 51604 46002
rect 51548 45948 51604 45950
rect 51884 46284 51940 46340
rect 51548 45388 51604 45444
rect 51324 43372 51380 43428
rect 51212 42978 51268 42980
rect 51212 42926 51214 42978
rect 51214 42926 51266 42978
rect 51266 42926 51268 42978
rect 51212 42924 51268 42926
rect 51996 45724 52052 45780
rect 51884 45666 51940 45668
rect 51884 45614 51886 45666
rect 51886 45614 51938 45666
rect 51938 45614 51940 45666
rect 51884 45612 51940 45614
rect 51548 42700 51604 42756
rect 51884 45388 51940 45444
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 51548 42140 51604 42196
rect 50540 41858 50596 41860
rect 50540 41806 50542 41858
rect 50542 41806 50594 41858
rect 50594 41806 50596 41858
rect 50540 41804 50596 41806
rect 50764 40962 50820 40964
rect 50764 40910 50766 40962
rect 50766 40910 50818 40962
rect 50818 40910 50820 40962
rect 50764 40908 50820 40910
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50428 40348 50484 40404
rect 50316 39676 50372 39732
rect 50428 39618 50484 39620
rect 50428 39566 50430 39618
rect 50430 39566 50482 39618
rect 50482 39566 50484 39618
rect 50428 39564 50484 39566
rect 50316 39452 50372 39508
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50428 39004 50484 39060
rect 50316 38892 50372 38948
rect 49868 37884 49924 37940
rect 49868 37660 49924 37716
rect 50316 37378 50372 37380
rect 50316 37326 50318 37378
rect 50318 37326 50370 37378
rect 50370 37326 50372 37378
rect 50316 37324 50372 37326
rect 50764 38668 50820 38724
rect 50764 38050 50820 38052
rect 50764 37998 50766 38050
rect 50766 37998 50818 38050
rect 50818 37998 50820 38050
rect 50764 37996 50820 37998
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50204 36988 50260 37044
rect 50204 36764 50260 36820
rect 50540 36652 50596 36708
rect 49868 35308 49924 35364
rect 49980 34860 50036 34916
rect 50092 33404 50148 33460
rect 50204 34076 50260 34132
rect 51436 39564 51492 39620
rect 51772 43484 51828 43540
rect 51996 43708 52052 43764
rect 51772 42812 51828 42868
rect 51660 41804 51716 41860
rect 52108 42700 52164 42756
rect 51996 42082 52052 42084
rect 51996 42030 51998 42082
rect 51998 42030 52050 42082
rect 52050 42030 52052 42082
rect 51996 42028 52052 42030
rect 51996 41804 52052 41860
rect 53228 47740 53284 47796
rect 52892 46844 52948 46900
rect 52668 46284 52724 46340
rect 53340 45836 53396 45892
rect 52668 44940 52724 44996
rect 53340 45500 53396 45556
rect 53228 45052 53284 45108
rect 53340 44604 53396 44660
rect 52892 43932 52948 43988
rect 53116 44492 53172 44548
rect 53676 50092 53732 50148
rect 53788 49756 53844 49812
rect 53900 52332 53956 52388
rect 55020 57090 55076 57092
rect 55020 57038 55022 57090
rect 55022 57038 55074 57090
rect 55074 57038 55076 57090
rect 55020 57036 55076 57038
rect 54796 56812 54852 56868
rect 54796 56252 54852 56308
rect 54908 56588 54964 56644
rect 56700 57820 56756 57876
rect 55916 57708 55972 57764
rect 55468 57538 55524 57540
rect 55468 57486 55470 57538
rect 55470 57486 55522 57538
rect 55522 57486 55524 57538
rect 55468 57484 55524 57486
rect 55468 56588 55524 56644
rect 55804 57036 55860 57092
rect 55692 56866 55748 56868
rect 55692 56814 55694 56866
rect 55694 56814 55746 56866
rect 55746 56814 55748 56866
rect 55692 56812 55748 56814
rect 55580 56194 55636 56196
rect 55580 56142 55582 56194
rect 55582 56142 55634 56194
rect 55634 56142 55636 56194
rect 55580 56140 55636 56142
rect 55132 55468 55188 55524
rect 55468 55356 55524 55412
rect 56364 57036 56420 57092
rect 55916 55132 55972 55188
rect 54684 54514 54740 54516
rect 54684 54462 54686 54514
rect 54686 54462 54738 54514
rect 54738 54462 54740 54514
rect 54684 54460 54740 54462
rect 54348 54290 54404 54292
rect 54348 54238 54350 54290
rect 54350 54238 54402 54290
rect 54402 54238 54404 54290
rect 54348 54236 54404 54238
rect 54348 52834 54404 52836
rect 54348 52782 54350 52834
rect 54350 52782 54402 52834
rect 54402 52782 54404 52834
rect 54348 52780 54404 52782
rect 54348 52556 54404 52612
rect 54460 52444 54516 52500
rect 53788 49532 53844 49588
rect 54124 50988 54180 51044
rect 54236 51996 54292 52052
rect 55132 53730 55188 53732
rect 55132 53678 55134 53730
rect 55134 53678 55186 53730
rect 55186 53678 55188 53730
rect 55132 53676 55188 53678
rect 55132 53116 55188 53172
rect 55020 53058 55076 53060
rect 55020 53006 55022 53058
rect 55022 53006 55074 53058
rect 55074 53006 55076 53058
rect 55020 53004 55076 53006
rect 54796 52444 54852 52500
rect 54572 51378 54628 51380
rect 54572 51326 54574 51378
rect 54574 51326 54626 51378
rect 54626 51326 54628 51378
rect 54572 51324 54628 51326
rect 55356 53004 55412 53060
rect 54908 49980 54964 50036
rect 56476 56642 56532 56644
rect 56476 56590 56478 56642
rect 56478 56590 56530 56642
rect 56530 56590 56532 56642
rect 56476 56588 56532 56590
rect 56028 54796 56084 54852
rect 56140 55468 56196 55524
rect 55692 54684 55748 54740
rect 55580 53116 55636 53172
rect 55580 52722 55636 52724
rect 55580 52670 55582 52722
rect 55582 52670 55634 52722
rect 55634 52670 55636 52722
rect 55580 52668 55636 52670
rect 55468 52556 55524 52612
rect 56812 56252 56868 56308
rect 56476 55468 56532 55524
rect 56924 56924 56980 56980
rect 57820 56978 57876 56980
rect 57820 56926 57822 56978
rect 57822 56926 57874 56978
rect 57874 56926 57876 56978
rect 57820 56924 57876 56926
rect 57036 56812 57092 56868
rect 57260 56700 57316 56756
rect 58268 56754 58324 56756
rect 58268 56702 58270 56754
rect 58270 56702 58322 56754
rect 58322 56702 58324 56754
rect 58268 56700 58324 56702
rect 59052 56700 59108 56756
rect 57820 56194 57876 56196
rect 57820 56142 57822 56194
rect 57822 56142 57874 56194
rect 57874 56142 57876 56194
rect 57820 56140 57876 56142
rect 57260 55580 57316 55636
rect 56812 55356 56868 55412
rect 56588 54684 56644 54740
rect 56588 54348 56644 54404
rect 56700 53676 56756 53732
rect 56252 53116 56308 53172
rect 55916 51548 55972 51604
rect 55692 50594 55748 50596
rect 55692 50542 55694 50594
rect 55694 50542 55746 50594
rect 55746 50542 55748 50594
rect 55692 50540 55748 50542
rect 55244 49980 55300 50036
rect 54236 49810 54292 49812
rect 54236 49758 54238 49810
rect 54238 49758 54290 49810
rect 54290 49758 54292 49810
rect 54236 49756 54292 49758
rect 55356 49644 55412 49700
rect 54572 49250 54628 49252
rect 54572 49198 54574 49250
rect 54574 49198 54626 49250
rect 54626 49198 54628 49250
rect 54572 49196 54628 49198
rect 53900 47180 53956 47236
rect 53676 46898 53732 46900
rect 53676 46846 53678 46898
rect 53678 46846 53730 46898
rect 53730 46846 53732 46898
rect 53676 46844 53732 46846
rect 53788 46508 53844 46564
rect 53564 45500 53620 45556
rect 54348 46396 54404 46452
rect 53676 45052 53732 45108
rect 52780 43708 52836 43764
rect 52892 43538 52948 43540
rect 52892 43486 52894 43538
rect 52894 43486 52946 43538
rect 52946 43486 52948 43538
rect 52892 43484 52948 43486
rect 52780 43036 52836 43092
rect 52892 42754 52948 42756
rect 52892 42702 52894 42754
rect 52894 42702 52946 42754
rect 52946 42702 52948 42754
rect 52892 42700 52948 42702
rect 53228 43820 53284 43876
rect 53564 43932 53620 43988
rect 53564 43260 53620 43316
rect 53452 42924 53508 42980
rect 53452 42700 53508 42756
rect 52332 42028 52388 42084
rect 52668 41916 52724 41972
rect 52332 41132 52388 41188
rect 51772 39340 51828 39396
rect 52108 39228 52164 39284
rect 51548 38780 51604 38836
rect 51212 38610 51268 38612
rect 51212 38558 51214 38610
rect 51214 38558 51266 38610
rect 51266 38558 51268 38610
rect 51212 38556 51268 38558
rect 51548 38556 51604 38612
rect 51100 37772 51156 37828
rect 51100 37266 51156 37268
rect 51100 37214 51102 37266
rect 51102 37214 51154 37266
rect 51154 37214 51156 37266
rect 51100 37212 51156 37214
rect 50876 36316 50932 36372
rect 50988 36764 51044 36820
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50428 35196 50484 35252
rect 50988 35532 51044 35588
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50428 34300 50484 34356
rect 51212 35196 51268 35252
rect 50988 33964 51044 34020
rect 50988 33068 51044 33124
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 49980 32060 50036 32116
rect 49756 29484 49812 29540
rect 49756 28924 49812 28980
rect 49868 28588 49924 28644
rect 49756 27298 49812 27300
rect 49756 27246 49758 27298
rect 49758 27246 49810 27298
rect 49810 27246 49812 27298
rect 49756 27244 49812 27246
rect 49756 26908 49812 26964
rect 49420 25506 49476 25508
rect 49420 25454 49422 25506
rect 49422 25454 49474 25506
rect 49474 25454 49476 25506
rect 49420 25452 49476 25454
rect 49308 25340 49364 25396
rect 50204 30044 50260 30100
rect 49980 27692 50036 27748
rect 50092 27916 50148 27972
rect 50204 27804 50260 27860
rect 50204 27468 50260 27524
rect 50316 27132 50372 27188
rect 50540 31948 50596 32004
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 51324 33292 51380 33348
rect 51212 32562 51268 32564
rect 51212 32510 51214 32562
rect 51214 32510 51266 32562
rect 51266 32510 51268 32562
rect 51212 32508 51268 32510
rect 51100 32060 51156 32116
rect 51548 36988 51604 37044
rect 51996 37996 52052 38052
rect 52108 38556 52164 38612
rect 52892 41186 52948 41188
rect 52892 41134 52894 41186
rect 52894 41134 52946 41186
rect 52946 41134 52948 41186
rect 52892 41132 52948 41134
rect 52444 38834 52500 38836
rect 52444 38782 52446 38834
rect 52446 38782 52498 38834
rect 52498 38782 52500 38834
rect 52444 38780 52500 38782
rect 53452 42194 53508 42196
rect 53452 42142 53454 42194
rect 53454 42142 53506 42194
rect 53506 42142 53508 42194
rect 53452 42140 53508 42142
rect 53228 41692 53284 41748
rect 53116 40962 53172 40964
rect 53116 40910 53118 40962
rect 53118 40910 53170 40962
rect 53170 40910 53172 40962
rect 53116 40908 53172 40910
rect 53228 40460 53284 40516
rect 54796 47628 54852 47684
rect 55692 49196 55748 49252
rect 55804 49420 55860 49476
rect 55468 48972 55524 49028
rect 54908 47404 54964 47460
rect 55020 48076 55076 48132
rect 55468 47740 55524 47796
rect 55244 47068 55300 47124
rect 55356 47628 55412 47684
rect 54796 46508 54852 46564
rect 55020 46396 55076 46452
rect 54684 45724 54740 45780
rect 54012 44380 54068 44436
rect 54572 44716 54628 44772
rect 54684 45052 54740 45108
rect 54460 44546 54516 44548
rect 54460 44494 54462 44546
rect 54462 44494 54514 44546
rect 54514 44494 54516 44546
rect 54460 44492 54516 44494
rect 53900 44044 53956 44100
rect 54012 44156 54068 44212
rect 53788 43932 53844 43988
rect 54012 43596 54068 43652
rect 53900 43260 53956 43316
rect 53900 43036 53956 43092
rect 53228 40012 53284 40068
rect 53564 39730 53620 39732
rect 53564 39678 53566 39730
rect 53566 39678 53618 39730
rect 53618 39678 53620 39730
rect 53564 39676 53620 39678
rect 53116 39004 53172 39060
rect 53004 38780 53060 38836
rect 52332 37884 52388 37940
rect 51884 37324 51940 37380
rect 52556 37266 52612 37268
rect 52556 37214 52558 37266
rect 52558 37214 52610 37266
rect 52610 37214 52612 37266
rect 52556 37212 52612 37214
rect 52892 36988 52948 37044
rect 53340 38668 53396 38724
rect 52220 36540 52276 36596
rect 52892 36540 52948 36596
rect 51884 36428 51940 36484
rect 52780 36482 52836 36484
rect 52780 36430 52782 36482
rect 52782 36430 52834 36482
rect 52834 36430 52836 36482
rect 52780 36428 52836 36430
rect 51772 36316 51828 36372
rect 52220 36204 52276 36260
rect 51772 35026 51828 35028
rect 51772 34974 51774 35026
rect 51774 34974 51826 35026
rect 51826 34974 51828 35026
rect 51772 34972 51828 34974
rect 51996 35698 52052 35700
rect 51996 35646 51998 35698
rect 51998 35646 52050 35698
rect 52050 35646 52052 35698
rect 51996 35644 52052 35646
rect 52668 35868 52724 35924
rect 51660 33964 51716 34020
rect 51996 33964 52052 34020
rect 51548 33346 51604 33348
rect 51548 33294 51550 33346
rect 51550 33294 51602 33346
rect 51602 33294 51604 33346
rect 51548 33292 51604 33294
rect 52108 33628 52164 33684
rect 51436 31164 51492 31220
rect 51996 32396 52052 32452
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50540 29372 50596 29428
rect 50540 28812 50596 28868
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50764 27804 50820 27860
rect 50540 27186 50596 27188
rect 50540 27134 50542 27186
rect 50542 27134 50594 27186
rect 50594 27134 50596 27186
rect 50540 27132 50596 27134
rect 51212 29484 51268 29540
rect 50988 28642 51044 28644
rect 50988 28590 50990 28642
rect 50990 28590 51042 28642
rect 51042 28590 51044 28642
rect 50988 28588 51044 28590
rect 51660 31948 51716 32004
rect 50876 27356 50932 27412
rect 50988 27074 51044 27076
rect 50988 27022 50990 27074
rect 50990 27022 51042 27074
rect 51042 27022 51044 27074
rect 50988 27020 51044 27022
rect 50092 26908 50148 26964
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50092 26402 50148 26404
rect 50092 26350 50094 26402
rect 50094 26350 50146 26402
rect 50146 26350 50148 26402
rect 50092 26348 50148 26350
rect 49644 26290 49700 26292
rect 49644 26238 49646 26290
rect 49646 26238 49698 26290
rect 49698 26238 49700 26290
rect 49644 26236 49700 26238
rect 49868 25788 49924 25844
rect 50540 25788 50596 25844
rect 50988 25676 51044 25732
rect 50092 25452 50148 25508
rect 49756 25282 49812 25284
rect 49756 25230 49758 25282
rect 49758 25230 49810 25282
rect 49810 25230 49812 25282
rect 49756 25228 49812 25230
rect 49868 24780 49924 24836
rect 50540 25394 50596 25396
rect 50540 25342 50542 25394
rect 50542 25342 50594 25394
rect 50594 25342 50596 25394
rect 50540 25340 50596 25342
rect 50876 25506 50932 25508
rect 50876 25454 50878 25506
rect 50878 25454 50930 25506
rect 50930 25454 50932 25506
rect 50876 25452 50932 25454
rect 50204 25004 50260 25060
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50092 24780 50148 24836
rect 50540 24892 50596 24948
rect 49532 24722 49588 24724
rect 49532 24670 49534 24722
rect 49534 24670 49586 24722
rect 49586 24670 49588 24722
rect 49532 24668 49588 24670
rect 49756 24722 49812 24724
rect 49756 24670 49758 24722
rect 49758 24670 49810 24722
rect 49810 24670 49812 24722
rect 49756 24668 49812 24670
rect 49420 23772 49476 23828
rect 49308 22204 49364 22260
rect 49420 21644 49476 21700
rect 49644 23996 49700 24052
rect 49644 23772 49700 23828
rect 49868 23154 49924 23156
rect 49868 23102 49870 23154
rect 49870 23102 49922 23154
rect 49922 23102 49924 23154
rect 49868 23100 49924 23102
rect 49980 22594 50036 22596
rect 49980 22542 49982 22594
rect 49982 22542 50034 22594
rect 50034 22542 50036 22594
rect 49980 22540 50036 22542
rect 49532 21532 49588 21588
rect 49644 21644 49700 21700
rect 49308 21308 49364 21364
rect 49644 21196 49700 21252
rect 49532 20914 49588 20916
rect 49532 20862 49534 20914
rect 49534 20862 49586 20914
rect 49586 20862 49588 20914
rect 49532 20860 49588 20862
rect 49308 20018 49364 20020
rect 49308 19966 49310 20018
rect 49310 19966 49362 20018
rect 49362 19966 49364 20018
rect 49308 19964 49364 19966
rect 49084 19180 49140 19236
rect 48860 18396 48916 18452
rect 48636 17836 48692 17892
rect 49084 17666 49140 17668
rect 49084 17614 49086 17666
rect 49086 17614 49138 17666
rect 49138 17614 49140 17666
rect 49084 17612 49140 17614
rect 49420 18844 49476 18900
rect 49644 18620 49700 18676
rect 49980 21474 50036 21476
rect 49980 21422 49982 21474
rect 49982 21422 50034 21474
rect 50034 21422 50036 21474
rect 49980 21420 50036 21422
rect 50540 24498 50596 24500
rect 50540 24446 50542 24498
rect 50542 24446 50594 24498
rect 50594 24446 50596 24498
rect 50540 24444 50596 24446
rect 50988 24444 51044 24500
rect 50540 24108 50596 24164
rect 50652 24220 50708 24276
rect 51100 23938 51156 23940
rect 51100 23886 51102 23938
rect 51102 23886 51154 23938
rect 51154 23886 51156 23938
rect 51100 23884 51156 23886
rect 50876 23826 50932 23828
rect 50876 23774 50878 23826
rect 50878 23774 50930 23826
rect 50930 23774 50932 23826
rect 50876 23772 50932 23774
rect 50092 21084 50148 21140
rect 50428 23660 50484 23716
rect 49868 20860 49924 20916
rect 50204 20636 50260 20692
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50540 23100 50596 23156
rect 51100 22316 51156 22372
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 52332 35420 52388 35476
rect 52220 32732 52276 32788
rect 52220 31948 52276 32004
rect 51772 30940 51828 30996
rect 51884 30210 51940 30212
rect 51884 30158 51886 30210
rect 51886 30158 51938 30210
rect 51938 30158 51940 30210
rect 51884 30156 51940 30158
rect 52108 29372 52164 29428
rect 51996 29314 52052 29316
rect 51996 29262 51998 29314
rect 51998 29262 52050 29314
rect 52050 29262 52052 29314
rect 51996 29260 52052 29262
rect 52780 35532 52836 35588
rect 53340 36876 53396 36932
rect 53228 36764 53284 36820
rect 53116 36482 53172 36484
rect 53116 36430 53118 36482
rect 53118 36430 53170 36482
rect 53170 36430 53172 36482
rect 53116 36428 53172 36430
rect 53228 36204 53284 36260
rect 53004 35868 53060 35924
rect 53116 36092 53172 36148
rect 52892 35644 52948 35700
rect 53340 35644 53396 35700
rect 53004 35138 53060 35140
rect 53004 35086 53006 35138
rect 53006 35086 53058 35138
rect 53058 35086 53060 35138
rect 53004 35084 53060 35086
rect 53788 42924 53844 42980
rect 54236 43820 54292 43876
rect 54348 43762 54404 43764
rect 54348 43710 54350 43762
rect 54350 43710 54402 43762
rect 54402 43710 54404 43762
rect 54348 43708 54404 43710
rect 54236 42140 54292 42196
rect 54572 42812 54628 42868
rect 55132 45052 55188 45108
rect 55244 46396 55300 46452
rect 55468 47458 55524 47460
rect 55468 47406 55470 47458
rect 55470 47406 55522 47458
rect 55522 47406 55524 47458
rect 55468 47404 55524 47406
rect 55580 46732 55636 46788
rect 56028 47740 56084 47796
rect 56924 55020 56980 55076
rect 56924 53788 56980 53844
rect 56588 52834 56644 52836
rect 56588 52782 56590 52834
rect 56590 52782 56642 52834
rect 56642 52782 56644 52834
rect 56588 52780 56644 52782
rect 57148 52722 57204 52724
rect 57148 52670 57150 52722
rect 57150 52670 57202 52722
rect 57202 52670 57204 52722
rect 57148 52668 57204 52670
rect 57036 51436 57092 51492
rect 57036 50876 57092 50932
rect 58156 55298 58212 55300
rect 58156 55246 58158 55298
rect 58158 55246 58210 55298
rect 58210 55246 58212 55298
rect 58156 55244 58212 55246
rect 58380 56306 58436 56308
rect 58380 56254 58382 56306
rect 58382 56254 58434 56306
rect 58434 56254 58436 56306
rect 58380 56252 58436 56254
rect 57596 54796 57652 54852
rect 57484 53058 57540 53060
rect 57484 53006 57486 53058
rect 57486 53006 57538 53058
rect 57538 53006 57540 53058
rect 57484 53004 57540 53006
rect 58716 55186 58772 55188
rect 58716 55134 58718 55186
rect 58718 55134 58770 55186
rect 58770 55134 58772 55186
rect 58716 55132 58772 55134
rect 57708 53954 57764 53956
rect 57708 53902 57710 53954
rect 57710 53902 57762 53954
rect 57762 53902 57764 53954
rect 57708 53900 57764 53902
rect 57932 53452 57988 53508
rect 58044 53730 58100 53732
rect 58044 53678 58046 53730
rect 58046 53678 58098 53730
rect 58098 53678 58100 53730
rect 58044 53676 58100 53678
rect 58492 53676 58548 53732
rect 59276 56306 59332 56308
rect 59276 56254 59278 56306
rect 59278 56254 59330 56306
rect 59330 56254 59332 56306
rect 59276 56252 59332 56254
rect 62748 55244 62804 55300
rect 59388 55132 59444 55188
rect 58940 53788 58996 53844
rect 59052 53730 59108 53732
rect 59052 53678 59054 53730
rect 59054 53678 59106 53730
rect 59106 53678 59108 53730
rect 59052 53676 59108 53678
rect 59612 53506 59668 53508
rect 59612 53454 59614 53506
rect 59614 53454 59666 53506
rect 59666 53454 59668 53506
rect 59612 53452 59668 53454
rect 57260 50764 57316 50820
rect 57484 51436 57540 51492
rect 57036 50652 57092 50708
rect 56700 50204 56756 50260
rect 56588 50034 56644 50036
rect 56588 49982 56590 50034
rect 56590 49982 56642 50034
rect 56642 49982 56644 50034
rect 56588 49980 56644 49982
rect 56700 48860 56756 48916
rect 56924 50482 56980 50484
rect 56924 50430 56926 50482
rect 56926 50430 56978 50482
rect 56978 50430 56980 50482
rect 56924 50428 56980 50430
rect 56924 49810 56980 49812
rect 56924 49758 56926 49810
rect 56926 49758 56978 49810
rect 56978 49758 56980 49810
rect 56924 49756 56980 49758
rect 56364 48748 56420 48804
rect 57820 51266 57876 51268
rect 57820 51214 57822 51266
rect 57822 51214 57874 51266
rect 57874 51214 57876 51266
rect 57820 51212 57876 51214
rect 57708 51100 57764 51156
rect 57932 51100 57988 51156
rect 57484 50092 57540 50148
rect 57148 49868 57204 49924
rect 57148 49084 57204 49140
rect 57036 48636 57092 48692
rect 56700 48466 56756 48468
rect 56700 48414 56702 48466
rect 56702 48414 56754 48466
rect 56754 48414 56756 48466
rect 56700 48412 56756 48414
rect 57036 48300 57092 48356
rect 56924 47852 56980 47908
rect 56252 47068 56308 47124
rect 55580 46172 55636 46228
rect 54908 44268 54964 44324
rect 54796 43820 54852 43876
rect 55356 43932 55412 43988
rect 55020 43538 55076 43540
rect 55020 43486 55022 43538
rect 55022 43486 55074 43538
rect 55074 43486 55076 43538
rect 55020 43484 55076 43486
rect 55356 41804 55412 41860
rect 54572 41132 54628 41188
rect 55132 40796 55188 40852
rect 54572 40684 54628 40740
rect 54236 40514 54292 40516
rect 54236 40462 54238 40514
rect 54238 40462 54290 40514
rect 54290 40462 54292 40514
rect 54236 40460 54292 40462
rect 53788 40236 53844 40292
rect 54348 40124 54404 40180
rect 53788 38780 53844 38836
rect 53900 37938 53956 37940
rect 53900 37886 53902 37938
rect 53902 37886 53954 37938
rect 53954 37886 53956 37938
rect 53900 37884 53956 37886
rect 54012 37490 54068 37492
rect 54012 37438 54014 37490
rect 54014 37438 54066 37490
rect 54066 37438 54068 37490
rect 54012 37436 54068 37438
rect 54236 37266 54292 37268
rect 54236 37214 54238 37266
rect 54238 37214 54290 37266
rect 54290 37214 54292 37266
rect 54236 37212 54292 37214
rect 54124 37154 54180 37156
rect 54124 37102 54126 37154
rect 54126 37102 54178 37154
rect 54178 37102 54180 37154
rect 54124 37100 54180 37102
rect 54012 36988 54068 37044
rect 53788 36764 53844 36820
rect 53564 36092 53620 36148
rect 53564 35138 53620 35140
rect 53564 35086 53566 35138
rect 53566 35086 53618 35138
rect 53618 35086 53620 35138
rect 53564 35084 53620 35086
rect 53452 34972 53508 35028
rect 53788 35196 53844 35252
rect 53676 34860 53732 34916
rect 54012 36482 54068 36484
rect 54012 36430 54014 36482
rect 54014 36430 54066 36482
rect 54066 36430 54068 36482
rect 54012 36428 54068 36430
rect 54012 35586 54068 35588
rect 54012 35534 54014 35586
rect 54014 35534 54066 35586
rect 54066 35534 54068 35586
rect 54012 35532 54068 35534
rect 54684 40348 54740 40404
rect 54796 39900 54852 39956
rect 55132 40124 55188 40180
rect 54796 38556 54852 38612
rect 54908 37996 54964 38052
rect 55020 37884 55076 37940
rect 55356 41244 55412 41300
rect 55916 45218 55972 45220
rect 55916 45166 55918 45218
rect 55918 45166 55970 45218
rect 55970 45166 55972 45218
rect 55916 45164 55972 45166
rect 55580 44940 55636 44996
rect 55916 44994 55972 44996
rect 55916 44942 55918 44994
rect 55918 44942 55970 44994
rect 55970 44942 55972 44994
rect 55916 44940 55972 44942
rect 55916 44380 55972 44436
rect 55580 44044 55636 44100
rect 55468 40908 55524 40964
rect 55804 43650 55860 43652
rect 55804 43598 55806 43650
rect 55806 43598 55858 43650
rect 55858 43598 55860 43650
rect 55804 43596 55860 43598
rect 55916 43036 55972 43092
rect 56700 47292 56756 47348
rect 56588 44604 56644 44660
rect 56476 44380 56532 44436
rect 56252 44156 56308 44212
rect 58044 50594 58100 50596
rect 58044 50542 58046 50594
rect 58046 50542 58098 50594
rect 58098 50542 58100 50594
rect 58044 50540 58100 50542
rect 57932 49644 57988 49700
rect 57820 49532 57876 49588
rect 58044 49308 58100 49364
rect 57484 49196 57540 49252
rect 57260 46732 57316 46788
rect 57820 48300 57876 48356
rect 57596 46732 57652 46788
rect 57932 48242 57988 48244
rect 57932 48190 57934 48242
rect 57934 48190 57986 48242
rect 57986 48190 57988 48242
rect 57932 48188 57988 48190
rect 57708 47068 57764 47124
rect 57260 46396 57316 46452
rect 56924 45276 56980 45332
rect 57036 44268 57092 44324
rect 56812 44210 56868 44212
rect 56812 44158 56814 44210
rect 56814 44158 56866 44210
rect 56866 44158 56868 44210
rect 56812 44156 56868 44158
rect 56700 43820 56756 43876
rect 56028 42812 56084 42868
rect 55916 42754 55972 42756
rect 55916 42702 55918 42754
rect 55918 42702 55970 42754
rect 55970 42702 55972 42754
rect 55916 42700 55972 42702
rect 55692 40684 55748 40740
rect 55804 41356 55860 41412
rect 55580 39900 55636 39956
rect 55916 41244 55972 41300
rect 55916 41074 55972 41076
rect 55916 41022 55918 41074
rect 55918 41022 55970 41074
rect 55970 41022 55972 41074
rect 55916 41020 55972 41022
rect 55804 40514 55860 40516
rect 55804 40462 55806 40514
rect 55806 40462 55858 40514
rect 55858 40462 55860 40514
rect 55804 40460 55860 40462
rect 56028 40236 56084 40292
rect 55916 39900 55972 39956
rect 55356 39564 55412 39620
rect 55580 39452 55636 39508
rect 54908 36652 54964 36708
rect 54348 35644 54404 35700
rect 54796 36370 54852 36372
rect 54796 36318 54798 36370
rect 54798 36318 54850 36370
rect 54850 36318 54852 36370
rect 54796 36316 54852 36318
rect 54460 35420 54516 35476
rect 54796 35308 54852 35364
rect 55916 38834 55972 38836
rect 55916 38782 55918 38834
rect 55918 38782 55970 38834
rect 55970 38782 55972 38834
rect 55916 38780 55972 38782
rect 55804 38274 55860 38276
rect 55804 38222 55806 38274
rect 55806 38222 55858 38274
rect 55858 38222 55860 38274
rect 55804 38220 55860 38222
rect 55916 38050 55972 38052
rect 55916 37998 55918 38050
rect 55918 37998 55970 38050
rect 55970 37998 55972 38050
rect 55916 37996 55972 37998
rect 56364 42978 56420 42980
rect 56364 42926 56366 42978
rect 56366 42926 56418 42978
rect 56418 42926 56420 42978
rect 56364 42924 56420 42926
rect 56476 42866 56532 42868
rect 56476 42814 56478 42866
rect 56478 42814 56530 42866
rect 56530 42814 56532 42866
rect 56476 42812 56532 42814
rect 56252 41804 56308 41860
rect 56476 41410 56532 41412
rect 56476 41358 56478 41410
rect 56478 41358 56530 41410
rect 56530 41358 56532 41410
rect 56476 41356 56532 41358
rect 56588 40908 56644 40964
rect 56812 41356 56868 41412
rect 56364 40348 56420 40404
rect 56700 40460 56756 40516
rect 56364 39788 56420 39844
rect 55132 36652 55188 36708
rect 54572 34860 54628 34916
rect 54348 34524 54404 34580
rect 53788 34130 53844 34132
rect 53788 34078 53790 34130
rect 53790 34078 53842 34130
rect 53842 34078 53844 34130
rect 53788 34076 53844 34078
rect 54012 34130 54068 34132
rect 54012 34078 54014 34130
rect 54014 34078 54066 34130
rect 54066 34078 54068 34130
rect 54012 34076 54068 34078
rect 53228 33628 53284 33684
rect 53900 34018 53956 34020
rect 53900 33966 53902 34018
rect 53902 33966 53954 34018
rect 53954 33966 53956 34018
rect 53900 33964 53956 33966
rect 54236 33516 54292 33572
rect 52892 33292 52948 33348
rect 53340 33346 53396 33348
rect 53340 33294 53342 33346
rect 53342 33294 53394 33346
rect 53394 33294 53396 33346
rect 53340 33292 53396 33294
rect 53900 33346 53956 33348
rect 53900 33294 53902 33346
rect 53902 33294 53954 33346
rect 53954 33294 53956 33346
rect 53900 33292 53956 33294
rect 54684 33292 54740 33348
rect 52780 33180 52836 33236
rect 52780 32396 52836 32452
rect 52668 31836 52724 31892
rect 53004 32060 53060 32116
rect 53564 31948 53620 32004
rect 53676 32396 53732 32452
rect 53340 31836 53396 31892
rect 54124 32450 54180 32452
rect 54124 32398 54126 32450
rect 54126 32398 54178 32450
rect 54178 32398 54180 32450
rect 54124 32396 54180 32398
rect 54572 31836 54628 31892
rect 54460 31554 54516 31556
rect 54460 31502 54462 31554
rect 54462 31502 54514 31554
rect 54514 31502 54516 31554
rect 54460 31500 54516 31502
rect 52668 31276 52724 31332
rect 52332 29538 52388 29540
rect 52332 29486 52334 29538
rect 52334 29486 52386 29538
rect 52386 29486 52388 29538
rect 52332 29484 52388 29486
rect 51772 28700 51828 28756
rect 52108 28700 52164 28756
rect 52108 28252 52164 28308
rect 51996 28140 52052 28196
rect 51996 27858 52052 27860
rect 51996 27806 51998 27858
rect 51998 27806 52050 27858
rect 52050 27806 52052 27858
rect 51996 27804 52052 27806
rect 51324 27746 51380 27748
rect 51324 27694 51326 27746
rect 51326 27694 51378 27746
rect 51378 27694 51380 27746
rect 51324 27692 51380 27694
rect 51436 27580 51492 27636
rect 51660 27244 51716 27300
rect 52220 27580 52276 27636
rect 51884 26796 51940 26852
rect 51324 25340 51380 25396
rect 51436 24892 51492 24948
rect 52220 26012 52276 26068
rect 51548 24220 51604 24276
rect 51436 23996 51492 24052
rect 51324 23714 51380 23716
rect 51324 23662 51326 23714
rect 51326 23662 51378 23714
rect 51378 23662 51380 23714
rect 51324 23660 51380 23662
rect 51548 23154 51604 23156
rect 51548 23102 51550 23154
rect 51550 23102 51602 23154
rect 51602 23102 51604 23154
rect 51548 23100 51604 23102
rect 51660 22876 51716 22932
rect 51212 20860 51268 20916
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 51548 22258 51604 22260
rect 51548 22206 51550 22258
rect 51550 22206 51602 22258
rect 51602 22206 51604 22258
rect 51548 22204 51604 22206
rect 51436 21308 51492 21364
rect 51548 21868 51604 21924
rect 51436 20524 51492 20580
rect 50876 20076 50932 20132
rect 50988 20412 51044 20468
rect 51884 24556 51940 24612
rect 51996 24722 52052 24724
rect 51996 24670 51998 24722
rect 51998 24670 52050 24722
rect 52050 24670 52052 24722
rect 51996 24668 52052 24670
rect 51996 23772 52052 23828
rect 51996 23324 52052 23380
rect 51884 21980 51940 22036
rect 51996 22652 52052 22708
rect 52108 22316 52164 22372
rect 52108 22146 52164 22148
rect 52108 22094 52110 22146
rect 52110 22094 52162 22146
rect 52162 22094 52164 22146
rect 52108 22092 52164 22094
rect 51772 20188 51828 20244
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 49308 17500 49364 17556
rect 49532 17554 49588 17556
rect 49532 17502 49534 17554
rect 49534 17502 49586 17554
rect 49586 17502 49588 17554
rect 49532 17500 49588 17502
rect 50092 18338 50148 18340
rect 50092 18286 50094 18338
rect 50094 18286 50146 18338
rect 50146 18286 50148 18338
rect 50092 18284 50148 18286
rect 50204 17836 50260 17892
rect 49196 17388 49252 17444
rect 49980 17276 50036 17332
rect 48860 17052 48916 17108
rect 48748 16940 48804 16996
rect 47740 16716 47796 16772
rect 47628 16044 47684 16100
rect 47404 15036 47460 15092
rect 47516 14252 47572 14308
rect 48188 16098 48244 16100
rect 48188 16046 48190 16098
rect 48190 16046 48242 16098
rect 48242 16046 48244 16098
rect 48188 16044 48244 16046
rect 47852 15986 47908 15988
rect 47852 15934 47854 15986
rect 47854 15934 47906 15986
rect 47906 15934 47908 15986
rect 47852 15932 47908 15934
rect 47516 13916 47572 13972
rect 47964 15820 48020 15876
rect 47852 15426 47908 15428
rect 47852 15374 47854 15426
rect 47854 15374 47906 15426
rect 47906 15374 47908 15426
rect 47852 15372 47908 15374
rect 47740 14252 47796 14308
rect 47964 14812 48020 14868
rect 48188 15036 48244 15092
rect 48076 13804 48132 13860
rect 48636 16716 48692 16772
rect 48972 17164 49028 17220
rect 50988 18620 51044 18676
rect 52220 20130 52276 20132
rect 52220 20078 52222 20130
rect 52222 20078 52274 20130
rect 52274 20078 52276 20130
rect 52220 20076 52276 20078
rect 52108 19964 52164 20020
rect 50204 17052 50260 17108
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50428 16940 50484 16996
rect 49756 16716 49812 16772
rect 49084 16322 49140 16324
rect 49084 16270 49086 16322
rect 49086 16270 49138 16322
rect 49138 16270 49140 16322
rect 49084 16268 49140 16270
rect 48972 16156 49028 16212
rect 48636 15820 48692 15876
rect 49308 15596 49364 15652
rect 48748 15372 48804 15428
rect 48524 15148 48580 15204
rect 48860 15314 48916 15316
rect 48860 15262 48862 15314
rect 48862 15262 48914 15314
rect 48914 15262 48916 15314
rect 48860 15260 48916 15262
rect 49084 13916 49140 13972
rect 47628 13692 47684 13748
rect 49532 16268 49588 16324
rect 50204 16322 50260 16324
rect 50204 16270 50206 16322
rect 50206 16270 50258 16322
rect 50258 16270 50260 16322
rect 50204 16268 50260 16270
rect 49868 16210 49924 16212
rect 49868 16158 49870 16210
rect 49870 16158 49922 16210
rect 49922 16158 49924 16210
rect 49868 16156 49924 16158
rect 50876 15986 50932 15988
rect 50876 15934 50878 15986
rect 50878 15934 50930 15986
rect 50930 15934 50932 15986
rect 50876 15932 50932 15934
rect 50092 15596 50148 15652
rect 50092 15426 50148 15428
rect 50092 15374 50094 15426
rect 50094 15374 50146 15426
rect 50146 15374 50148 15426
rect 50092 15372 50148 15374
rect 49756 15260 49812 15316
rect 49868 15148 49924 15204
rect 49532 15036 49588 15092
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 51660 19516 51716 19572
rect 52780 31052 52836 31108
rect 52444 28140 52500 28196
rect 52668 30156 52724 30212
rect 53564 31106 53620 31108
rect 53564 31054 53566 31106
rect 53566 31054 53618 31106
rect 53618 31054 53620 31106
rect 53564 31052 53620 31054
rect 53228 30156 53284 30212
rect 53340 30098 53396 30100
rect 53340 30046 53342 30098
rect 53342 30046 53394 30098
rect 53394 30046 53396 30098
rect 53340 30044 53396 30046
rect 53004 28140 53060 28196
rect 52668 27970 52724 27972
rect 52668 27918 52670 27970
rect 52670 27918 52722 27970
rect 52722 27918 52724 27970
rect 52668 27916 52724 27918
rect 52556 27020 52612 27076
rect 52892 27746 52948 27748
rect 52892 27694 52894 27746
rect 52894 27694 52946 27746
rect 52946 27694 52948 27746
rect 52892 27692 52948 27694
rect 53676 28812 53732 28868
rect 52780 26850 52836 26852
rect 52780 26798 52782 26850
rect 52782 26798 52834 26850
rect 52834 26798 52836 26850
rect 52780 26796 52836 26798
rect 53340 28252 53396 28308
rect 53676 28140 53732 28196
rect 53564 27916 53620 27972
rect 53900 28140 53956 28196
rect 54124 30156 54180 30212
rect 54572 31052 54628 31108
rect 54460 30210 54516 30212
rect 54460 30158 54462 30210
rect 54462 30158 54514 30210
rect 54514 30158 54516 30210
rect 54460 30156 54516 30158
rect 54236 30044 54292 30100
rect 54348 28588 54404 28644
rect 54572 29426 54628 29428
rect 54572 29374 54574 29426
rect 54574 29374 54626 29426
rect 54626 29374 54628 29426
rect 54572 29372 54628 29374
rect 55244 35308 55300 35364
rect 54908 34972 54964 35028
rect 56028 36594 56084 36596
rect 56028 36542 56030 36594
rect 56030 36542 56082 36594
rect 56082 36542 56084 36594
rect 56028 36540 56084 36542
rect 55692 35474 55748 35476
rect 55692 35422 55694 35474
rect 55694 35422 55746 35474
rect 55746 35422 55748 35474
rect 55692 35420 55748 35422
rect 55468 35196 55524 35252
rect 55580 35138 55636 35140
rect 55580 35086 55582 35138
rect 55582 35086 55634 35138
rect 55634 35086 55636 35138
rect 55580 35084 55636 35086
rect 55804 35196 55860 35252
rect 55916 35308 55972 35364
rect 55692 34972 55748 35028
rect 55020 33628 55076 33684
rect 54908 33516 54964 33572
rect 55020 31500 55076 31556
rect 55020 30882 55076 30884
rect 55020 30830 55022 30882
rect 55022 30830 55074 30882
rect 55074 30830 55076 30882
rect 55020 30828 55076 30830
rect 55132 30156 55188 30212
rect 55020 29986 55076 29988
rect 55020 29934 55022 29986
rect 55022 29934 55074 29986
rect 55074 29934 55076 29986
rect 55020 29932 55076 29934
rect 54908 29314 54964 29316
rect 54908 29262 54910 29314
rect 54910 29262 54962 29314
rect 54962 29262 54964 29314
rect 54908 29260 54964 29262
rect 55692 33516 55748 33572
rect 55468 33458 55524 33460
rect 55468 33406 55470 33458
rect 55470 33406 55522 33458
rect 55522 33406 55524 33458
rect 55468 33404 55524 33406
rect 56028 34860 56084 34916
rect 57036 42812 57092 42868
rect 57036 42364 57092 42420
rect 56924 40572 56980 40628
rect 57036 41020 57092 41076
rect 57036 40460 57092 40516
rect 56700 38668 56756 38724
rect 57260 43484 57316 43540
rect 58156 49196 58212 49252
rect 58828 52162 58884 52164
rect 58828 52110 58830 52162
rect 58830 52110 58882 52162
rect 58882 52110 58884 52162
rect 58828 52108 58884 52110
rect 58380 51436 58436 51492
rect 58828 51324 58884 51380
rect 58716 50988 58772 51044
rect 58492 50482 58548 50484
rect 58492 50430 58494 50482
rect 58494 50430 58546 50482
rect 58546 50430 58548 50482
rect 58492 50428 58548 50430
rect 58156 49026 58212 49028
rect 58156 48974 58158 49026
rect 58158 48974 58210 49026
rect 58210 48974 58212 49026
rect 58156 48972 58212 48974
rect 58380 49138 58436 49140
rect 58380 49086 58382 49138
rect 58382 49086 58434 49138
rect 58434 49086 58436 49138
rect 58380 49084 58436 49086
rect 58716 49196 58772 49252
rect 58492 48860 58548 48916
rect 58044 48076 58100 48132
rect 58716 48802 58772 48804
rect 58716 48750 58718 48802
rect 58718 48750 58770 48802
rect 58770 48750 58772 48802
rect 58716 48748 58772 48750
rect 59052 52108 59108 52164
rect 59612 52162 59668 52164
rect 59612 52110 59614 52162
rect 59614 52110 59666 52162
rect 59666 52110 59668 52162
rect 59612 52108 59668 52110
rect 59388 51548 59444 51604
rect 59164 51212 59220 51268
rect 61068 55186 61124 55188
rect 61068 55134 61070 55186
rect 61070 55134 61122 55186
rect 61122 55134 61124 55186
rect 61068 55132 61124 55134
rect 60060 51212 60116 51268
rect 60396 51266 60452 51268
rect 60396 51214 60398 51266
rect 60398 51214 60450 51266
rect 60450 51214 60452 51266
rect 60396 51212 60452 51214
rect 59052 49756 59108 49812
rect 59276 49138 59332 49140
rect 59276 49086 59278 49138
rect 59278 49086 59330 49138
rect 59330 49086 59332 49138
rect 59276 49084 59332 49086
rect 59052 49026 59108 49028
rect 59052 48974 59054 49026
rect 59054 48974 59106 49026
rect 59106 48974 59108 49026
rect 59052 48972 59108 48974
rect 58044 47292 58100 47348
rect 57820 46844 57876 46900
rect 57932 45836 57988 45892
rect 57708 45164 57764 45220
rect 57372 42924 57428 42980
rect 57596 44156 57652 44212
rect 57372 41858 57428 41860
rect 57372 41806 57374 41858
rect 57374 41806 57426 41858
rect 57426 41806 57428 41858
rect 57372 41804 57428 41806
rect 57820 43650 57876 43652
rect 57820 43598 57822 43650
rect 57822 43598 57874 43650
rect 57874 43598 57876 43650
rect 57820 43596 57876 43598
rect 58940 48300 58996 48356
rect 58492 48076 58548 48132
rect 58380 47516 58436 47572
rect 58492 47740 58548 47796
rect 58268 47404 58324 47460
rect 58380 46284 58436 46340
rect 58156 44716 58212 44772
rect 57820 42194 57876 42196
rect 57820 42142 57822 42194
rect 57822 42142 57874 42194
rect 57874 42142 57876 42194
rect 57820 42140 57876 42142
rect 58044 42252 58100 42308
rect 58716 46172 58772 46228
rect 59164 48748 59220 48804
rect 58940 45612 58996 45668
rect 58828 44882 58884 44884
rect 58828 44830 58830 44882
rect 58830 44830 58882 44882
rect 58882 44830 58884 44882
rect 58828 44828 58884 44830
rect 58716 43596 58772 43652
rect 57260 40236 57316 40292
rect 57260 39676 57316 39732
rect 56588 37884 56644 37940
rect 57148 39452 57204 39508
rect 56812 38220 56868 38276
rect 57260 39340 57316 39396
rect 56700 37378 56756 37380
rect 56700 37326 56702 37378
rect 56702 37326 56754 37378
rect 56754 37326 56756 37378
rect 56700 37324 56756 37326
rect 56700 36482 56756 36484
rect 56700 36430 56702 36482
rect 56702 36430 56754 36482
rect 56754 36430 56756 36482
rect 56700 36428 56756 36430
rect 56476 36092 56532 36148
rect 56924 37266 56980 37268
rect 56924 37214 56926 37266
rect 56926 37214 56978 37266
rect 56978 37214 56980 37266
rect 56924 37212 56980 37214
rect 57820 40402 57876 40404
rect 57820 40350 57822 40402
rect 57822 40350 57874 40402
rect 57874 40350 57876 40402
rect 57820 40348 57876 40350
rect 57820 39004 57876 39060
rect 57932 40124 57988 40180
rect 58156 39340 58212 39396
rect 58268 40572 58324 40628
rect 58828 41970 58884 41972
rect 58828 41918 58830 41970
rect 58830 41918 58882 41970
rect 58882 41918 58884 41970
rect 58828 41916 58884 41918
rect 59276 47682 59332 47684
rect 59276 47630 59278 47682
rect 59278 47630 59330 47682
rect 59330 47630 59332 47682
rect 59276 47628 59332 47630
rect 59612 49026 59668 49028
rect 59612 48974 59614 49026
rect 59614 48974 59666 49026
rect 59666 48974 59668 49026
rect 59612 48972 59668 48974
rect 59948 50764 60004 50820
rect 60732 53506 60788 53508
rect 60732 53454 60734 53506
rect 60734 53454 60786 53506
rect 60786 53454 60788 53506
rect 60732 53452 60788 53454
rect 61068 53452 61124 53508
rect 60732 53170 60788 53172
rect 60732 53118 60734 53170
rect 60734 53118 60786 53170
rect 60786 53118 60788 53170
rect 60732 53116 60788 53118
rect 60732 52274 60788 52276
rect 60732 52222 60734 52274
rect 60734 52222 60786 52274
rect 60786 52222 60788 52274
rect 60732 52220 60788 52222
rect 60844 51490 60900 51492
rect 60844 51438 60846 51490
rect 60846 51438 60898 51490
rect 60898 51438 60900 51490
rect 60844 51436 60900 51438
rect 60620 50876 60676 50932
rect 59948 49308 60004 49364
rect 59836 48748 59892 48804
rect 59724 48412 59780 48468
rect 59276 47068 59332 47124
rect 59612 45948 59668 46004
rect 59836 45052 59892 45108
rect 59164 42140 59220 42196
rect 59276 43260 59332 43316
rect 59052 40796 59108 40852
rect 58268 39788 58324 39844
rect 58044 38556 58100 38612
rect 58492 39004 58548 39060
rect 59052 39004 59108 39060
rect 58940 38108 58996 38164
rect 58828 38050 58884 38052
rect 58828 37998 58830 38050
rect 58830 37998 58882 38050
rect 58882 37998 58884 38050
rect 58828 37996 58884 37998
rect 57708 37884 57764 37940
rect 59500 42364 59556 42420
rect 60284 49698 60340 49700
rect 60284 49646 60286 49698
rect 60286 49646 60338 49698
rect 60338 49646 60340 49698
rect 60284 49644 60340 49646
rect 60620 50706 60676 50708
rect 60620 50654 60622 50706
rect 60622 50654 60674 50706
rect 60674 50654 60676 50706
rect 60620 50652 60676 50654
rect 61516 52274 61572 52276
rect 61516 52222 61518 52274
rect 61518 52222 61570 52274
rect 61570 52222 61572 52274
rect 61516 52220 61572 52222
rect 61404 51100 61460 51156
rect 61516 50876 61572 50932
rect 60508 48860 60564 48916
rect 60284 47068 60340 47124
rect 60732 48748 60788 48804
rect 61180 50316 61236 50372
rect 60956 48188 61012 48244
rect 62188 53506 62244 53508
rect 62188 53454 62190 53506
rect 62190 53454 62242 53506
rect 62242 53454 62244 53506
rect 62188 53452 62244 53454
rect 61740 51100 61796 51156
rect 61740 50876 61796 50932
rect 61852 50204 61908 50260
rect 61628 48748 61684 48804
rect 62636 52220 62692 52276
rect 61740 48860 61796 48916
rect 60956 47740 61012 47796
rect 61292 47628 61348 47684
rect 60620 47458 60676 47460
rect 60620 47406 60622 47458
rect 60622 47406 60674 47458
rect 60674 47406 60676 47458
rect 60620 47404 60676 47406
rect 60732 47292 60788 47348
rect 60620 47234 60676 47236
rect 60620 47182 60622 47234
rect 60622 47182 60674 47234
rect 60674 47182 60676 47234
rect 60620 47180 60676 47182
rect 60732 46956 60788 47012
rect 60620 46002 60676 46004
rect 60620 45950 60622 46002
rect 60622 45950 60674 46002
rect 60674 45950 60676 46002
rect 60620 45948 60676 45950
rect 60844 45836 60900 45892
rect 60060 42700 60116 42756
rect 59612 42028 59668 42084
rect 59724 42252 59780 42308
rect 59500 41858 59556 41860
rect 59500 41806 59502 41858
rect 59502 41806 59554 41858
rect 59554 41806 59556 41858
rect 59500 41804 59556 41806
rect 59724 41074 59780 41076
rect 59724 41022 59726 41074
rect 59726 41022 59778 41074
rect 59778 41022 59780 41074
rect 59724 41020 59780 41022
rect 59612 40796 59668 40852
rect 59500 39730 59556 39732
rect 59500 39678 59502 39730
rect 59502 39678 59554 39730
rect 59554 39678 59556 39730
rect 59500 39676 59556 39678
rect 59836 39618 59892 39620
rect 59836 39566 59838 39618
rect 59838 39566 59890 39618
rect 59890 39566 59892 39618
rect 59836 39564 59892 39566
rect 59724 39004 59780 39060
rect 59612 38892 59668 38948
rect 59276 38556 59332 38612
rect 57372 36706 57428 36708
rect 57372 36654 57374 36706
rect 57374 36654 57426 36706
rect 57426 36654 57428 36706
rect 57372 36652 57428 36654
rect 57260 36428 57316 36484
rect 57260 35868 57316 35924
rect 56252 35084 56308 35140
rect 56700 35532 56756 35588
rect 56588 34802 56644 34804
rect 56588 34750 56590 34802
rect 56590 34750 56642 34802
rect 56642 34750 56644 34802
rect 56588 34748 56644 34750
rect 56252 34690 56308 34692
rect 56252 34638 56254 34690
rect 56254 34638 56306 34690
rect 56306 34638 56308 34690
rect 56252 34636 56308 34638
rect 56140 33628 56196 33684
rect 55804 33180 55860 33236
rect 56252 33292 56308 33348
rect 56476 32508 56532 32564
rect 55692 31836 55748 31892
rect 56252 31500 56308 31556
rect 54460 27804 54516 27860
rect 54460 27468 54516 27524
rect 55468 30268 55524 30324
rect 55020 28700 55076 28756
rect 55020 28028 55076 28084
rect 54796 27916 54852 27972
rect 54684 27580 54740 27636
rect 52780 25506 52836 25508
rect 52780 25454 52782 25506
rect 52782 25454 52834 25506
rect 52834 25454 52836 25506
rect 52780 25452 52836 25454
rect 52892 25394 52948 25396
rect 52892 25342 52894 25394
rect 52894 25342 52946 25394
rect 52946 25342 52948 25394
rect 52892 25340 52948 25342
rect 53004 24722 53060 24724
rect 53004 24670 53006 24722
rect 53006 24670 53058 24722
rect 53058 24670 53060 24722
rect 53004 24668 53060 24670
rect 52892 24444 52948 24500
rect 52668 24108 52724 24164
rect 52668 22988 52724 23044
rect 52780 23996 52836 24052
rect 53340 24556 53396 24612
rect 54348 26348 54404 26404
rect 54236 25788 54292 25844
rect 53788 25676 53844 25732
rect 53676 25282 53732 25284
rect 53676 25230 53678 25282
rect 53678 25230 53730 25282
rect 53730 25230 53732 25282
rect 53676 25228 53732 25230
rect 54684 26348 54740 26404
rect 53788 25116 53844 25172
rect 54012 25004 54068 25060
rect 54684 24722 54740 24724
rect 54684 24670 54686 24722
rect 54686 24670 54738 24722
rect 54738 24670 54740 24722
rect 54684 24668 54740 24670
rect 53788 24556 53844 24612
rect 53452 23436 53508 23492
rect 53004 23212 53060 23268
rect 52892 23154 52948 23156
rect 52892 23102 52894 23154
rect 52894 23102 52946 23154
rect 52946 23102 52948 23154
rect 52892 23100 52948 23102
rect 52668 22204 52724 22260
rect 53452 22988 53508 23044
rect 52444 21644 52500 21700
rect 52668 20972 52724 21028
rect 52892 20188 52948 20244
rect 53004 21196 53060 21252
rect 52108 19404 52164 19460
rect 51548 19010 51604 19012
rect 51548 18958 51550 19010
rect 51550 18958 51602 19010
rect 51602 18958 51604 19010
rect 51548 18956 51604 18958
rect 51772 18508 51828 18564
rect 51884 18284 51940 18340
rect 51884 17948 51940 18004
rect 51660 17724 51716 17780
rect 51436 16716 51492 16772
rect 51212 16268 51268 16324
rect 50204 14924 50260 14980
rect 49756 14812 49812 14868
rect 49532 14364 49588 14420
rect 48300 13468 48356 13524
rect 48300 12850 48356 12852
rect 48300 12798 48302 12850
rect 48302 12798 48354 12850
rect 48354 12798 48356 12850
rect 48300 12796 48356 12798
rect 44604 9212 44660 9268
rect 44044 8764 44100 8820
rect 43932 8652 43988 8708
rect 44156 7756 44212 7812
rect 44492 7756 44548 7812
rect 47628 11394 47684 11396
rect 47628 11342 47630 11394
rect 47630 11342 47682 11394
rect 47682 11342 47684 11394
rect 47628 11340 47684 11342
rect 47404 11282 47460 11284
rect 47404 11230 47406 11282
rect 47406 11230 47458 11282
rect 47458 11230 47460 11282
rect 47404 11228 47460 11230
rect 47516 11170 47572 11172
rect 47516 11118 47518 11170
rect 47518 11118 47570 11170
rect 47570 11118 47572 11170
rect 47516 11116 47572 11118
rect 47628 11004 47684 11060
rect 47404 10780 47460 10836
rect 45388 9826 45444 9828
rect 45388 9774 45390 9826
rect 45390 9774 45442 9826
rect 45442 9774 45444 9826
rect 45388 9772 45444 9774
rect 45164 8988 45220 9044
rect 45276 9212 45332 9268
rect 44940 8930 44996 8932
rect 44940 8878 44942 8930
rect 44942 8878 44994 8930
rect 44994 8878 44996 8930
rect 44940 8876 44996 8878
rect 45052 8764 45108 8820
rect 44940 8652 44996 8708
rect 44492 7586 44548 7588
rect 44492 7534 44494 7586
rect 44494 7534 44546 7586
rect 44546 7534 44548 7586
rect 44492 7532 44548 7534
rect 44156 7420 44212 7476
rect 45052 8428 45108 8484
rect 45500 9154 45556 9156
rect 45500 9102 45502 9154
rect 45502 9102 45554 9154
rect 45554 9102 45556 9154
rect 45500 9100 45556 9102
rect 45612 9042 45668 9044
rect 45612 8990 45614 9042
rect 45614 8990 45666 9042
rect 45666 8990 45668 9042
rect 45612 8988 45668 8990
rect 45612 8316 45668 8372
rect 44156 6748 44212 6804
rect 44268 6524 44324 6580
rect 44156 6076 44212 6132
rect 45052 6300 45108 6356
rect 44828 5852 44884 5908
rect 44156 5628 44212 5684
rect 45052 5964 45108 6020
rect 44940 5628 44996 5684
rect 44940 5010 44996 5012
rect 44940 4958 44942 5010
rect 44942 4958 44994 5010
rect 44994 4958 44996 5010
rect 44940 4956 44996 4958
rect 44604 4508 44660 4564
rect 44268 3612 44324 3668
rect 45836 9602 45892 9604
rect 45836 9550 45838 9602
rect 45838 9550 45890 9602
rect 45890 9550 45892 9602
rect 45836 9548 45892 9550
rect 46060 9266 46116 9268
rect 46060 9214 46062 9266
rect 46062 9214 46114 9266
rect 46114 9214 46116 9266
rect 46060 9212 46116 9214
rect 45724 7868 45780 7924
rect 46060 8540 46116 8596
rect 45612 7474 45668 7476
rect 45612 7422 45614 7474
rect 45614 7422 45666 7474
rect 45666 7422 45668 7474
rect 45612 7420 45668 7422
rect 45388 6972 45444 7028
rect 45500 6860 45556 6916
rect 45276 6636 45332 6692
rect 45948 6748 46004 6804
rect 45724 6690 45780 6692
rect 45724 6638 45726 6690
rect 45726 6638 45778 6690
rect 45778 6638 45780 6690
rect 45724 6636 45780 6638
rect 46172 7196 46228 7252
rect 46172 6972 46228 7028
rect 46620 9548 46676 9604
rect 46732 9436 46788 9492
rect 47292 10610 47348 10612
rect 47292 10558 47294 10610
rect 47294 10558 47346 10610
rect 47346 10558 47348 10610
rect 47292 10556 47348 10558
rect 47404 10050 47460 10052
rect 47404 9998 47406 10050
rect 47406 9998 47458 10050
rect 47458 9998 47460 10050
rect 47404 9996 47460 9998
rect 46956 9660 47012 9716
rect 47180 9100 47236 9156
rect 46732 9042 46788 9044
rect 46732 8990 46734 9042
rect 46734 8990 46786 9042
rect 46786 8990 46788 9042
rect 46732 8988 46788 8990
rect 46956 8988 47012 9044
rect 46284 6860 46340 6916
rect 46508 6636 46564 6692
rect 45612 5964 45668 6020
rect 45836 5906 45892 5908
rect 45836 5854 45838 5906
rect 45838 5854 45890 5906
rect 45890 5854 45892 5906
rect 45836 5852 45892 5854
rect 45724 5628 45780 5684
rect 45724 4508 45780 4564
rect 46620 7084 46676 7140
rect 46396 6076 46452 6132
rect 46172 5906 46228 5908
rect 46172 5854 46174 5906
rect 46174 5854 46226 5906
rect 46226 5854 46228 5906
rect 46172 5852 46228 5854
rect 47404 7474 47460 7476
rect 47404 7422 47406 7474
rect 47406 7422 47458 7474
rect 47458 7422 47460 7474
rect 47404 7420 47460 7422
rect 47516 7196 47572 7252
rect 47068 6076 47124 6132
rect 47292 6188 47348 6244
rect 46844 5122 46900 5124
rect 46844 5070 46846 5122
rect 46846 5070 46898 5122
rect 46898 5070 46900 5122
rect 46844 5068 46900 5070
rect 46732 4338 46788 4340
rect 46732 4286 46734 4338
rect 46734 4286 46786 4338
rect 46786 4286 46788 4338
rect 46732 4284 46788 4286
rect 46508 3666 46564 3668
rect 46508 3614 46510 3666
rect 46510 3614 46562 3666
rect 46562 3614 46564 3666
rect 46508 3612 46564 3614
rect 46956 4508 47012 4564
rect 47292 5292 47348 5348
rect 48076 11452 48132 11508
rect 47852 10892 47908 10948
rect 48188 11340 48244 11396
rect 48300 11170 48356 11172
rect 48300 11118 48302 11170
rect 48302 11118 48354 11170
rect 48354 11118 48356 11170
rect 48300 11116 48356 11118
rect 48748 11452 48804 11508
rect 49196 12850 49252 12852
rect 49196 12798 49198 12850
rect 49198 12798 49250 12850
rect 49250 12798 49252 12850
rect 49196 12796 49252 12798
rect 49420 12460 49476 12516
rect 48972 11394 49028 11396
rect 48972 11342 48974 11394
rect 48974 11342 49026 11394
rect 49026 11342 49028 11394
rect 48972 11340 49028 11342
rect 49420 11506 49476 11508
rect 49420 11454 49422 11506
rect 49422 11454 49474 11506
rect 49474 11454 49476 11506
rect 49420 11452 49476 11454
rect 49308 11340 49364 11396
rect 48860 11116 48916 11172
rect 48524 10892 48580 10948
rect 48860 10892 48916 10948
rect 48188 10780 48244 10836
rect 47964 10668 48020 10724
rect 48972 10610 49028 10612
rect 48972 10558 48974 10610
rect 48974 10558 49026 10610
rect 49026 10558 49028 10610
rect 48972 10556 49028 10558
rect 47964 8988 48020 9044
rect 47852 8930 47908 8932
rect 47852 8878 47854 8930
rect 47854 8878 47906 8930
rect 47906 8878 47908 8930
rect 47852 8876 47908 8878
rect 47740 8482 47796 8484
rect 47740 8430 47742 8482
rect 47742 8430 47794 8482
rect 47794 8430 47796 8482
rect 47740 8428 47796 8430
rect 48860 9714 48916 9716
rect 48860 9662 48862 9714
rect 48862 9662 48914 9714
rect 48914 9662 48916 9714
rect 48860 9660 48916 9662
rect 48748 9042 48804 9044
rect 48748 8990 48750 9042
rect 48750 8990 48802 9042
rect 48802 8990 48804 9042
rect 48748 8988 48804 8990
rect 48748 8428 48804 8484
rect 47964 7532 48020 7588
rect 47740 7308 47796 7364
rect 47740 6636 47796 6692
rect 47852 6748 47908 6804
rect 48188 7362 48244 7364
rect 48188 7310 48190 7362
rect 48190 7310 48242 7362
rect 48242 7310 48244 7362
rect 48188 7308 48244 7310
rect 48412 6860 48468 6916
rect 48860 8258 48916 8260
rect 48860 8206 48862 8258
rect 48862 8206 48914 8258
rect 48914 8206 48916 8258
rect 48860 8204 48916 8206
rect 50428 15314 50484 15316
rect 50428 15262 50430 15314
rect 50430 15262 50482 15314
rect 50482 15262 50484 15314
rect 50428 15260 50484 15262
rect 50092 13692 50148 13748
rect 49980 13074 50036 13076
rect 49980 13022 49982 13074
rect 49982 13022 50034 13074
rect 50034 13022 50036 13074
rect 49980 13020 50036 13022
rect 50652 14700 50708 14756
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50652 13970 50708 13972
rect 50652 13918 50654 13970
rect 50654 13918 50706 13970
rect 50706 13918 50708 13970
rect 50652 13916 50708 13918
rect 50428 13692 50484 13748
rect 50092 12348 50148 12404
rect 50204 13468 50260 13524
rect 49868 11116 49924 11172
rect 49532 10556 49588 10612
rect 49308 10332 49364 10388
rect 49420 10444 49476 10500
rect 49420 8204 49476 8260
rect 49308 8092 49364 8148
rect 49196 8034 49252 8036
rect 49196 7982 49198 8034
rect 49198 7982 49250 8034
rect 49250 7982 49252 8034
rect 49196 7980 49252 7982
rect 49196 7756 49252 7812
rect 48860 7362 48916 7364
rect 48860 7310 48862 7362
rect 48862 7310 48914 7362
rect 48914 7310 48916 7362
rect 48860 7308 48916 7310
rect 48188 6076 48244 6132
rect 48076 6018 48132 6020
rect 48076 5966 48078 6018
rect 48078 5966 48130 6018
rect 48130 5966 48132 6018
rect 48076 5964 48132 5966
rect 49084 6412 49140 6468
rect 49308 6972 49364 7028
rect 48748 6018 48804 6020
rect 48748 5966 48750 6018
rect 48750 5966 48802 6018
rect 48802 5966 48804 6018
rect 48748 5964 48804 5966
rect 48524 4956 48580 5012
rect 47964 4620 48020 4676
rect 48076 4450 48132 4452
rect 48076 4398 48078 4450
rect 48078 4398 48130 4450
rect 48130 4398 48132 4450
rect 48076 4396 48132 4398
rect 49644 8930 49700 8932
rect 49644 8878 49646 8930
rect 49646 8878 49698 8930
rect 49698 8878 49700 8930
rect 49644 8876 49700 8878
rect 49980 7586 50036 7588
rect 49980 7534 49982 7586
rect 49982 7534 50034 7586
rect 50034 7534 50036 7586
rect 49980 7532 50036 7534
rect 51548 16492 51604 16548
rect 52556 18508 52612 18564
rect 52220 18226 52276 18228
rect 52220 18174 52222 18226
rect 52222 18174 52274 18226
rect 52274 18174 52276 18226
rect 52220 18172 52276 18174
rect 52108 17836 52164 17892
rect 52892 18396 52948 18452
rect 53228 21868 53284 21924
rect 53340 21756 53396 21812
rect 55580 30098 55636 30100
rect 55580 30046 55582 30098
rect 55582 30046 55634 30098
rect 55634 30046 55636 30098
rect 55580 30044 55636 30046
rect 55468 29426 55524 29428
rect 55468 29374 55470 29426
rect 55470 29374 55522 29426
rect 55522 29374 55524 29426
rect 55468 29372 55524 29374
rect 55468 29036 55524 29092
rect 55244 28364 55300 28420
rect 55356 27746 55412 27748
rect 55356 27694 55358 27746
rect 55358 27694 55410 27746
rect 55410 27694 55412 27746
rect 55356 27692 55412 27694
rect 56028 30210 56084 30212
rect 56028 30158 56030 30210
rect 56030 30158 56082 30210
rect 56082 30158 56084 30210
rect 56028 30156 56084 30158
rect 55804 29986 55860 29988
rect 55804 29934 55806 29986
rect 55806 29934 55858 29986
rect 55858 29934 55860 29986
rect 55804 29932 55860 29934
rect 56028 29932 56084 29988
rect 55916 29538 55972 29540
rect 55916 29486 55918 29538
rect 55918 29486 55970 29538
rect 55970 29486 55972 29538
rect 55916 29484 55972 29486
rect 55804 29148 55860 29204
rect 56588 31500 56644 31556
rect 56588 31276 56644 31332
rect 56252 28924 56308 28980
rect 56476 30210 56532 30212
rect 56476 30158 56478 30210
rect 56478 30158 56530 30210
rect 56530 30158 56532 30210
rect 56476 30156 56532 30158
rect 55804 28530 55860 28532
rect 55804 28478 55806 28530
rect 55806 28478 55858 28530
rect 55858 28478 55860 28530
rect 55804 28476 55860 28478
rect 55468 27580 55524 27636
rect 55580 28140 55636 28196
rect 55356 27244 55412 27300
rect 55804 27244 55860 27300
rect 54908 25676 54964 25732
rect 55132 26236 55188 26292
rect 55132 25618 55188 25620
rect 55132 25566 55134 25618
rect 55134 25566 55186 25618
rect 55186 25566 55188 25618
rect 55132 25564 55188 25566
rect 55132 25340 55188 25396
rect 55580 26572 55636 26628
rect 55804 26402 55860 26404
rect 55804 26350 55806 26402
rect 55806 26350 55858 26402
rect 55858 26350 55860 26402
rect 55804 26348 55860 26350
rect 54796 24220 54852 24276
rect 54796 23938 54852 23940
rect 54796 23886 54798 23938
rect 54798 23886 54850 23938
rect 54850 23886 54852 23938
rect 54796 23884 54852 23886
rect 53788 23660 53844 23716
rect 54236 23660 54292 23716
rect 54348 23324 54404 23380
rect 54572 23212 54628 23268
rect 54796 23042 54852 23044
rect 54796 22990 54798 23042
rect 54798 22990 54850 23042
rect 54850 22990 54852 23042
rect 54796 22988 54852 22990
rect 54012 21868 54068 21924
rect 55692 25564 55748 25620
rect 55692 24220 55748 24276
rect 55468 23884 55524 23940
rect 53452 21308 53508 21364
rect 53676 21308 53732 21364
rect 53900 21420 53956 21476
rect 54012 21196 54068 21252
rect 54460 21362 54516 21364
rect 54460 21310 54462 21362
rect 54462 21310 54514 21362
rect 54514 21310 54516 21362
rect 54460 21308 54516 21310
rect 55356 21810 55412 21812
rect 55356 21758 55358 21810
rect 55358 21758 55410 21810
rect 55410 21758 55412 21810
rect 55356 21756 55412 21758
rect 55020 21586 55076 21588
rect 55020 21534 55022 21586
rect 55022 21534 55074 21586
rect 55074 21534 55076 21586
rect 55020 21532 55076 21534
rect 55244 21644 55300 21700
rect 54684 21196 54740 21252
rect 54348 20860 54404 20916
rect 54124 20748 54180 20804
rect 53676 20018 53732 20020
rect 53676 19966 53678 20018
rect 53678 19966 53730 20018
rect 53730 19966 53732 20018
rect 53676 19964 53732 19966
rect 54460 20076 54516 20132
rect 54572 20636 54628 20692
rect 55020 20188 55076 20244
rect 54572 19852 54628 19908
rect 53116 19068 53172 19124
rect 53228 18956 53284 19012
rect 53116 18284 53172 18340
rect 53340 18172 53396 18228
rect 53228 17554 53284 17556
rect 53228 17502 53230 17554
rect 53230 17502 53282 17554
rect 53282 17502 53284 17554
rect 53228 17500 53284 17502
rect 51996 16828 52052 16884
rect 51884 16380 51940 16436
rect 51548 15932 51604 15988
rect 51772 16268 51828 16324
rect 51212 15484 51268 15540
rect 50988 15426 51044 15428
rect 50988 15374 50990 15426
rect 50990 15374 51042 15426
rect 51042 15374 51044 15426
rect 50988 15372 51044 15374
rect 51548 15426 51604 15428
rect 51548 15374 51550 15426
rect 51550 15374 51602 15426
rect 51602 15374 51604 15426
rect 51548 15372 51604 15374
rect 51660 14140 51716 14196
rect 50652 12850 50708 12852
rect 50652 12798 50654 12850
rect 50654 12798 50706 12850
rect 50706 12798 50708 12850
rect 50652 12796 50708 12798
rect 50428 12738 50484 12740
rect 50428 12686 50430 12738
rect 50430 12686 50482 12738
rect 50482 12686 50484 12738
rect 50428 12684 50484 12686
rect 50316 12460 50372 12516
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 51884 15148 51940 15204
rect 53116 15820 53172 15876
rect 52780 15484 52836 15540
rect 53116 15372 53172 15428
rect 52332 15202 52388 15204
rect 52332 15150 52334 15202
rect 52334 15150 52386 15202
rect 52386 15150 52388 15202
rect 52332 15148 52388 15150
rect 51212 12290 51268 12292
rect 51212 12238 51214 12290
rect 51214 12238 51266 12290
rect 51266 12238 51268 12290
rect 51212 12236 51268 12238
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50428 10108 50484 10164
rect 50652 10610 50708 10612
rect 50652 10558 50654 10610
rect 50654 10558 50706 10610
rect 50706 10558 50708 10610
rect 50652 10556 50708 10558
rect 50876 9660 50932 9716
rect 50988 11340 51044 11396
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 51212 11116 51268 11172
rect 51436 11004 51492 11060
rect 51772 9772 51828 9828
rect 51660 9714 51716 9716
rect 51660 9662 51662 9714
rect 51662 9662 51714 9714
rect 51714 9662 51716 9714
rect 51660 9660 51716 9662
rect 51548 8988 51604 9044
rect 50428 8092 50484 8148
rect 50204 7308 50260 7364
rect 49532 6412 49588 6468
rect 49420 6188 49476 6244
rect 52892 14140 52948 14196
rect 52108 13916 52164 13972
rect 51996 11340 52052 11396
rect 51996 9826 52052 9828
rect 51996 9774 51998 9826
rect 51998 9774 52050 9826
rect 52050 9774 52052 9826
rect 51996 9772 52052 9774
rect 51660 7980 51716 8036
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 51660 7698 51716 7700
rect 51660 7646 51662 7698
rect 51662 7646 51714 7698
rect 51714 7646 51716 7698
rect 51660 7644 51716 7646
rect 51100 7420 51156 7476
rect 50764 6690 50820 6692
rect 50764 6638 50766 6690
rect 50766 6638 50818 6690
rect 50818 6638 50820 6690
rect 50764 6636 50820 6638
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 50316 6130 50372 6132
rect 50316 6078 50318 6130
rect 50318 6078 50370 6130
rect 50370 6078 50372 6130
rect 50316 6076 50372 6078
rect 50764 5180 50820 5236
rect 50204 5122 50260 5124
rect 50204 5070 50206 5122
rect 50206 5070 50258 5122
rect 50258 5070 50260 5122
rect 50204 5068 50260 5070
rect 51212 7084 51268 7140
rect 51660 6972 51716 7028
rect 51100 5068 51156 5124
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 48524 3666 48580 3668
rect 48524 3614 48526 3666
rect 48526 3614 48578 3666
rect 48578 3614 48580 3666
rect 48524 3612 48580 3614
rect 49308 4226 49364 4228
rect 49308 4174 49310 4226
rect 49310 4174 49362 4226
rect 49362 4174 49364 4226
rect 49308 4172 49364 4174
rect 46844 3500 46900 3556
rect 47516 3554 47572 3556
rect 47516 3502 47518 3554
rect 47518 3502 47570 3554
rect 47570 3502 47572 3554
rect 47516 3500 47572 3502
rect 49308 3500 49364 3556
rect 51996 8370 52052 8372
rect 51996 8318 51998 8370
rect 51998 8318 52050 8370
rect 52050 8318 52052 8370
rect 51996 8316 52052 8318
rect 52332 13858 52388 13860
rect 52332 13806 52334 13858
rect 52334 13806 52386 13858
rect 52386 13806 52388 13858
rect 52332 13804 52388 13806
rect 52556 13746 52612 13748
rect 52556 13694 52558 13746
rect 52558 13694 52610 13746
rect 52610 13694 52612 13746
rect 52556 13692 52612 13694
rect 52220 11004 52276 11060
rect 53004 12012 53060 12068
rect 52780 11170 52836 11172
rect 52780 11118 52782 11170
rect 52782 11118 52834 11170
rect 52834 11118 52836 11170
rect 52780 11116 52836 11118
rect 52892 11004 52948 11060
rect 52444 10556 52500 10612
rect 52556 10386 52612 10388
rect 52556 10334 52558 10386
rect 52558 10334 52610 10386
rect 52610 10334 52612 10386
rect 52556 10332 52612 10334
rect 52780 10556 52836 10612
rect 53116 11340 53172 11396
rect 52780 9826 52836 9828
rect 52780 9774 52782 9826
rect 52782 9774 52834 9826
rect 52834 9774 52836 9826
rect 52780 9772 52836 9774
rect 52668 9042 52724 9044
rect 52668 8990 52670 9042
rect 52670 8990 52722 9042
rect 52722 8990 52724 9042
rect 52668 8988 52724 8990
rect 53340 16940 53396 16996
rect 54348 19068 54404 19124
rect 53676 18844 53732 18900
rect 53788 18674 53844 18676
rect 53788 18622 53790 18674
rect 53790 18622 53842 18674
rect 53842 18622 53844 18674
rect 53788 18620 53844 18622
rect 53564 18284 53620 18340
rect 53564 17836 53620 17892
rect 53676 17948 53732 18004
rect 53788 17724 53844 17780
rect 53788 17106 53844 17108
rect 53788 17054 53790 17106
rect 53790 17054 53842 17106
rect 53842 17054 53844 17106
rect 53788 17052 53844 17054
rect 53452 16156 53508 16212
rect 53452 15932 53508 15988
rect 53564 15426 53620 15428
rect 53564 15374 53566 15426
rect 53566 15374 53618 15426
rect 53618 15374 53620 15426
rect 53564 15372 53620 15374
rect 53676 15148 53732 15204
rect 53340 14252 53396 14308
rect 54348 18226 54404 18228
rect 54348 18174 54350 18226
rect 54350 18174 54402 18226
rect 54402 18174 54404 18226
rect 54348 18172 54404 18174
rect 54012 16044 54068 16100
rect 53340 13746 53396 13748
rect 53340 13694 53342 13746
rect 53342 13694 53394 13746
rect 53394 13694 53396 13746
rect 53340 13692 53396 13694
rect 53900 14364 53956 14420
rect 54012 14028 54068 14084
rect 53788 13468 53844 13524
rect 53340 13074 53396 13076
rect 53340 13022 53342 13074
rect 53342 13022 53394 13074
rect 53394 13022 53396 13074
rect 53340 13020 53396 13022
rect 53340 12684 53396 12740
rect 53340 9212 53396 9268
rect 53004 8316 53060 8372
rect 53676 8764 53732 8820
rect 55580 22988 55636 23044
rect 54684 19180 54740 19236
rect 54908 18450 54964 18452
rect 54908 18398 54910 18450
rect 54910 18398 54962 18450
rect 54962 18398 54964 18450
rect 54908 18396 54964 18398
rect 56252 28754 56308 28756
rect 56252 28702 56254 28754
rect 56254 28702 56306 28754
rect 56306 28702 56308 28754
rect 56252 28700 56308 28702
rect 57260 35308 57316 35364
rect 56812 35196 56868 35252
rect 58380 36204 58436 36260
rect 57484 35196 57540 35252
rect 58044 35084 58100 35140
rect 56924 34914 56980 34916
rect 56924 34862 56926 34914
rect 56926 34862 56978 34914
rect 56978 34862 56980 34914
rect 56924 34860 56980 34862
rect 58492 35980 58548 36036
rect 58828 35698 58884 35700
rect 58828 35646 58830 35698
rect 58830 35646 58882 35698
rect 58882 35646 58884 35698
rect 58828 35644 58884 35646
rect 58716 35084 58772 35140
rect 56924 34636 56980 34692
rect 56812 33346 56868 33348
rect 56812 33294 56814 33346
rect 56814 33294 56866 33346
rect 56866 33294 56868 33346
rect 56812 33292 56868 33294
rect 56812 32732 56868 32788
rect 57036 34524 57092 34580
rect 58268 34636 58324 34692
rect 57148 34300 57204 34356
rect 57036 33852 57092 33908
rect 59500 38108 59556 38164
rect 59500 37436 59556 37492
rect 59276 36764 59332 36820
rect 59500 37100 59556 37156
rect 59612 36988 59668 37044
rect 60060 36428 60116 36484
rect 59612 34860 59668 34916
rect 59388 34188 59444 34244
rect 57148 33516 57204 33572
rect 56812 32060 56868 32116
rect 58156 33346 58212 33348
rect 58156 33294 58158 33346
rect 58158 33294 58210 33346
rect 58210 33294 58212 33346
rect 58156 33292 58212 33294
rect 57484 32786 57540 32788
rect 57484 32734 57486 32786
rect 57486 32734 57538 32786
rect 57538 32734 57540 32786
rect 57484 32732 57540 32734
rect 57148 31500 57204 31556
rect 56812 30380 56868 30436
rect 57036 30268 57092 30324
rect 56924 30044 56980 30100
rect 56700 29372 56756 29428
rect 56924 29484 56980 29540
rect 56588 29036 56644 29092
rect 56588 28812 56644 28868
rect 56476 28476 56532 28532
rect 56476 28252 56532 28308
rect 56028 26290 56084 26292
rect 56028 26238 56030 26290
rect 56030 26238 56082 26290
rect 56082 26238 56084 26290
rect 56028 26236 56084 26238
rect 56028 26012 56084 26068
rect 56028 25788 56084 25844
rect 56028 22988 56084 23044
rect 55804 22316 55860 22372
rect 56028 22204 56084 22260
rect 55804 20972 55860 21028
rect 55692 19964 55748 20020
rect 55804 19068 55860 19124
rect 56364 28028 56420 28084
rect 56812 28588 56868 28644
rect 57484 31890 57540 31892
rect 57484 31838 57486 31890
rect 57486 31838 57538 31890
rect 57538 31838 57540 31890
rect 57484 31836 57540 31838
rect 57596 31500 57652 31556
rect 57820 31724 57876 31780
rect 57932 31276 57988 31332
rect 58492 32562 58548 32564
rect 58492 32510 58494 32562
rect 58494 32510 58546 32562
rect 58546 32510 58548 32562
rect 58492 32508 58548 32510
rect 57708 30380 57764 30436
rect 57260 29202 57316 29204
rect 57260 29150 57262 29202
rect 57262 29150 57314 29202
rect 57314 29150 57316 29202
rect 57260 29148 57316 29150
rect 57148 28364 57204 28420
rect 57596 29426 57652 29428
rect 57596 29374 57598 29426
rect 57598 29374 57650 29426
rect 57650 29374 57652 29426
rect 57596 29372 57652 29374
rect 57036 28252 57092 28308
rect 56812 27244 56868 27300
rect 56476 26908 56532 26964
rect 56700 26572 56756 26628
rect 57036 26908 57092 26964
rect 57148 26796 57204 26852
rect 56476 25676 56532 25732
rect 56924 25788 56980 25844
rect 56588 24220 56644 24276
rect 56364 23714 56420 23716
rect 56364 23662 56366 23714
rect 56366 23662 56418 23714
rect 56418 23662 56420 23714
rect 56364 23660 56420 23662
rect 56812 25228 56868 25284
rect 57260 26348 57316 26404
rect 58044 29426 58100 29428
rect 58044 29374 58046 29426
rect 58046 29374 58098 29426
rect 58098 29374 58100 29426
rect 58044 29372 58100 29374
rect 57708 28140 57764 28196
rect 57932 28588 57988 28644
rect 57596 27916 57652 27972
rect 57596 27468 57652 27524
rect 57484 26460 57540 26516
rect 57372 26236 57428 26292
rect 57260 25228 57316 25284
rect 57260 25004 57316 25060
rect 57036 24946 57092 24948
rect 57036 24894 57038 24946
rect 57038 24894 57090 24946
rect 57090 24894 57092 24946
rect 57036 24892 57092 24894
rect 57148 24834 57204 24836
rect 57148 24782 57150 24834
rect 57150 24782 57202 24834
rect 57202 24782 57204 24834
rect 57148 24780 57204 24782
rect 56924 24444 56980 24500
rect 56924 24220 56980 24276
rect 56588 23436 56644 23492
rect 57148 24050 57204 24052
rect 57148 23998 57150 24050
rect 57150 23998 57202 24050
rect 57202 23998 57204 24050
rect 57148 23996 57204 23998
rect 57036 23772 57092 23828
rect 57260 23436 57316 23492
rect 57036 22988 57092 23044
rect 56252 20860 56308 20916
rect 57260 22876 57316 22932
rect 57036 21980 57092 22036
rect 57148 22092 57204 22148
rect 56140 20188 56196 20244
rect 56588 20636 56644 20692
rect 57036 20018 57092 20020
rect 57036 19966 57038 20018
rect 57038 19966 57090 20018
rect 57090 19966 57092 20018
rect 57036 19964 57092 19966
rect 56588 19906 56644 19908
rect 56588 19854 56590 19906
rect 56590 19854 56642 19906
rect 56642 19854 56644 19906
rect 56588 19852 56644 19854
rect 56252 19234 56308 19236
rect 56252 19182 56254 19234
rect 56254 19182 56306 19234
rect 56306 19182 56308 19234
rect 56252 19180 56308 19182
rect 56252 18620 56308 18676
rect 56700 19180 56756 19236
rect 55692 18172 55748 18228
rect 55580 18060 55636 18116
rect 54460 17554 54516 17556
rect 54460 17502 54462 17554
rect 54462 17502 54514 17554
rect 54514 17502 54516 17554
rect 54460 17500 54516 17502
rect 54348 17442 54404 17444
rect 54348 17390 54350 17442
rect 54350 17390 54402 17442
rect 54402 17390 54404 17442
rect 54348 17388 54404 17390
rect 54572 17106 54628 17108
rect 54572 17054 54574 17106
rect 54574 17054 54626 17106
rect 54626 17054 54628 17106
rect 54572 17052 54628 17054
rect 54460 16770 54516 16772
rect 54460 16718 54462 16770
rect 54462 16718 54514 16770
rect 54514 16718 54516 16770
rect 54460 16716 54516 16718
rect 54796 16044 54852 16100
rect 54908 16716 54964 16772
rect 55468 16716 55524 16772
rect 55356 15932 55412 15988
rect 55356 15260 55412 15316
rect 56364 18396 56420 18452
rect 55916 16994 55972 16996
rect 55916 16942 55918 16994
rect 55918 16942 55970 16994
rect 55970 16942 55972 16994
rect 55916 16940 55972 16942
rect 55804 16156 55860 16212
rect 56140 16716 56196 16772
rect 56252 18060 56308 18116
rect 56140 16156 56196 16212
rect 56140 15260 56196 15316
rect 56588 18172 56644 18228
rect 56476 17164 56532 17220
rect 56252 14700 56308 14756
rect 56364 15372 56420 15428
rect 55020 14364 55076 14420
rect 55916 14252 55972 14308
rect 54236 13020 54292 13076
rect 54124 12962 54180 12964
rect 54124 12910 54126 12962
rect 54126 12910 54178 12962
rect 54178 12910 54180 12962
rect 54124 12908 54180 12910
rect 54124 12684 54180 12740
rect 54348 11004 54404 11060
rect 54124 10610 54180 10612
rect 54124 10558 54126 10610
rect 54126 10558 54178 10610
rect 54178 10558 54180 10610
rect 54124 10556 54180 10558
rect 55356 13746 55412 13748
rect 55356 13694 55358 13746
rect 55358 13694 55410 13746
rect 55410 13694 55412 13746
rect 55356 13692 55412 13694
rect 55804 13020 55860 13076
rect 55244 12908 55300 12964
rect 55692 12908 55748 12964
rect 55020 12684 55076 12740
rect 55468 12402 55524 12404
rect 55468 12350 55470 12402
rect 55470 12350 55522 12402
rect 55522 12350 55524 12402
rect 55468 12348 55524 12350
rect 55804 12348 55860 12404
rect 56252 12850 56308 12852
rect 56252 12798 56254 12850
rect 56254 12798 56306 12850
rect 56306 12798 56308 12850
rect 56252 12796 56308 12798
rect 56812 19068 56868 19124
rect 57484 23212 57540 23268
rect 57708 27356 57764 27412
rect 58044 28476 58100 28532
rect 58380 31500 58436 31556
rect 59612 33906 59668 33908
rect 59612 33854 59614 33906
rect 59614 33854 59666 33906
rect 59666 33854 59668 33906
rect 59612 33852 59668 33854
rect 60284 44940 60340 44996
rect 60620 44716 60676 44772
rect 61068 47516 61124 47572
rect 61516 47628 61572 47684
rect 61516 46956 61572 47012
rect 62076 48354 62132 48356
rect 62076 48302 62078 48354
rect 62078 48302 62130 48354
rect 62130 48302 62132 48354
rect 62076 48300 62132 48302
rect 61740 46844 61796 46900
rect 61964 48188 62020 48244
rect 62076 47852 62132 47908
rect 61964 46956 62020 47012
rect 61404 46620 61460 46676
rect 61292 46562 61348 46564
rect 61292 46510 61294 46562
rect 61294 46510 61346 46562
rect 61346 46510 61348 46562
rect 61292 46508 61348 46510
rect 61516 46284 61572 46340
rect 61740 46284 61796 46340
rect 61292 45890 61348 45892
rect 61292 45838 61294 45890
rect 61294 45838 61346 45890
rect 61346 45838 61348 45890
rect 61292 45836 61348 45838
rect 61628 45666 61684 45668
rect 61628 45614 61630 45666
rect 61630 45614 61682 45666
rect 61682 45614 61684 45666
rect 61628 45612 61684 45614
rect 61628 45218 61684 45220
rect 61628 45166 61630 45218
rect 61630 45166 61682 45218
rect 61682 45166 61684 45218
rect 61628 45164 61684 45166
rect 61404 45052 61460 45108
rect 60844 44268 60900 44324
rect 60508 41186 60564 41188
rect 60508 41134 60510 41186
rect 60510 41134 60562 41186
rect 60562 41134 60564 41186
rect 60508 41132 60564 41134
rect 60620 40514 60676 40516
rect 60620 40462 60622 40514
rect 60622 40462 60674 40514
rect 60674 40462 60676 40514
rect 60620 40460 60676 40462
rect 60396 40236 60452 40292
rect 60508 40124 60564 40180
rect 60956 42812 61012 42868
rect 61292 42700 61348 42756
rect 61516 43596 61572 43652
rect 62188 47346 62244 47348
rect 62188 47294 62190 47346
rect 62190 47294 62242 47346
rect 62242 47294 62244 47346
rect 62188 47292 62244 47294
rect 61964 43484 62020 43540
rect 62188 45890 62244 45892
rect 62188 45838 62190 45890
rect 62190 45838 62242 45890
rect 62242 45838 62244 45890
rect 62188 45836 62244 45838
rect 62076 44828 62132 44884
rect 61964 43314 62020 43316
rect 61964 43262 61966 43314
rect 61966 43262 62018 43314
rect 62018 43262 62020 43314
rect 61964 43260 62020 43262
rect 61516 42812 61572 42868
rect 61628 42700 61684 42756
rect 61292 42364 61348 42420
rect 61180 41916 61236 41972
rect 60956 41356 61012 41412
rect 61068 41804 61124 41860
rect 61180 41468 61236 41524
rect 60956 40962 61012 40964
rect 60956 40910 60958 40962
rect 60958 40910 61010 40962
rect 61010 40910 61012 40962
rect 60956 40908 61012 40910
rect 61068 40796 61124 40852
rect 61068 40348 61124 40404
rect 61180 40572 61236 40628
rect 60956 39788 61012 39844
rect 60508 38946 60564 38948
rect 60508 38894 60510 38946
rect 60510 38894 60562 38946
rect 60562 38894 60564 38946
rect 60508 38892 60564 38894
rect 60956 38892 61012 38948
rect 60732 38834 60788 38836
rect 60732 38782 60734 38834
rect 60734 38782 60786 38834
rect 60786 38782 60788 38834
rect 60732 38780 60788 38782
rect 59724 32284 59780 32340
rect 58828 31724 58884 31780
rect 59612 30994 59668 30996
rect 59612 30942 59614 30994
rect 59614 30942 59666 30994
rect 59666 30942 59668 30994
rect 59612 30940 59668 30942
rect 59276 30492 59332 30548
rect 60172 31724 60228 31780
rect 60508 38050 60564 38052
rect 60508 37998 60510 38050
rect 60510 37998 60562 38050
rect 60562 37998 60564 38050
rect 60508 37996 60564 37998
rect 60956 37996 61012 38052
rect 60844 37938 60900 37940
rect 60844 37886 60846 37938
rect 60846 37886 60898 37938
rect 60898 37886 60900 37938
rect 60844 37884 60900 37886
rect 60396 37436 60452 37492
rect 60620 37324 60676 37380
rect 60620 36988 60676 37044
rect 60508 36258 60564 36260
rect 60508 36206 60510 36258
rect 60510 36206 60562 36258
rect 60562 36206 60564 36258
rect 60508 36204 60564 36206
rect 61068 37436 61124 37492
rect 61068 36540 61124 36596
rect 60956 36428 61012 36484
rect 60844 36092 60900 36148
rect 60732 35980 60788 36036
rect 60732 34914 60788 34916
rect 60732 34862 60734 34914
rect 60734 34862 60786 34914
rect 60786 34862 60788 34914
rect 60732 34860 60788 34862
rect 60732 34242 60788 34244
rect 60732 34190 60734 34242
rect 60734 34190 60786 34242
rect 60786 34190 60788 34242
rect 60732 34188 60788 34190
rect 60508 33516 60564 33572
rect 60732 33346 60788 33348
rect 60732 33294 60734 33346
rect 60734 33294 60786 33346
rect 60786 33294 60788 33346
rect 60732 33292 60788 33294
rect 60508 33234 60564 33236
rect 60508 33182 60510 33234
rect 60510 33182 60562 33234
rect 60562 33182 60564 33234
rect 60508 33180 60564 33182
rect 60508 32562 60564 32564
rect 60508 32510 60510 32562
rect 60510 32510 60562 32562
rect 60562 32510 60564 32562
rect 60508 32508 60564 32510
rect 61628 41858 61684 41860
rect 61628 41806 61630 41858
rect 61630 41806 61682 41858
rect 61682 41806 61684 41858
rect 61628 41804 61684 41806
rect 61404 41020 61460 41076
rect 61404 40460 61460 40516
rect 61628 41356 61684 41412
rect 61516 40348 61572 40404
rect 61404 39228 61460 39284
rect 61404 38834 61460 38836
rect 61404 38782 61406 38834
rect 61406 38782 61458 38834
rect 61458 38782 61460 38834
rect 61404 38780 61460 38782
rect 61292 38050 61348 38052
rect 61292 37998 61294 38050
rect 61294 37998 61346 38050
rect 61346 37998 61348 38050
rect 61292 37996 61348 37998
rect 61292 36482 61348 36484
rect 61292 36430 61294 36482
rect 61294 36430 61346 36482
rect 61346 36430 61348 36482
rect 61292 36428 61348 36430
rect 61292 35196 61348 35252
rect 61740 41244 61796 41300
rect 61740 40684 61796 40740
rect 61740 40460 61796 40516
rect 62076 41970 62132 41972
rect 62076 41918 62078 41970
rect 62078 41918 62130 41970
rect 62130 41918 62132 41970
rect 62076 41916 62132 41918
rect 62076 40402 62132 40404
rect 62076 40350 62078 40402
rect 62078 40350 62130 40402
rect 62130 40350 62132 40402
rect 62076 40348 62132 40350
rect 62300 41692 62356 41748
rect 62300 40572 62356 40628
rect 62412 42140 62468 42196
rect 62188 40236 62244 40292
rect 61964 40124 62020 40180
rect 61628 37436 61684 37492
rect 61852 38892 61908 38948
rect 62076 37266 62132 37268
rect 62076 37214 62078 37266
rect 62078 37214 62130 37266
rect 62130 37214 62132 37266
rect 62076 37212 62132 37214
rect 61516 36370 61572 36372
rect 61516 36318 61518 36370
rect 61518 36318 61570 36370
rect 61570 36318 61572 36370
rect 61516 36316 61572 36318
rect 61628 36092 61684 36148
rect 61740 36764 61796 36820
rect 61964 36764 62020 36820
rect 61964 36540 62020 36596
rect 62188 35922 62244 35924
rect 62188 35870 62190 35922
rect 62190 35870 62242 35922
rect 62242 35870 62244 35922
rect 62188 35868 62244 35870
rect 61740 34242 61796 34244
rect 61740 34190 61742 34242
rect 61742 34190 61794 34242
rect 61794 34190 61796 34242
rect 61740 34188 61796 34190
rect 61740 33346 61796 33348
rect 61740 33294 61742 33346
rect 61742 33294 61794 33346
rect 61794 33294 61796 33346
rect 61740 33292 61796 33294
rect 61180 32508 61236 32564
rect 60508 31276 60564 31332
rect 60284 30716 60340 30772
rect 59948 30492 60004 30548
rect 59724 30044 59780 30100
rect 60284 30156 60340 30212
rect 59612 29596 59668 29652
rect 58828 29484 58884 29540
rect 58716 28476 58772 28532
rect 58828 29148 58884 29204
rect 58604 27916 58660 27972
rect 59276 28530 59332 28532
rect 59276 28478 59278 28530
rect 59278 28478 59330 28530
rect 59330 28478 59332 28530
rect 59276 28476 59332 28478
rect 58268 27298 58324 27300
rect 58268 27246 58270 27298
rect 58270 27246 58322 27298
rect 58322 27246 58324 27298
rect 58268 27244 58324 27246
rect 59052 27132 59108 27188
rect 58268 26796 58324 26852
rect 58044 26012 58100 26068
rect 57708 25900 57764 25956
rect 57820 24834 57876 24836
rect 57820 24782 57822 24834
rect 57822 24782 57874 24834
rect 57874 24782 57876 24834
rect 57820 24780 57876 24782
rect 57820 22204 57876 22260
rect 57708 22092 57764 22148
rect 57260 21308 57316 21364
rect 57372 21644 57428 21700
rect 57708 21532 57764 21588
rect 57596 20242 57652 20244
rect 57596 20190 57598 20242
rect 57598 20190 57650 20242
rect 57650 20190 57652 20242
rect 57596 20188 57652 20190
rect 57596 19852 57652 19908
rect 57148 18396 57204 18452
rect 57036 17948 57092 18004
rect 57148 18172 57204 18228
rect 57036 17666 57092 17668
rect 57036 17614 57038 17666
rect 57038 17614 57090 17666
rect 57090 17614 57092 17666
rect 57036 17612 57092 17614
rect 56588 16156 56644 16212
rect 56588 14140 56644 14196
rect 56588 13468 56644 13524
rect 57372 17724 57428 17780
rect 57708 17388 57764 17444
rect 57596 16994 57652 16996
rect 57596 16942 57598 16994
rect 57598 16942 57650 16994
rect 57650 16942 57652 16994
rect 57596 16940 57652 16942
rect 57036 15820 57092 15876
rect 56812 15148 56868 15204
rect 56700 13356 56756 13412
rect 56588 12402 56644 12404
rect 56588 12350 56590 12402
rect 56590 12350 56642 12402
rect 56642 12350 56644 12402
rect 56588 12348 56644 12350
rect 56924 13132 56980 13188
rect 57932 21532 57988 21588
rect 57932 21196 57988 21252
rect 58604 26402 58660 26404
rect 58604 26350 58606 26402
rect 58606 26350 58658 26402
rect 58658 26350 58660 26402
rect 58604 26348 58660 26350
rect 58492 25788 58548 25844
rect 58156 24668 58212 24724
rect 58604 24892 58660 24948
rect 58156 23996 58212 24052
rect 58156 22370 58212 22372
rect 58156 22318 58158 22370
rect 58158 22318 58210 22370
rect 58210 22318 58212 22370
rect 58156 22316 58212 22318
rect 58604 23154 58660 23156
rect 58604 23102 58606 23154
rect 58606 23102 58658 23154
rect 58658 23102 58660 23154
rect 58604 23100 58660 23102
rect 59276 25116 59332 25172
rect 58716 23436 58772 23492
rect 59500 24444 59556 24500
rect 58828 22764 58884 22820
rect 58156 19740 58212 19796
rect 58380 20972 58436 21028
rect 58380 20802 58436 20804
rect 58380 20750 58382 20802
rect 58382 20750 58434 20802
rect 58434 20750 58436 20802
rect 58380 20748 58436 20750
rect 58268 19964 58324 20020
rect 58044 19516 58100 19572
rect 58156 19234 58212 19236
rect 58156 19182 58158 19234
rect 58158 19182 58210 19234
rect 58210 19182 58212 19234
rect 58156 19180 58212 19182
rect 58828 21084 58884 21140
rect 58604 21026 58660 21028
rect 58604 20974 58606 21026
rect 58606 20974 58658 21026
rect 58658 20974 58660 21026
rect 58604 20972 58660 20974
rect 59052 22540 59108 22596
rect 59388 22092 59444 22148
rect 59724 28924 59780 28980
rect 61068 30156 61124 30212
rect 60508 29986 60564 29988
rect 60508 29934 60510 29986
rect 60510 29934 60562 29986
rect 60562 29934 60564 29986
rect 60508 29932 60564 29934
rect 60284 29426 60340 29428
rect 60284 29374 60286 29426
rect 60286 29374 60338 29426
rect 60338 29374 60340 29426
rect 60284 29372 60340 29374
rect 59836 28588 59892 28644
rect 60060 28812 60116 28868
rect 59724 27858 59780 27860
rect 59724 27806 59726 27858
rect 59726 27806 59778 27858
rect 59778 27806 59780 27858
rect 59724 27804 59780 27806
rect 59724 27468 59780 27524
rect 59836 27132 59892 27188
rect 59724 25788 59780 25844
rect 59052 21586 59108 21588
rect 59052 21534 59054 21586
rect 59054 21534 59106 21586
rect 59106 21534 59108 21586
rect 59052 21532 59108 21534
rect 59052 20972 59108 21028
rect 59052 20802 59108 20804
rect 59052 20750 59054 20802
rect 59054 20750 59106 20802
rect 59106 20750 59108 20802
rect 59052 20748 59108 20750
rect 59500 21474 59556 21476
rect 59500 21422 59502 21474
rect 59502 21422 59554 21474
rect 59554 21422 59556 21474
rect 59500 21420 59556 21422
rect 59276 21308 59332 21364
rect 59052 20524 59108 20580
rect 58044 18732 58100 18788
rect 57820 16492 57876 16548
rect 57596 15932 57652 15988
rect 58716 19740 58772 19796
rect 58492 18732 58548 18788
rect 58156 16044 58212 16100
rect 57932 15932 57988 15988
rect 58044 15820 58100 15876
rect 57708 14418 57764 14420
rect 57708 14366 57710 14418
rect 57710 14366 57762 14418
rect 57762 14366 57764 14418
rect 57708 14364 57764 14366
rect 57148 13746 57204 13748
rect 57148 13694 57150 13746
rect 57150 13694 57202 13746
rect 57202 13694 57204 13746
rect 57148 13692 57204 13694
rect 57596 13634 57652 13636
rect 57596 13582 57598 13634
rect 57598 13582 57650 13634
rect 57650 13582 57652 13634
rect 57596 13580 57652 13582
rect 57596 13020 57652 13076
rect 57148 12572 57204 12628
rect 57148 12124 57204 12180
rect 57372 12066 57428 12068
rect 57372 12014 57374 12066
rect 57374 12014 57426 12066
rect 57426 12014 57428 12066
rect 57372 12012 57428 12014
rect 54460 9212 54516 9268
rect 55020 8652 55076 8708
rect 54572 8540 54628 8596
rect 55916 8540 55972 8596
rect 54012 7644 54068 7700
rect 54124 8034 54180 8036
rect 54124 7982 54126 8034
rect 54126 7982 54178 8034
rect 54178 7982 54180 8034
rect 54124 7980 54180 7982
rect 54124 7420 54180 7476
rect 52444 7362 52500 7364
rect 52444 7310 52446 7362
rect 52446 7310 52498 7362
rect 52498 7310 52500 7362
rect 52444 7308 52500 7310
rect 52892 6972 52948 7028
rect 52108 6076 52164 6132
rect 57932 13468 57988 13524
rect 57820 13356 57876 13412
rect 58044 13244 58100 13300
rect 58156 14700 58212 14756
rect 58156 13692 58212 13748
rect 58492 18226 58548 18228
rect 58492 18174 58494 18226
rect 58494 18174 58546 18226
rect 58546 18174 58548 18226
rect 58492 18172 58548 18174
rect 58380 16716 58436 16772
rect 58604 16268 58660 16324
rect 60396 29484 60452 29540
rect 60956 29986 61012 29988
rect 60956 29934 60958 29986
rect 60958 29934 61010 29986
rect 61010 29934 61012 29986
rect 60956 29932 61012 29934
rect 61628 31778 61684 31780
rect 61628 31726 61630 31778
rect 61630 31726 61682 31778
rect 61682 31726 61684 31778
rect 61628 31724 61684 31726
rect 61516 31554 61572 31556
rect 61516 31502 61518 31554
rect 61518 31502 61570 31554
rect 61570 31502 61572 31554
rect 61516 31500 61572 31502
rect 62636 46396 62692 46452
rect 62972 52108 63028 52164
rect 62636 45164 62692 45220
rect 62860 46508 62916 46564
rect 62524 40796 62580 40852
rect 62860 34188 62916 34244
rect 62972 34636 63028 34692
rect 62412 33292 62468 33348
rect 62076 32396 62132 32452
rect 61628 30268 61684 30324
rect 62076 31612 62132 31668
rect 61404 30044 61460 30100
rect 60732 29372 60788 29428
rect 61180 29260 61236 29316
rect 60620 28812 60676 28868
rect 60732 29036 60788 29092
rect 61068 28588 61124 28644
rect 60284 28252 60340 28308
rect 60284 27468 60340 27524
rect 60620 27186 60676 27188
rect 60620 27134 60622 27186
rect 60622 27134 60674 27186
rect 60674 27134 60676 27186
rect 60620 27132 60676 27134
rect 61628 28642 61684 28644
rect 61628 28590 61630 28642
rect 61630 28590 61682 28642
rect 61682 28590 61684 28642
rect 61628 28588 61684 28590
rect 61404 28364 61460 28420
rect 61292 27916 61348 27972
rect 61516 28476 61572 28532
rect 61180 27132 61236 27188
rect 61516 27132 61572 27188
rect 60172 27020 60228 27076
rect 61404 27074 61460 27076
rect 61404 27022 61406 27074
rect 61406 27022 61458 27074
rect 61458 27022 61460 27074
rect 61404 27020 61460 27022
rect 61964 30882 62020 30884
rect 61964 30830 61966 30882
rect 61966 30830 62018 30882
rect 62018 30830 62020 30882
rect 61964 30828 62020 30830
rect 62636 30268 62692 30324
rect 62188 30098 62244 30100
rect 62188 30046 62190 30098
rect 62190 30046 62242 30098
rect 62242 30046 62244 30098
rect 62188 30044 62244 30046
rect 62412 29372 62468 29428
rect 62188 28364 62244 28420
rect 61964 28140 62020 28196
rect 60172 26796 60228 26852
rect 61180 26850 61236 26852
rect 61180 26798 61182 26850
rect 61182 26798 61234 26850
rect 61234 26798 61236 26850
rect 61180 26796 61236 26798
rect 61740 26572 61796 26628
rect 61628 26514 61684 26516
rect 61628 26462 61630 26514
rect 61630 26462 61682 26514
rect 61682 26462 61684 26514
rect 61628 26460 61684 26462
rect 60396 26348 60452 26404
rect 60620 25394 60676 25396
rect 60620 25342 60622 25394
rect 60622 25342 60674 25394
rect 60674 25342 60676 25394
rect 60620 25340 60676 25342
rect 60956 24444 61012 24500
rect 60060 24162 60116 24164
rect 60060 24110 60062 24162
rect 60062 24110 60114 24162
rect 60114 24110 60116 24162
rect 60060 24108 60116 24110
rect 60956 24108 61012 24164
rect 60620 23826 60676 23828
rect 60620 23774 60622 23826
rect 60622 23774 60674 23826
rect 60674 23774 60676 23826
rect 60620 23772 60676 23774
rect 59836 21084 59892 21140
rect 59948 20972 60004 21028
rect 59836 20860 59892 20916
rect 59836 20300 59892 20356
rect 58828 18284 58884 18340
rect 59052 19628 59108 19684
rect 58940 17500 58996 17556
rect 58828 16098 58884 16100
rect 58828 16046 58830 16098
rect 58830 16046 58882 16098
rect 58882 16046 58884 16098
rect 58828 16044 58884 16046
rect 58268 13020 58324 13076
rect 58604 14924 58660 14980
rect 58604 14588 58660 14644
rect 59836 19458 59892 19460
rect 59836 19406 59838 19458
rect 59838 19406 59890 19458
rect 59890 19406 59892 19458
rect 59836 19404 59892 19406
rect 59388 18508 59444 18564
rect 59500 17836 59556 17892
rect 59276 16210 59332 16212
rect 59276 16158 59278 16210
rect 59278 16158 59330 16210
rect 59330 16158 59332 16210
rect 59276 16156 59332 16158
rect 59052 15484 59108 15540
rect 59500 15932 59556 15988
rect 59388 14924 59444 14980
rect 58828 14476 58884 14532
rect 58492 14028 58548 14084
rect 58828 12402 58884 12404
rect 58828 12350 58830 12402
rect 58830 12350 58882 12402
rect 58882 12350 58884 12402
rect 58828 12348 58884 12350
rect 58268 12178 58324 12180
rect 58268 12126 58270 12178
rect 58270 12126 58322 12178
rect 58322 12126 58324 12178
rect 58268 12124 58324 12126
rect 59164 13074 59220 13076
rect 59164 13022 59166 13074
rect 59166 13022 59218 13074
rect 59218 13022 59220 13074
rect 59164 13020 59220 13022
rect 59164 12066 59220 12068
rect 59164 12014 59166 12066
rect 59166 12014 59218 12066
rect 59218 12014 59220 12066
rect 59164 12012 59220 12014
rect 59948 19068 60004 19124
rect 59836 19010 59892 19012
rect 59836 18958 59838 19010
rect 59838 18958 59890 19010
rect 59890 18958 59892 19010
rect 59836 18956 59892 18958
rect 59948 18562 60004 18564
rect 59948 18510 59950 18562
rect 59950 18510 60002 18562
rect 60002 18510 60004 18562
rect 59948 18508 60004 18510
rect 59836 18396 59892 18452
rect 60620 22594 60676 22596
rect 60620 22542 60622 22594
rect 60622 22542 60674 22594
rect 60674 22542 60676 22594
rect 60620 22540 60676 22542
rect 60956 23266 61012 23268
rect 60956 23214 60958 23266
rect 60958 23214 61010 23266
rect 61010 23214 61012 23266
rect 60956 23212 61012 23214
rect 61180 23100 61236 23156
rect 60508 21756 60564 21812
rect 60396 21532 60452 21588
rect 60172 21362 60228 21364
rect 60172 21310 60174 21362
rect 60174 21310 60226 21362
rect 60226 21310 60228 21362
rect 60172 21308 60228 21310
rect 60060 18396 60116 18452
rect 60172 21084 60228 21140
rect 59836 16492 59892 16548
rect 60284 20076 60340 20132
rect 60284 18956 60340 19012
rect 60172 17052 60228 17108
rect 60620 20860 60676 20916
rect 60508 20636 60564 20692
rect 60508 19180 60564 19236
rect 60732 20802 60788 20804
rect 60732 20750 60734 20802
rect 60734 20750 60786 20802
rect 60786 20750 60788 20802
rect 60732 20748 60788 20750
rect 61516 24108 61572 24164
rect 61292 21308 61348 21364
rect 60956 20748 61012 20804
rect 61068 20578 61124 20580
rect 61068 20526 61070 20578
rect 61070 20526 61122 20578
rect 61122 20526 61124 20578
rect 61068 20524 61124 20526
rect 61180 20412 61236 20468
rect 60508 18732 60564 18788
rect 60844 18674 60900 18676
rect 60844 18622 60846 18674
rect 60846 18622 60898 18674
rect 60898 18622 60900 18674
rect 60844 18620 60900 18622
rect 61404 20188 61460 20244
rect 61628 21026 61684 21028
rect 61628 20974 61630 21026
rect 61630 20974 61682 21026
rect 61682 20974 61684 21026
rect 61628 20972 61684 20974
rect 61404 20018 61460 20020
rect 61404 19966 61406 20018
rect 61406 19966 61458 20018
rect 61458 19966 61460 20018
rect 61404 19964 61460 19966
rect 62076 27580 62132 27636
rect 62188 27186 62244 27188
rect 62188 27134 62190 27186
rect 62190 27134 62242 27186
rect 62242 27134 62244 27186
rect 62188 27132 62244 27134
rect 62188 26402 62244 26404
rect 62188 26350 62190 26402
rect 62190 26350 62242 26402
rect 62242 26350 62244 26402
rect 62188 26348 62244 26350
rect 62188 21980 62244 22036
rect 61964 20860 62020 20916
rect 62076 20300 62132 20356
rect 61964 19852 62020 19908
rect 61628 19180 61684 19236
rect 61404 19122 61460 19124
rect 61404 19070 61406 19122
rect 61406 19070 61458 19122
rect 61458 19070 61460 19122
rect 61404 19068 61460 19070
rect 61404 18844 61460 18900
rect 61628 18956 61684 19012
rect 60620 17890 60676 17892
rect 60620 17838 60622 17890
rect 60622 17838 60674 17890
rect 60674 17838 60676 17890
rect 60620 17836 60676 17838
rect 60508 17724 60564 17780
rect 60732 17724 60788 17780
rect 60844 17500 60900 17556
rect 61292 18284 61348 18340
rect 61404 17388 61460 17444
rect 60620 16716 60676 16772
rect 61180 16380 61236 16436
rect 61068 15874 61124 15876
rect 61068 15822 61070 15874
rect 61070 15822 61122 15874
rect 61122 15822 61124 15874
rect 61068 15820 61124 15822
rect 60396 15538 60452 15540
rect 60396 15486 60398 15538
rect 60398 15486 60450 15538
rect 60450 15486 60452 15538
rect 60396 15484 60452 15486
rect 60844 15538 60900 15540
rect 60844 15486 60846 15538
rect 60846 15486 60898 15538
rect 60898 15486 60900 15538
rect 60844 15484 60900 15486
rect 61068 14700 61124 14756
rect 60620 14530 60676 14532
rect 60620 14478 60622 14530
rect 60622 14478 60674 14530
rect 60674 14478 60676 14530
rect 60620 14476 60676 14478
rect 61068 14364 61124 14420
rect 59612 13916 59668 13972
rect 60284 13970 60340 13972
rect 60284 13918 60286 13970
rect 60286 13918 60338 13970
rect 60338 13918 60340 13970
rect 60284 13916 60340 13918
rect 61628 17724 61684 17780
rect 61516 16492 61572 16548
rect 61404 15538 61460 15540
rect 61404 15486 61406 15538
rect 61406 15486 61458 15538
rect 61458 15486 61460 15538
rect 61404 15484 61460 15486
rect 61852 19516 61908 19572
rect 62188 18732 62244 18788
rect 61852 18284 61908 18340
rect 62076 18450 62132 18452
rect 62076 18398 62078 18450
rect 62078 18398 62130 18450
rect 62130 18398 62132 18450
rect 62076 18396 62132 18398
rect 61852 17666 61908 17668
rect 61852 17614 61854 17666
rect 61854 17614 61906 17666
rect 61906 17614 61908 17666
rect 61852 17612 61908 17614
rect 62076 17442 62132 17444
rect 62076 17390 62078 17442
rect 62078 17390 62130 17442
rect 62130 17390 62132 17442
rect 62076 17388 62132 17390
rect 61852 16604 61908 16660
rect 61964 16940 62020 16996
rect 61292 14588 61348 14644
rect 61628 14642 61684 14644
rect 61628 14590 61630 14642
rect 61630 14590 61682 14642
rect 61682 14590 61684 14642
rect 61628 14588 61684 14590
rect 60732 13858 60788 13860
rect 60732 13806 60734 13858
rect 60734 13806 60786 13858
rect 60786 13806 60788 13858
rect 60732 13804 60788 13806
rect 59836 13746 59892 13748
rect 59836 13694 59838 13746
rect 59838 13694 59890 13746
rect 59890 13694 59892 13746
rect 59836 13692 59892 13694
rect 59500 12796 59556 12852
rect 61964 16210 62020 16212
rect 61964 16158 61966 16210
rect 61966 16158 62018 16210
rect 62018 16158 62020 16210
rect 61964 16156 62020 16158
rect 62188 17106 62244 17108
rect 62188 17054 62190 17106
rect 62190 17054 62242 17106
rect 62242 17054 62244 17106
rect 62188 17052 62244 17054
rect 62188 15538 62244 15540
rect 62188 15486 62190 15538
rect 62190 15486 62242 15538
rect 62242 15486 62244 15538
rect 62188 15484 62244 15486
rect 62524 25900 62580 25956
rect 62524 16716 62580 16772
rect 62972 30268 63028 30324
rect 62860 29932 62916 29988
rect 62860 19404 62916 19460
rect 62972 27580 63028 27636
rect 62972 17724 63028 17780
rect 62636 15484 62692 15540
rect 62412 14700 62468 14756
rect 61180 12348 61236 12404
rect 59276 11676 59332 11732
rect 57148 10834 57204 10836
rect 57148 10782 57150 10834
rect 57150 10782 57202 10834
rect 57202 10782 57204 10834
rect 57148 10780 57204 10782
rect 56700 7980 56756 8036
rect 56364 4508 56420 4564
rect 51772 3276 51828 3332
rect 46396 3164 46452 3220
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 11442 60508 11452 60564
rect 11508 60508 25340 60564
rect 25396 60508 25406 60564
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 16146 60172 16156 60228
rect 16212 60172 17948 60228
rect 18004 60172 18014 60228
rect 47730 60172 47740 60228
rect 47796 60172 48972 60228
rect 49028 60172 49038 60228
rect 29586 59948 29596 60004
rect 29652 59948 33964 60004
rect 34020 59948 34972 60004
rect 35028 59948 35038 60004
rect 13570 59836 13580 59892
rect 13636 59836 14028 59892
rect 14084 59836 19964 59892
rect 20020 59836 20860 59892
rect 20916 59836 20926 59892
rect 22530 59836 22540 59892
rect 22596 59836 23212 59892
rect 23268 59836 27356 59892
rect 27412 59836 27422 59892
rect 29698 59836 29708 59892
rect 29764 59836 31164 59892
rect 31220 59836 32732 59892
rect 32788 59836 33068 59892
rect 33124 59836 33134 59892
rect 20290 59724 20300 59780
rect 20356 59724 28140 59780
rect 28196 59724 28206 59780
rect 30034 59724 30044 59780
rect 30100 59724 32396 59780
rect 32452 59724 33180 59780
rect 33236 59724 33246 59780
rect 22082 59612 22092 59668
rect 22148 59612 25228 59668
rect 25284 59612 26348 59668
rect 26404 59612 26414 59668
rect 29138 59612 29148 59668
rect 29204 59612 33740 59668
rect 33796 59612 33806 59668
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 14802 59388 14812 59444
rect 14868 59388 16156 59444
rect 16212 59388 16222 59444
rect 26226 59388 26236 59444
rect 26292 59388 27468 59444
rect 27524 59388 27534 59444
rect 48402 59388 48412 59444
rect 48468 59388 49756 59444
rect 49812 59388 49822 59444
rect 14130 59276 14140 59332
rect 14196 59276 14924 59332
rect 14980 59276 17948 59332
rect 18004 59276 18014 59332
rect 29810 59276 29820 59332
rect 29876 59276 34188 59332
rect 34244 59276 34748 59332
rect 34804 59276 34814 59332
rect 20850 59164 20860 59220
rect 20916 59164 23660 59220
rect 23716 59164 23726 59220
rect 24546 59164 24556 59220
rect 24612 59164 25004 59220
rect 25060 59164 25564 59220
rect 25620 59164 25630 59220
rect 27794 59164 27804 59220
rect 27860 59164 32284 59220
rect 32340 59164 32350 59220
rect 16258 59052 16268 59108
rect 16324 59052 21756 59108
rect 21812 59052 21822 59108
rect 27906 59052 27916 59108
rect 27972 59052 29820 59108
rect 29876 59052 29886 59108
rect 34066 59052 34076 59108
rect 34132 59052 35532 59108
rect 35588 59052 35598 59108
rect 12898 58940 12908 58996
rect 12964 58940 13804 58996
rect 13860 58940 13870 58996
rect 21410 58940 21420 58996
rect 21476 58940 23436 58996
rect 23492 58940 23502 58996
rect 26114 58940 26124 58996
rect 26180 58940 26796 58996
rect 26852 58940 27804 58996
rect 27860 58940 27870 58996
rect 31154 58940 31164 58996
rect 31220 58940 32172 58996
rect 32228 58940 33180 58996
rect 33236 58940 33246 58996
rect 15092 58828 15260 58884
rect 15316 58828 19516 58884
rect 19572 58828 19582 58884
rect 20962 58828 20972 58884
rect 21028 58828 23884 58884
rect 23940 58828 23950 58884
rect 24546 58828 24556 58884
rect 24612 58828 30268 58884
rect 30324 58828 30334 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 15092 58772 15148 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 13794 58716 13804 58772
rect 13860 58716 15148 58772
rect 28354 58716 28364 58772
rect 28420 58716 29148 58772
rect 29204 58716 29214 58772
rect 29586 58716 29596 58772
rect 29652 58716 30380 58772
rect 30436 58716 31276 58772
rect 31332 58716 31342 58772
rect 32610 58716 32620 58772
rect 32676 58716 33516 58772
rect 33572 58716 33582 58772
rect 13458 58604 13468 58660
rect 13524 58604 15932 58660
rect 15988 58604 15998 58660
rect 28018 58604 28028 58660
rect 28084 58604 29484 58660
rect 29540 58604 29550 58660
rect 63200 58548 64000 58576
rect 14466 58492 14476 58548
rect 14532 58492 15820 58548
rect 15876 58492 15886 58548
rect 20066 58492 20076 58548
rect 20132 58492 21980 58548
rect 22036 58492 23884 58548
rect 23940 58492 25004 58548
rect 25060 58492 25070 58548
rect 48066 58492 48076 58548
rect 48132 58492 51660 58548
rect 51716 58492 52108 58548
rect 52164 58492 52174 58548
rect 62178 58492 62188 58548
rect 62244 58492 64000 58548
rect 63200 58464 64000 58492
rect 14130 58380 14140 58436
rect 14196 58380 15372 58436
rect 15428 58380 16044 58436
rect 16100 58380 19628 58436
rect 19684 58380 19694 58436
rect 26852 58380 27020 58436
rect 27076 58380 27086 58436
rect 27794 58380 27804 58436
rect 27860 58380 28588 58436
rect 28644 58380 29596 58436
rect 29652 58380 29662 58436
rect 30146 58380 30156 58436
rect 30212 58380 32172 58436
rect 32228 58380 32508 58436
rect 32564 58380 32574 58436
rect 43698 58380 43708 58436
rect 43764 58380 50316 58436
rect 50372 58380 51324 58436
rect 51380 58380 51390 58436
rect 26852 58212 26908 58380
rect 47506 58268 47516 58324
rect 47572 58268 50764 58324
rect 50820 58268 51548 58324
rect 51604 58268 51614 58324
rect 14802 58156 14812 58212
rect 14868 58156 15484 58212
rect 15540 58156 15550 58212
rect 16930 58156 16940 58212
rect 16996 58156 24668 58212
rect 24724 58156 26908 58212
rect 28802 58156 28812 58212
rect 28868 58156 36092 58212
rect 36148 58156 40012 58212
rect 40068 58156 40684 58212
rect 40740 58156 41132 58212
rect 41188 58156 41198 58212
rect 44482 58156 44492 58212
rect 44548 58156 45612 58212
rect 45668 58156 46060 58212
rect 46116 58156 46126 58212
rect 48066 58156 48076 58212
rect 48132 58156 48524 58212
rect 48580 58156 49196 58212
rect 49252 58156 49262 58212
rect 50372 58156 51324 58212
rect 51380 58156 51660 58212
rect 51716 58156 51726 58212
rect 50372 58100 50428 58156
rect 18834 58044 18844 58100
rect 18900 58044 19628 58100
rect 19684 58044 19694 58100
rect 21522 58044 21532 58100
rect 21588 58044 26460 58100
rect 26516 58044 26526 58100
rect 40226 58044 40236 58100
rect 40292 58044 48972 58100
rect 49028 58044 50428 58100
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 16370 57932 16380 57988
rect 16436 57932 17164 57988
rect 17220 57932 19180 57988
rect 19236 57932 19246 57988
rect 25106 57932 25116 57988
rect 25172 57932 37100 57988
rect 37156 57932 48412 57988
rect 48468 57932 48478 57988
rect 19180 57876 19236 57932
rect 13570 57820 13580 57876
rect 13636 57820 14588 57876
rect 14644 57820 14654 57876
rect 15474 57820 15484 57876
rect 15540 57820 18844 57876
rect 18900 57820 18910 57876
rect 19180 57820 19964 57876
rect 20020 57820 20030 57876
rect 28466 57820 28476 57876
rect 28532 57820 39564 57876
rect 39620 57820 39630 57876
rect 40562 57820 40572 57876
rect 40628 57820 42252 57876
rect 42308 57820 55356 57876
rect 55412 57820 56700 57876
rect 56756 57820 56766 57876
rect 14028 57708 16940 57764
rect 16996 57708 17006 57764
rect 17938 57708 17948 57764
rect 18004 57708 19404 57764
rect 19460 57708 19470 57764
rect 19730 57708 19740 57764
rect 19796 57708 21196 57764
rect 21252 57708 21262 57764
rect 24322 57708 24332 57764
rect 24388 57708 28028 57764
rect 28084 57708 28094 57764
rect 36418 57708 36428 57764
rect 36484 57708 48076 57764
rect 48132 57708 48142 57764
rect 52098 57708 52108 57764
rect 52164 57708 53788 57764
rect 53844 57708 55916 57764
rect 55972 57708 55982 57764
rect 14028 57540 14084 57708
rect 15026 57596 15036 57652
rect 15092 57540 15148 57652
rect 15922 57596 15932 57652
rect 15988 57596 21868 57652
rect 21924 57596 21934 57652
rect 22082 57596 22092 57652
rect 22148 57596 24108 57652
rect 24164 57596 24174 57652
rect 24994 57596 25004 57652
rect 25060 57596 26012 57652
rect 26068 57596 26078 57652
rect 29250 57596 29260 57652
rect 29316 57596 30156 57652
rect 30212 57596 30222 57652
rect 32834 57596 32844 57652
rect 32900 57596 33740 57652
rect 33796 57596 33806 57652
rect 47954 57596 47964 57652
rect 48020 57596 48860 57652
rect 48916 57596 48926 57652
rect 51874 57596 51884 57652
rect 51940 57596 52892 57652
rect 52948 57596 52958 57652
rect 53218 57596 53228 57652
rect 53284 57596 54012 57652
rect 54068 57596 54078 57652
rect 14018 57484 14028 57540
rect 14084 57484 14094 57540
rect 15092 57484 19292 57540
rect 19348 57484 19358 57540
rect 19618 57484 19628 57540
rect 19684 57484 20748 57540
rect 20804 57484 28476 57540
rect 28532 57484 28542 57540
rect 29474 57484 29484 57540
rect 29540 57484 37324 57540
rect 37380 57484 37390 57540
rect 37986 57484 37996 57540
rect 38052 57484 41244 57540
rect 41300 57484 47628 57540
rect 47684 57484 47694 57540
rect 50372 57484 52780 57540
rect 52836 57484 52846 57540
rect 55010 57484 55020 57540
rect 55076 57484 55468 57540
rect 55524 57484 55534 57540
rect 19628 57428 19684 57484
rect 50372 57428 50428 57484
rect 12114 57372 12124 57428
rect 12180 57372 12684 57428
rect 12740 57372 19684 57428
rect 23202 57372 23212 57428
rect 23268 57372 24108 57428
rect 24164 57372 24780 57428
rect 24836 57372 24846 57428
rect 46610 57372 46620 57428
rect 46676 57372 50428 57428
rect 52322 57372 52332 57428
rect 52388 57372 53564 57428
rect 53620 57372 53630 57428
rect 19394 57260 19404 57316
rect 19460 57260 20524 57316
rect 20580 57260 20590 57316
rect 24658 57260 24668 57316
rect 24724 57260 26460 57316
rect 26516 57260 26526 57316
rect 44034 57260 44044 57316
rect 44100 57260 44940 57316
rect 44996 57260 47068 57316
rect 47124 57260 47134 57316
rect 51090 57260 51100 57316
rect 51156 57260 53116 57316
rect 53172 57260 53676 57316
rect 53732 57260 53742 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 10098 57148 10108 57204
rect 10164 57148 16156 57204
rect 16212 57148 16222 57204
rect 17826 57148 17836 57204
rect 17892 57148 22092 57204
rect 22148 57148 22158 57204
rect 24434 57148 24444 57204
rect 24500 57148 28476 57204
rect 28532 57148 29148 57204
rect 29204 57148 29214 57204
rect 29810 57148 29820 57204
rect 29876 57148 32732 57204
rect 32788 57148 32798 57204
rect 38434 57148 38444 57204
rect 38500 57148 54852 57204
rect 20524 57092 20580 57148
rect 13132 57036 14028 57092
rect 14084 57036 14094 57092
rect 15586 57036 15596 57092
rect 15652 57036 18508 57092
rect 18564 57036 18574 57092
rect 20524 57036 20636 57092
rect 20692 57036 20702 57092
rect 20962 57036 20972 57092
rect 21028 57036 25228 57092
rect 25284 57036 25294 57092
rect 13132 56980 13188 57036
rect 54796 56980 54852 57148
rect 55010 57036 55020 57092
rect 55076 57036 55804 57092
rect 55860 57036 56364 57092
rect 56420 57036 56430 57092
rect 5730 56924 5740 56980
rect 5796 56924 13132 56980
rect 13188 56924 13198 56980
rect 13906 56924 13916 56980
rect 13972 56924 15036 56980
rect 15092 56924 16492 56980
rect 16548 56924 18172 56980
rect 18228 56924 18238 56980
rect 23538 56924 23548 56980
rect 23604 56924 25676 56980
rect 25732 56924 27692 56980
rect 27748 56924 27758 56980
rect 39554 56924 39564 56980
rect 39620 56924 40908 56980
rect 40964 56924 41356 56980
rect 41412 56924 41422 56980
rect 54796 56924 56924 56980
rect 56980 56924 57820 56980
rect 57876 56924 57886 56980
rect 13010 56812 13020 56868
rect 13076 56812 13580 56868
rect 13636 56812 18340 56868
rect 18498 56812 18508 56868
rect 18564 56812 20188 56868
rect 20244 56812 21644 56868
rect 21700 56812 21710 56868
rect 23986 56812 23996 56868
rect 24052 56812 27020 56868
rect 27076 56812 27580 56868
rect 27636 56812 27646 56868
rect 45164 56812 50428 56868
rect 54786 56812 54796 56868
rect 54852 56812 55692 56868
rect 55748 56812 57036 56868
rect 57092 56812 57102 56868
rect 18284 56756 18340 56812
rect 45164 56756 45220 56812
rect 50372 56756 50428 56812
rect 14690 56700 14700 56756
rect 14756 56700 17052 56756
rect 17108 56700 17118 56756
rect 18284 56700 19012 56756
rect 19170 56700 19180 56756
rect 19236 56700 19740 56756
rect 19796 56700 23660 56756
rect 23716 56700 23726 56756
rect 23884 56700 24556 56756
rect 24612 56700 25116 56756
rect 25172 56700 25182 56756
rect 31378 56700 31388 56756
rect 31444 56700 32060 56756
rect 32116 56700 32126 56756
rect 37090 56700 37100 56756
rect 37156 56700 39340 56756
rect 39396 56700 40236 56756
rect 40292 56700 40302 56756
rect 40450 56700 40460 56756
rect 40516 56700 42252 56756
rect 42308 56700 42318 56756
rect 45154 56700 45164 56756
rect 45220 56700 45230 56756
rect 45826 56700 45836 56756
rect 45892 56700 46508 56756
rect 46564 56700 47628 56756
rect 47684 56700 47694 56756
rect 50372 56700 57260 56756
rect 57316 56700 58268 56756
rect 58324 56700 59052 56756
rect 59108 56700 59118 56756
rect 18956 56644 19012 56700
rect 23884 56644 23940 56700
rect 15362 56588 15372 56644
rect 15428 56588 18284 56644
rect 18340 56588 18350 56644
rect 18956 56588 22764 56644
rect 22820 56588 23940 56644
rect 24434 56588 24444 56644
rect 24500 56588 30492 56644
rect 30548 56588 30558 56644
rect 31266 56588 31276 56644
rect 31332 56588 32396 56644
rect 32452 56588 32462 56644
rect 33058 56588 33068 56644
rect 33124 56588 34524 56644
rect 34580 56588 39004 56644
rect 39060 56588 39070 56644
rect 44258 56588 44268 56644
rect 44324 56588 46172 56644
rect 46228 56588 46238 56644
rect 52854 56588 52892 56644
rect 52948 56588 52958 56644
rect 54898 56588 54908 56644
rect 54964 56588 55468 56644
rect 55524 56588 56476 56644
rect 56532 56588 56542 56644
rect 33068 56532 33124 56588
rect 14130 56476 14140 56532
rect 14196 56476 15708 56532
rect 15764 56476 16828 56532
rect 16884 56476 16894 56532
rect 29698 56476 29708 56532
rect 29764 56476 31052 56532
rect 31108 56476 31118 56532
rect 31602 56476 31612 56532
rect 31668 56476 33124 56532
rect 34178 56476 34188 56532
rect 34244 56476 37772 56532
rect 37828 56476 37838 56532
rect 44706 56476 44716 56532
rect 44772 56476 45500 56532
rect 45556 56476 45948 56532
rect 46004 56476 50092 56532
rect 50148 56476 50158 56532
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 20178 56364 20188 56420
rect 20244 56364 24332 56420
rect 24388 56364 28812 56420
rect 28868 56364 28878 56420
rect 30706 56364 30716 56420
rect 30772 56364 31276 56420
rect 31332 56364 33964 56420
rect 34020 56364 34030 56420
rect 34626 56364 34636 56420
rect 34692 56364 38556 56420
rect 38612 56364 38622 56420
rect 14354 56252 14364 56308
rect 14420 56252 15596 56308
rect 15652 56252 15662 56308
rect 18946 56252 18956 56308
rect 19012 56252 21196 56308
rect 21252 56252 21262 56308
rect 25666 56252 25676 56308
rect 25732 56252 28588 56308
rect 28644 56252 28654 56308
rect 29138 56252 29148 56308
rect 29204 56252 38668 56308
rect 42578 56252 42588 56308
rect 42644 56252 42812 56308
rect 42868 56252 49084 56308
rect 49140 56252 49756 56308
rect 49812 56252 49822 56308
rect 50082 56252 50092 56308
rect 50148 56252 50316 56308
rect 50372 56252 50382 56308
rect 51650 56252 51660 56308
rect 51716 56252 53788 56308
rect 53844 56252 54796 56308
rect 54852 56252 54862 56308
rect 56802 56252 56812 56308
rect 56868 56252 58380 56308
rect 58436 56252 59276 56308
rect 59332 56252 59342 56308
rect 38612 56196 38668 56252
rect 50092 56196 50148 56252
rect 12562 56140 12572 56196
rect 12628 56140 20188 56196
rect 20244 56140 20254 56196
rect 20514 56140 20524 56196
rect 20580 56140 23548 56196
rect 23604 56140 23614 56196
rect 24210 56140 24220 56196
rect 24276 56140 25564 56196
rect 25620 56140 29596 56196
rect 29652 56140 29662 56196
rect 30594 56140 30604 56196
rect 30660 56140 32172 56196
rect 32228 56140 32238 56196
rect 38612 56140 40460 56196
rect 40516 56140 40526 56196
rect 48066 56140 48076 56196
rect 48132 56140 50148 56196
rect 55570 56140 55580 56196
rect 55636 56140 57820 56196
rect 57876 56140 57886 56196
rect 15922 56028 15932 56084
rect 15988 56028 16716 56084
rect 16772 56028 18508 56084
rect 18564 56028 18574 56084
rect 23090 56028 23100 56084
rect 23156 56028 25900 56084
rect 25956 56028 25966 56084
rect 29922 56028 29932 56084
rect 29988 56028 31948 56084
rect 32004 56028 32014 56084
rect 35410 56028 35420 56084
rect 35476 56028 36092 56084
rect 36148 56028 37100 56084
rect 37156 56028 37166 56084
rect 48178 56028 48188 56084
rect 48244 56028 48972 56084
rect 49028 56028 49038 56084
rect 49746 56028 49756 56084
rect 49812 56028 50988 56084
rect 51044 56028 51054 56084
rect 49756 55972 49812 56028
rect 12562 55916 12572 55972
rect 12628 55916 13356 55972
rect 13412 55916 13422 55972
rect 14690 55916 14700 55972
rect 14756 55916 15148 55972
rect 24434 55916 24444 55972
rect 24500 55916 24892 55972
rect 24948 55916 27860 55972
rect 32162 55916 32172 55972
rect 32228 55916 33292 55972
rect 33348 55916 37660 55972
rect 37716 55916 38332 55972
rect 38388 55916 38668 55972
rect 38994 55916 39004 55972
rect 39060 55916 39452 55972
rect 39508 55916 40460 55972
rect 40516 55916 40526 55972
rect 41458 55916 41468 55972
rect 41524 55916 43596 55972
rect 43652 55916 43662 55972
rect 46834 55916 46844 55972
rect 46900 55916 49812 55972
rect 15092 55860 15148 55916
rect 15092 55804 16156 55860
rect 16212 55804 16222 55860
rect 24322 55804 24332 55860
rect 24388 55804 27468 55860
rect 27524 55804 27534 55860
rect 27804 55748 27860 55916
rect 33068 55804 35588 55860
rect 27794 55692 27804 55748
rect 27860 55692 28140 55748
rect 28196 55692 28206 55748
rect 30818 55692 30828 55748
rect 30884 55692 32732 55748
rect 32788 55692 32798 55748
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 33068 55636 33124 55804
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 35532 55636 35588 55804
rect 38612 55748 38668 55916
rect 38612 55692 39004 55748
rect 39060 55692 39070 55748
rect 41010 55692 41020 55748
rect 41076 55692 42252 55748
rect 42308 55692 46900 55748
rect 47618 55692 47628 55748
rect 47684 55692 48636 55748
rect 48692 55692 49420 55748
rect 49476 55692 49486 55748
rect 46844 55636 46900 55692
rect 17266 55580 17276 55636
rect 17332 55580 22652 55636
rect 22708 55580 22718 55636
rect 27570 55580 27580 55636
rect 27636 55580 33124 55636
rect 35532 55580 38892 55636
rect 38948 55580 38958 55636
rect 45042 55580 45052 55636
rect 45108 55580 46620 55636
rect 46676 55580 46686 55636
rect 46844 55580 52220 55636
rect 52276 55580 57260 55636
rect 57316 55580 57326 55636
rect 11666 55468 11676 55524
rect 11732 55468 14252 55524
rect 14308 55468 14588 55524
rect 14644 55468 14654 55524
rect 17938 55468 17948 55524
rect 18004 55468 18014 55524
rect 18274 55468 18284 55524
rect 18340 55468 20188 55524
rect 20244 55468 20254 55524
rect 27906 55468 27916 55524
rect 27972 55468 30716 55524
rect 30772 55468 30782 55524
rect 31042 55468 31052 55524
rect 31108 55468 31500 55524
rect 31556 55468 31566 55524
rect 32610 55468 32620 55524
rect 32676 55468 35308 55524
rect 35364 55468 36876 55524
rect 36932 55468 36942 55524
rect 41010 55468 41020 55524
rect 41076 55468 55132 55524
rect 55188 55468 55198 55524
rect 56130 55468 56140 55524
rect 56196 55468 56476 55524
rect 56532 55468 56542 55524
rect 17948 55412 18004 55468
rect 15250 55356 15260 55412
rect 15316 55356 15484 55412
rect 15540 55356 19516 55412
rect 19572 55356 19582 55412
rect 23734 55356 23772 55412
rect 23828 55356 23838 55412
rect 25330 55356 25340 55412
rect 25396 55356 26572 55412
rect 26628 55356 26638 55412
rect 27356 55356 27468 55412
rect 27524 55356 28252 55412
rect 28308 55356 28318 55412
rect 30146 55356 30156 55412
rect 30212 55356 33068 55412
rect 33124 55356 33134 55412
rect 33282 55356 33292 55412
rect 33348 55356 35644 55412
rect 35700 55356 37212 55412
rect 37268 55356 37278 55412
rect 45378 55356 45388 55412
rect 45444 55356 46172 55412
rect 46228 55356 46238 55412
rect 47730 55356 47740 55412
rect 47796 55356 50540 55412
rect 50596 55356 50988 55412
rect 51044 55356 51436 55412
rect 51492 55356 51502 55412
rect 55458 55356 55468 55412
rect 55524 55356 56812 55412
rect 56868 55356 56878 55412
rect 18722 55244 18732 55300
rect 18788 55244 21868 55300
rect 21924 55244 22764 55300
rect 22820 55244 22830 55300
rect 23874 55244 23884 55300
rect 23940 55244 24780 55300
rect 24836 55244 27132 55300
rect 27188 55244 27198 55300
rect 27356 55188 27412 55356
rect 30706 55244 30716 55300
rect 30772 55244 32620 55300
rect 32676 55244 33180 55300
rect 33236 55244 33246 55300
rect 36306 55244 36316 55300
rect 36372 55244 36652 55300
rect 36708 55244 36988 55300
rect 37044 55244 37054 55300
rect 37762 55244 37772 55300
rect 37828 55244 39676 55300
rect 39732 55244 39742 55300
rect 40786 55244 40796 55300
rect 40852 55244 42588 55300
rect 42644 55244 42654 55300
rect 47954 55244 47964 55300
rect 48020 55244 49868 55300
rect 49924 55244 49934 55300
rect 53218 55244 53228 55300
rect 53284 55244 53900 55300
rect 53956 55244 53966 55300
rect 58146 55244 58156 55300
rect 58212 55244 62748 55300
rect 62804 55244 62814 55300
rect 12674 55132 12684 55188
rect 12740 55132 14140 55188
rect 14196 55132 14206 55188
rect 15474 55132 15484 55188
rect 15540 55132 16268 55188
rect 16324 55132 18620 55188
rect 18676 55132 18686 55188
rect 19730 55132 19740 55188
rect 19796 55132 20860 55188
rect 20916 55132 20926 55188
rect 22978 55132 22988 55188
rect 23044 55132 24220 55188
rect 24276 55132 26684 55188
rect 26740 55132 27412 55188
rect 28028 55132 31948 55188
rect 32004 55132 33740 55188
rect 33796 55132 33806 55188
rect 33954 55132 33964 55188
rect 34020 55132 37324 55188
rect 37380 55132 37390 55188
rect 42914 55132 42924 55188
rect 42980 55132 44716 55188
rect 44772 55132 44782 55188
rect 46498 55132 46508 55188
rect 46564 55132 49196 55188
rect 49252 55132 49262 55188
rect 55906 55132 55916 55188
rect 55972 55132 58716 55188
rect 58772 55132 58782 55188
rect 59378 55132 59388 55188
rect 59444 55132 61068 55188
rect 61124 55132 61134 55188
rect 28028 55076 28084 55132
rect 1698 55020 1708 55076
rect 1764 55020 2492 55076
rect 2548 55020 2558 55076
rect 8642 55020 8652 55076
rect 8708 55020 10556 55076
rect 10612 55020 11004 55076
rect 11060 55020 11070 55076
rect 11778 55020 11788 55076
rect 11844 55020 12348 55076
rect 12404 55020 12414 55076
rect 13906 55020 13916 55076
rect 13972 55020 17668 55076
rect 18162 55020 18172 55076
rect 18228 55020 21980 55076
rect 22036 55020 22046 55076
rect 23090 55020 23100 55076
rect 23156 55020 25452 55076
rect 25508 55020 25676 55076
rect 25732 55020 25742 55076
rect 26898 55020 26908 55076
rect 26964 55020 28084 55076
rect 28242 55020 28252 55076
rect 28308 55020 30604 55076
rect 30660 55020 30670 55076
rect 35858 55020 35868 55076
rect 35924 55020 37996 55076
rect 38052 55020 38062 55076
rect 43894 55020 43932 55076
rect 43988 55020 43998 55076
rect 47142 55020 47180 55076
rect 47236 55020 47246 55076
rect 47394 55020 47404 55076
rect 47460 55020 49588 55076
rect 50082 55020 50092 55076
rect 50148 55020 50876 55076
rect 50932 55020 50942 55076
rect 51174 55020 51212 55076
rect 51268 55020 51278 55076
rect 51986 55020 51996 55076
rect 52052 55020 53452 55076
rect 53508 55020 53518 55076
rect 53666 55020 53676 55076
rect 53732 55020 56924 55076
rect 56980 55020 56990 55076
rect 11004 54964 11060 55020
rect 11004 54908 15932 54964
rect 15988 54908 17388 54964
rect 17444 54908 17454 54964
rect 17612 54852 17668 55020
rect 22082 54908 22092 54964
rect 22148 54908 25228 54964
rect 25284 54908 25294 54964
rect 36418 54908 36428 54964
rect 36484 54908 36764 54964
rect 36820 54908 38892 54964
rect 38948 54908 38958 54964
rect 45042 54908 45052 54964
rect 45108 54908 46396 54964
rect 46452 54908 46462 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 9538 54796 9548 54852
rect 9604 54796 11228 54852
rect 11284 54796 13916 54852
rect 13972 54796 13982 54852
rect 17612 54796 18060 54852
rect 18116 54796 18126 54852
rect 18274 54796 18284 54852
rect 18340 54796 19684 54852
rect 19628 54740 19684 54796
rect 30604 54796 32508 54852
rect 32564 54796 32574 54852
rect 46274 54796 46284 54852
rect 46340 54796 48972 54852
rect 49028 54796 49308 54852
rect 49364 54796 49374 54852
rect 13234 54684 13244 54740
rect 13300 54684 18508 54740
rect 18564 54684 19180 54740
rect 19236 54684 19246 54740
rect 19628 54684 22204 54740
rect 22260 54684 23212 54740
rect 23268 54684 23278 54740
rect 29474 54684 29484 54740
rect 29540 54684 30156 54740
rect 30212 54684 30222 54740
rect 30604 54628 30660 54796
rect 49532 54740 49588 55020
rect 51650 54908 51660 54964
rect 51716 54908 53564 54964
rect 53620 54908 53630 54964
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 56018 54796 56028 54852
rect 56084 54796 57596 54852
rect 57652 54796 57662 54852
rect 34514 54684 34524 54740
rect 34580 54684 36540 54740
rect 36596 54684 36606 54740
rect 42242 54684 42252 54740
rect 42308 54684 45892 54740
rect 49532 54684 50428 54740
rect 50866 54684 50876 54740
rect 50932 54684 52668 54740
rect 52724 54684 52734 54740
rect 55682 54684 55692 54740
rect 55748 54684 56588 54740
rect 56644 54684 56654 54740
rect 45836 54628 45892 54684
rect 9986 54572 9996 54628
rect 10052 54572 11676 54628
rect 11732 54572 12852 54628
rect 13010 54572 13020 54628
rect 13076 54572 13804 54628
rect 13860 54572 13870 54628
rect 16146 54572 16156 54628
rect 16212 54572 17612 54628
rect 17668 54572 17678 54628
rect 19506 54572 19516 54628
rect 19572 54572 20972 54628
rect 21028 54572 21038 54628
rect 27794 54572 27804 54628
rect 27860 54572 28476 54628
rect 28532 54572 28542 54628
rect 30594 54572 30604 54628
rect 30660 54572 30670 54628
rect 32162 54572 32172 54628
rect 32228 54572 35868 54628
rect 35924 54572 35934 54628
rect 36866 54572 36876 54628
rect 36932 54572 37212 54628
rect 37268 54572 37278 54628
rect 38434 54572 38444 54628
rect 38500 54572 40124 54628
rect 40180 54572 40190 54628
rect 44482 54572 44492 54628
rect 44548 54572 45612 54628
rect 45668 54572 45678 54628
rect 45836 54572 49980 54628
rect 50036 54572 50046 54628
rect 0 54516 800 54544
rect 12796 54516 12852 54572
rect 50372 54516 50428 54684
rect 52098 54572 52108 54628
rect 52164 54572 52780 54628
rect 52836 54572 53676 54628
rect 53732 54572 53742 54628
rect 0 54460 1708 54516
rect 1764 54460 1774 54516
rect 12786 54460 12796 54516
rect 12852 54460 13132 54516
rect 13188 54460 13198 54516
rect 13906 54460 13916 54516
rect 13972 54460 14252 54516
rect 14308 54460 14318 54516
rect 15820 54460 17948 54516
rect 18004 54460 18014 54516
rect 18610 54460 18620 54516
rect 18676 54460 20132 54516
rect 20738 54460 20748 54516
rect 20804 54460 21532 54516
rect 21588 54460 22540 54516
rect 22596 54460 22606 54516
rect 26226 54460 26236 54516
rect 26292 54460 29148 54516
rect 29204 54460 29214 54516
rect 29922 54460 29932 54516
rect 29988 54460 31276 54516
rect 31332 54460 31612 54516
rect 31668 54460 31678 54516
rect 45378 54460 45388 54516
rect 45444 54460 45724 54516
rect 45780 54460 46620 54516
rect 46676 54460 46686 54516
rect 50372 54460 51660 54516
rect 51716 54460 51726 54516
rect 53778 54460 53788 54516
rect 53844 54460 54684 54516
rect 54740 54460 54750 54516
rect 0 54432 800 54460
rect 15820 54404 15876 54460
rect 9650 54348 9660 54404
rect 9716 54348 10892 54404
rect 10948 54348 10958 54404
rect 12114 54348 12124 54404
rect 12180 54348 14812 54404
rect 14868 54348 15820 54404
rect 15876 54348 15886 54404
rect 16258 54348 16268 54404
rect 16324 54348 17836 54404
rect 17892 54348 19852 54404
rect 19908 54348 19918 54404
rect 20076 54292 20132 54460
rect 25106 54348 25116 54404
rect 25172 54348 31444 54404
rect 31826 54348 31836 54404
rect 31892 54348 33852 54404
rect 33908 54348 33918 54404
rect 34626 54348 34636 54404
rect 34692 54348 34702 54404
rect 42130 54348 42140 54404
rect 42196 54348 44940 54404
rect 44996 54348 45006 54404
rect 45602 54348 45612 54404
rect 45668 54348 46284 54404
rect 46340 54348 46350 54404
rect 52098 54348 52108 54404
rect 52164 54348 52444 54404
rect 52500 54348 52510 54404
rect 53218 54348 53228 54404
rect 53284 54348 56588 54404
rect 56644 54348 56654 54404
rect 31388 54292 31444 54348
rect 34636 54292 34692 54348
rect 10994 54236 11004 54292
rect 11060 54236 11340 54292
rect 11396 54236 11788 54292
rect 11844 54236 11854 54292
rect 12226 54236 12236 54292
rect 12292 54236 16156 54292
rect 16212 54236 16222 54292
rect 17612 54236 19516 54292
rect 19572 54236 19582 54292
rect 20076 54236 27244 54292
rect 27300 54236 27310 54292
rect 30370 54236 30380 54292
rect 30436 54236 30940 54292
rect 30996 54236 31006 54292
rect 31388 54236 34692 54292
rect 48850 54236 48860 54292
rect 48916 54236 49084 54292
rect 49140 54236 52892 54292
rect 52948 54236 52958 54292
rect 54338 54236 54348 54292
rect 54404 54236 54414 54292
rect 17612 54180 17668 54236
rect 49308 54180 49364 54236
rect 54348 54180 54404 54236
rect 10882 54124 10892 54180
rect 10948 54124 13692 54180
rect 13748 54124 17668 54180
rect 17826 54124 17836 54180
rect 17892 54124 18508 54180
rect 18564 54124 18574 54180
rect 19842 54124 19852 54180
rect 19908 54124 20636 54180
rect 20692 54124 20702 54180
rect 27682 54124 27692 54180
rect 27748 54124 30828 54180
rect 30884 54124 30894 54180
rect 31938 54124 31948 54180
rect 32004 54124 34076 54180
rect 34132 54124 34142 54180
rect 38882 54124 38892 54180
rect 38948 54124 46620 54180
rect 46676 54124 46686 54180
rect 49298 54124 49308 54180
rect 49364 54124 49374 54180
rect 52434 54124 52444 54180
rect 52500 54124 54404 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 13542 54012 13580 54068
rect 13636 54012 13646 54068
rect 13794 54012 13804 54068
rect 13860 54012 17500 54068
rect 17556 54012 17566 54068
rect 18050 54012 18060 54068
rect 18116 54012 23548 54068
rect 23604 54012 23614 54068
rect 43362 54012 43372 54068
rect 43428 54012 47852 54068
rect 47908 54012 47918 54068
rect 1586 53900 1596 53956
rect 1652 53900 12460 53956
rect 12516 53900 12526 53956
rect 13682 53900 13692 53956
rect 13748 53900 16380 53956
rect 16436 53900 16446 53956
rect 22754 53900 22764 53956
rect 22820 53900 23996 53956
rect 24052 53900 25452 53956
rect 25508 53900 25518 53956
rect 26562 53900 26572 53956
rect 26628 53900 27692 53956
rect 27748 53900 27758 53956
rect 30818 53900 30828 53956
rect 30884 53900 31276 53956
rect 31332 53900 31342 53956
rect 40450 53900 40460 53956
rect 40516 53900 57708 53956
rect 57764 53900 57774 53956
rect 11442 53788 11452 53844
rect 11508 53788 13524 53844
rect 13468 53732 13524 53788
rect 13916 53788 15932 53844
rect 15988 53788 15998 53844
rect 17602 53788 17612 53844
rect 17668 53788 21308 53844
rect 21364 53788 21374 53844
rect 22530 53788 22540 53844
rect 22596 53788 22606 53844
rect 25890 53788 25900 53844
rect 25956 53788 27356 53844
rect 27412 53788 27422 53844
rect 33170 53788 33180 53844
rect 33236 53788 35084 53844
rect 35140 53788 41356 53844
rect 41412 53788 41422 53844
rect 43922 53788 43932 53844
rect 43988 53788 45388 53844
rect 45444 53788 45454 53844
rect 46284 53788 46956 53844
rect 47012 53788 48188 53844
rect 48244 53788 48254 53844
rect 51874 53788 51884 53844
rect 51940 53788 51950 53844
rect 56914 53788 56924 53844
rect 56980 53788 58940 53844
rect 58996 53788 59006 53844
rect 13916 53732 13972 53788
rect 22540 53732 22596 53788
rect 46284 53732 46340 53788
rect 51884 53732 51940 53788
rect 11554 53676 11564 53732
rect 11620 53676 12908 53732
rect 12964 53676 12974 53732
rect 13468 53676 13972 53732
rect 15586 53676 15596 53732
rect 15652 53676 16044 53732
rect 16100 53676 16110 53732
rect 16258 53676 16268 53732
rect 16324 53676 17276 53732
rect 17332 53676 17342 53732
rect 18834 53676 18844 53732
rect 18900 53676 21532 53732
rect 21588 53676 21598 53732
rect 22540 53676 26684 53732
rect 26740 53676 26750 53732
rect 26852 53676 28588 53732
rect 28644 53676 28654 53732
rect 30594 53676 30604 53732
rect 30660 53676 31724 53732
rect 31780 53676 32620 53732
rect 32676 53676 32686 53732
rect 32834 53676 32844 53732
rect 32900 53676 36988 53732
rect 37044 53676 37054 53732
rect 26852 53620 26908 53676
rect 38612 53620 38668 53732
rect 38724 53676 38734 53732
rect 40002 53676 40012 53732
rect 40068 53676 42252 53732
rect 42308 53676 42318 53732
rect 42690 53676 42700 53732
rect 42756 53676 43708 53732
rect 43764 53676 43774 53732
rect 44258 53676 44268 53732
rect 44324 53676 45836 53732
rect 45892 53676 46340 53732
rect 46498 53676 46508 53732
rect 46564 53676 47516 53732
rect 47572 53676 47582 53732
rect 47730 53676 47740 53732
rect 47796 53676 49756 53732
rect 49812 53676 49822 53732
rect 51884 53676 52892 53732
rect 52948 53676 52958 53732
rect 53778 53676 53788 53732
rect 53844 53676 55132 53732
rect 55188 53676 56700 53732
rect 56756 53676 56766 53732
rect 58034 53676 58044 53732
rect 58100 53676 58492 53732
rect 58548 53676 59052 53732
rect 59108 53676 59118 53732
rect 9650 53564 9660 53620
rect 9716 53564 11900 53620
rect 11956 53564 11966 53620
rect 12338 53564 12348 53620
rect 12404 53564 14364 53620
rect 14420 53564 14430 53620
rect 15474 53564 15484 53620
rect 15540 53564 16828 53620
rect 16884 53564 16894 53620
rect 17154 53564 17164 53620
rect 17220 53564 19404 53620
rect 19460 53564 19470 53620
rect 20066 53564 20076 53620
rect 20132 53564 22204 53620
rect 22260 53564 22270 53620
rect 22642 53564 22652 53620
rect 22708 53564 22876 53620
rect 22932 53564 25228 53620
rect 25284 53564 26908 53620
rect 28130 53564 28140 53620
rect 28196 53564 32396 53620
rect 32452 53564 32462 53620
rect 34290 53564 34300 53620
rect 34356 53564 37660 53620
rect 37716 53564 38668 53620
rect 1474 53452 1484 53508
rect 1540 53452 8652 53508
rect 8708 53452 8718 53508
rect 9090 53452 9100 53508
rect 9156 53452 10220 53508
rect 10276 53452 10286 53508
rect 10546 53452 10556 53508
rect 10612 53452 11228 53508
rect 11284 53452 11294 53508
rect 11900 53396 11956 53564
rect 13570 53452 13580 53508
rect 13636 53452 16940 53508
rect 16996 53452 17006 53508
rect 17164 53396 17220 53564
rect 40012 53508 40068 53676
rect 18050 53452 18060 53508
rect 18116 53452 19180 53508
rect 19236 53452 19246 53508
rect 19404 53452 20300 53508
rect 20356 53452 22316 53508
rect 22372 53452 22382 53508
rect 26450 53452 26460 53508
rect 26516 53452 28252 53508
rect 28308 53452 28318 53508
rect 29698 53452 29708 53508
rect 29764 53452 30380 53508
rect 30436 53452 30446 53508
rect 31714 53452 31724 53508
rect 31780 53452 32508 53508
rect 32564 53452 32574 53508
rect 34514 53452 34524 53508
rect 34580 53452 35420 53508
rect 35476 53452 36204 53508
rect 36260 53452 36270 53508
rect 37202 53452 37212 53508
rect 37268 53452 40068 53508
rect 43708 53508 43764 53676
rect 45014 53564 45052 53620
rect 45108 53564 45118 53620
rect 45714 53564 45724 53620
rect 45780 53564 46844 53620
rect 46900 53564 51212 53620
rect 51268 53564 51278 53620
rect 51650 53564 51660 53620
rect 51716 53564 52556 53620
rect 52612 53564 52622 53620
rect 43708 53452 46060 53508
rect 46116 53452 46126 53508
rect 47506 53452 47516 53508
rect 47572 53452 49084 53508
rect 49140 53452 49150 53508
rect 49522 53452 49532 53508
rect 49588 53452 51436 53508
rect 51492 53452 51502 53508
rect 57922 53452 57932 53508
rect 57988 53452 59612 53508
rect 59668 53452 59678 53508
rect 60722 53452 60732 53508
rect 60788 53452 61068 53508
rect 61124 53452 62188 53508
rect 62244 53452 62254 53508
rect 19404 53396 19460 53452
rect 11900 53340 13804 53396
rect 13860 53340 13870 53396
rect 15138 53340 15148 53396
rect 15204 53340 17220 53396
rect 18498 53340 18508 53396
rect 18564 53340 19460 53396
rect 25330 53340 25340 53396
rect 25396 53340 38444 53396
rect 38500 53340 38668 53396
rect 42354 53340 42364 53396
rect 42420 53340 42812 53396
rect 42868 53340 44716 53396
rect 44772 53340 44782 53396
rect 46498 53340 46508 53396
rect 46564 53340 49980 53396
rect 50036 53340 50046 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 38612 53284 38668 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 8530 53228 8540 53284
rect 8596 53228 9884 53284
rect 9940 53228 13580 53284
rect 13636 53228 14700 53284
rect 14756 53228 14766 53284
rect 17042 53228 17052 53284
rect 17108 53228 18060 53284
rect 18116 53228 18126 53284
rect 21746 53228 21756 53284
rect 21812 53228 21822 53284
rect 26852 53228 30492 53284
rect 30548 53228 30558 53284
rect 30930 53228 30940 53284
rect 30996 53228 34524 53284
rect 34580 53228 34590 53284
rect 38612 53228 41132 53284
rect 41188 53228 41198 53284
rect 41906 53228 41916 53284
rect 41972 53228 47740 53284
rect 47796 53228 47806 53284
rect 48962 53228 48972 53284
rect 49028 53228 49196 53284
rect 49252 53228 49262 53284
rect 21756 53172 21812 53228
rect 26852 53172 26908 53228
rect 9090 53116 9100 53172
rect 9156 53116 14028 53172
rect 14084 53116 14094 53172
rect 14438 53116 14476 53172
rect 14532 53116 14542 53172
rect 15362 53116 15372 53172
rect 15428 53116 15438 53172
rect 19282 53116 19292 53172
rect 19348 53116 23212 53172
rect 23268 53116 23278 53172
rect 25778 53116 25788 53172
rect 25844 53116 26908 53172
rect 27010 53116 27020 53172
rect 27076 53116 28700 53172
rect 28756 53116 28766 53172
rect 29250 53116 29260 53172
rect 29316 53116 29708 53172
rect 29764 53116 29774 53172
rect 46386 53116 46396 53172
rect 46452 53116 47628 53172
rect 47684 53116 47694 53172
rect 48290 53116 48300 53172
rect 48356 53116 49420 53172
rect 49476 53116 52668 53172
rect 52724 53116 52734 53172
rect 53890 53116 53900 53172
rect 53956 53116 55132 53172
rect 55188 53116 55580 53172
rect 55636 53116 55646 53172
rect 56242 53116 56252 53172
rect 56308 53116 60732 53172
rect 60788 53116 60798 53172
rect 13234 53004 13244 53060
rect 13300 53004 15036 53060
rect 15092 53004 15102 53060
rect 6850 52892 6860 52948
rect 6916 52892 7756 52948
rect 7812 52892 14140 52948
rect 14196 52892 14206 52948
rect 14802 52892 14812 52948
rect 14868 52892 15148 52948
rect 15204 52892 15214 52948
rect 13682 52780 13692 52836
rect 13748 52780 15148 52836
rect 8306 52668 8316 52724
rect 8372 52668 11676 52724
rect 11732 52668 14812 52724
rect 14868 52668 14878 52724
rect 15092 52668 15148 52780
rect 15372 52724 15428 53116
rect 15922 53004 15932 53060
rect 15988 53004 16604 53060
rect 16660 53004 16670 53060
rect 17826 53004 17836 53060
rect 17892 53004 19964 53060
rect 20020 53004 20030 53060
rect 17490 52892 17500 52948
rect 17556 52892 21308 52948
rect 21364 52892 21374 52948
rect 21532 52836 21588 53116
rect 21746 53004 21756 53060
rect 21812 53004 22204 53060
rect 22260 53004 22270 53060
rect 27020 52948 27076 53116
rect 28578 53004 28588 53060
rect 28644 53004 34188 53060
rect 34244 53004 34254 53060
rect 38658 53004 38668 53060
rect 38724 53004 39340 53060
rect 39396 53004 40908 53060
rect 40964 53004 40974 53060
rect 45826 53004 45836 53060
rect 45892 53004 46732 53060
rect 46788 53004 48076 53060
rect 48132 53004 48142 53060
rect 55010 53004 55020 53060
rect 55076 53004 55356 53060
rect 55412 53004 57484 53060
rect 57540 53004 57550 53060
rect 24210 52892 24220 52948
rect 24276 52892 27076 52948
rect 29698 52892 29708 52948
rect 29764 52892 30492 52948
rect 30548 52892 30558 52948
rect 34178 52892 34188 52948
rect 34244 52892 35084 52948
rect 35140 52892 35150 52948
rect 44034 52892 44044 52948
rect 44100 52892 46508 52948
rect 46564 52892 46574 52948
rect 47730 52892 47740 52948
rect 47796 52892 49308 52948
rect 49364 52892 49374 52948
rect 49970 52892 49980 52948
rect 50036 52892 50988 52948
rect 51044 52892 53452 52948
rect 53508 52892 53518 52948
rect 19730 52780 19740 52836
rect 19796 52780 20524 52836
rect 20580 52780 20590 52836
rect 21532 52780 21756 52836
rect 21812 52780 21822 52836
rect 23538 52780 23548 52836
rect 23604 52780 25340 52836
rect 25396 52780 25406 52836
rect 29362 52780 29372 52836
rect 29428 52780 30156 52836
rect 30212 52780 31276 52836
rect 31332 52780 31342 52836
rect 31938 52780 31948 52836
rect 32004 52780 32396 52836
rect 32452 52780 32462 52836
rect 33282 52780 33292 52836
rect 33348 52780 36484 52836
rect 37426 52780 37436 52836
rect 37492 52780 38556 52836
rect 38612 52780 38622 52836
rect 44594 52780 44604 52836
rect 44660 52780 45388 52836
rect 45444 52780 45454 52836
rect 47954 52780 47964 52836
rect 48020 52780 49868 52836
rect 49924 52780 49934 52836
rect 54338 52780 54348 52836
rect 54404 52780 56588 52836
rect 56644 52780 56654 52836
rect 15204 52668 15214 52724
rect 15362 52668 15372 52724
rect 15428 52668 15438 52724
rect 16006 52668 16044 52724
rect 16100 52668 16110 52724
rect 19058 52668 19068 52724
rect 19124 52668 21420 52724
rect 21476 52668 21868 52724
rect 21924 52668 21934 52724
rect 26852 52668 28028 52724
rect 28084 52668 28094 52724
rect 31602 52668 31612 52724
rect 31668 52668 34636 52724
rect 34692 52668 34702 52724
rect 13794 52556 13804 52612
rect 13860 52556 15820 52612
rect 15876 52556 15886 52612
rect 16594 52556 16604 52612
rect 16660 52556 20636 52612
rect 20692 52556 20702 52612
rect 21522 52556 21532 52612
rect 21588 52556 23548 52612
rect 23604 52556 24220 52612
rect 24276 52556 24286 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 20636 52500 20692 52556
rect 14466 52444 14476 52500
rect 14532 52444 20580 52500
rect 20636 52444 26012 52500
rect 26068 52444 26572 52500
rect 26628 52444 26638 52500
rect 13458 52332 13468 52388
rect 13524 52332 14476 52388
rect 14532 52332 15148 52388
rect 17602 52332 17612 52388
rect 17668 52332 18172 52388
rect 18228 52332 18238 52388
rect 15092 52276 15148 52332
rect 20524 52276 20580 52444
rect 26852 52276 26908 52668
rect 27010 52556 27020 52612
rect 27076 52556 32844 52612
rect 32900 52556 32910 52612
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 36428 52500 36484 52780
rect 38098 52668 38108 52724
rect 38164 52668 38780 52724
rect 38836 52668 38846 52724
rect 48178 52668 48188 52724
rect 48244 52668 50204 52724
rect 50260 52668 50270 52724
rect 51538 52668 51548 52724
rect 51604 52668 53228 52724
rect 53284 52668 53294 52724
rect 55570 52668 55580 52724
rect 55636 52668 57148 52724
rect 57204 52668 57214 52724
rect 38546 52556 38556 52612
rect 38612 52556 44604 52612
rect 44660 52556 45052 52612
rect 45108 52556 45118 52612
rect 49186 52556 49196 52612
rect 49252 52556 50092 52612
rect 50148 52556 50158 52612
rect 54338 52556 54348 52612
rect 54404 52556 55468 52612
rect 55524 52556 55534 52612
rect 36418 52444 36428 52500
rect 36484 52444 38444 52500
rect 38500 52444 38510 52500
rect 43698 52444 43708 52500
rect 43764 52444 43820 52500
rect 43876 52444 43886 52500
rect 47282 52444 47292 52500
rect 47348 52444 52892 52500
rect 52948 52444 52958 52500
rect 53218 52444 53228 52500
rect 53284 52444 54460 52500
rect 54516 52444 54796 52500
rect 54852 52444 54862 52500
rect 30594 52332 30604 52388
rect 30660 52332 31612 52388
rect 31668 52332 31678 52388
rect 33506 52332 33516 52388
rect 33572 52332 37100 52388
rect 37156 52332 37166 52388
rect 42018 52332 42028 52388
rect 42084 52332 42700 52388
rect 42756 52332 43036 52388
rect 43092 52332 45948 52388
rect 46004 52332 46014 52388
rect 51314 52332 51324 52388
rect 51380 52332 53900 52388
rect 53956 52332 53966 52388
rect 8418 52220 8428 52276
rect 8484 52220 9100 52276
rect 9156 52220 9166 52276
rect 10210 52220 10220 52276
rect 10276 52220 14252 52276
rect 14308 52220 14318 52276
rect 15092 52220 15260 52276
rect 15316 52220 15326 52276
rect 20514 52220 20524 52276
rect 20580 52220 27580 52276
rect 27636 52220 27646 52276
rect 30370 52220 30380 52276
rect 30436 52220 31948 52276
rect 32004 52220 32844 52276
rect 32900 52220 32910 52276
rect 32844 52164 32900 52220
rect 34076 52164 34132 52332
rect 34290 52220 34300 52276
rect 34356 52220 34804 52276
rect 35410 52220 35420 52276
rect 35476 52220 36316 52276
rect 36372 52220 38388 52276
rect 43138 52220 43148 52276
rect 43204 52220 48300 52276
rect 48356 52220 48366 52276
rect 52210 52220 52220 52276
rect 52276 52220 54292 52276
rect 60722 52220 60732 52276
rect 60788 52220 61516 52276
rect 61572 52220 62636 52276
rect 62692 52220 62702 52276
rect 34748 52164 34804 52220
rect 38332 52164 38388 52220
rect 6178 52108 6188 52164
rect 6244 52108 7420 52164
rect 7476 52108 13692 52164
rect 13748 52108 13758 52164
rect 14690 52108 14700 52164
rect 14756 52108 15036 52164
rect 15092 52108 15102 52164
rect 16258 52108 16268 52164
rect 16324 52108 17388 52164
rect 17444 52108 17454 52164
rect 24322 52108 24332 52164
rect 24388 52108 25452 52164
rect 25508 52108 25518 52164
rect 27122 52108 27132 52164
rect 27188 52108 27804 52164
rect 27860 52108 27870 52164
rect 29250 52108 29260 52164
rect 29316 52108 30156 52164
rect 30212 52108 32172 52164
rect 32228 52108 32238 52164
rect 32844 52108 33516 52164
rect 33572 52108 33582 52164
rect 34076 52108 34580 52164
rect 34748 52108 34860 52164
rect 34916 52108 35532 52164
rect 35588 52108 35598 52164
rect 35858 52108 35868 52164
rect 35924 52108 35934 52164
rect 36194 52108 36204 52164
rect 36260 52108 36988 52164
rect 37044 52108 37054 52164
rect 38332 52108 38892 52164
rect 38948 52108 39228 52164
rect 39284 52108 39294 52164
rect 45154 52108 45164 52164
rect 45220 52108 45836 52164
rect 45892 52108 48076 52164
rect 48132 52108 48142 52164
rect 49970 52108 49980 52164
rect 50036 52108 50316 52164
rect 50372 52108 50382 52164
rect 51314 52108 51324 52164
rect 51380 52108 52780 52164
rect 52836 52108 52846 52164
rect 13906 51996 13916 52052
rect 13972 51996 16156 52052
rect 16212 51996 16222 52052
rect 17602 51996 17612 52052
rect 17668 51996 20412 52052
rect 20468 51996 20478 52052
rect 28914 51996 28924 52052
rect 28980 51996 29148 52052
rect 29204 51996 29214 52052
rect 30258 51996 30268 52052
rect 30324 51996 31836 52052
rect 31892 51996 33628 52052
rect 33684 51996 33694 52052
rect 34524 51940 34580 52108
rect 35868 52052 35924 52108
rect 38332 52052 38388 52108
rect 54236 52052 54292 52220
rect 58818 52108 58828 52164
rect 58884 52108 59052 52164
rect 59108 52108 59118 52164
rect 59602 52108 59612 52164
rect 59668 52108 62972 52164
rect 63028 52108 63038 52164
rect 34738 51996 34748 52052
rect 34804 51996 35924 52052
rect 38322 51996 38332 52052
rect 38388 51996 38398 52052
rect 41010 51996 41020 52052
rect 41076 51996 43036 52052
rect 43092 51996 43102 52052
rect 44594 51996 44604 52052
rect 44660 51996 46732 52052
rect 46788 51996 50316 52052
rect 50372 51996 50382 52052
rect 54226 51996 54236 52052
rect 54292 51996 54302 52052
rect 7186 51884 7196 51940
rect 7252 51884 8764 51940
rect 8820 51884 8830 51940
rect 10210 51884 10220 51940
rect 10276 51884 11676 51940
rect 11732 51884 13580 51940
rect 13636 51884 13646 51940
rect 14438 51884 14476 51940
rect 14532 51884 14542 51940
rect 17378 51884 17388 51940
rect 17444 51884 23996 51940
rect 24052 51884 24062 51940
rect 34524 51884 34972 51940
rect 35028 51884 35038 51940
rect 35410 51884 35420 51940
rect 35476 51884 36540 51940
rect 36596 51884 36606 51940
rect 52434 51884 52444 51940
rect 52500 51884 53676 51940
rect 53732 51884 53742 51940
rect 10098 51772 10108 51828
rect 10164 51772 12572 51828
rect 12628 51772 12638 51828
rect 12796 51772 13356 51828
rect 13412 51772 18844 51828
rect 18900 51772 18910 51828
rect 21410 51772 21420 51828
rect 21476 51772 26796 51828
rect 26852 51772 26862 51828
rect 34850 51772 34860 51828
rect 34916 51772 36428 51828
rect 36484 51772 36494 51828
rect 12796 51716 12852 51772
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 6514 51660 6524 51716
rect 6580 51660 12852 51716
rect 13458 51660 13468 51716
rect 13524 51660 17164 51716
rect 17220 51660 18396 51716
rect 18452 51660 18462 51716
rect 25414 51660 25452 51716
rect 25508 51660 25518 51716
rect 4834 51548 4844 51604
rect 4900 51548 5852 51604
rect 5908 51548 6860 51604
rect 6916 51548 6926 51604
rect 8642 51548 8652 51604
rect 8708 51548 11788 51604
rect 11844 51548 11854 51604
rect 14242 51548 14252 51604
rect 14308 51548 15148 51604
rect 15204 51548 15372 51604
rect 15428 51548 15438 51604
rect 16828 51548 17276 51604
rect 17332 51548 20076 51604
rect 20132 51548 20142 51604
rect 24434 51548 24444 51604
rect 24500 51548 25228 51604
rect 25284 51548 25294 51604
rect 25554 51548 25564 51604
rect 25620 51548 26348 51604
rect 26404 51548 26414 51604
rect 30482 51548 30492 51604
rect 30548 51548 32396 51604
rect 32452 51548 32462 51604
rect 34626 51548 34636 51604
rect 34692 51548 37212 51604
rect 37268 51548 37278 51604
rect 39890 51548 39900 51604
rect 39956 51548 40572 51604
rect 40628 51548 40638 51604
rect 43138 51548 43148 51604
rect 43204 51548 43708 51604
rect 43764 51548 43774 51604
rect 49532 51548 52948 51604
rect 55906 51548 55916 51604
rect 55972 51548 59388 51604
rect 59444 51548 59454 51604
rect 16828 51492 16884 51548
rect 16818 51436 16828 51492
rect 16884 51436 16894 51492
rect 18834 51436 18844 51492
rect 18900 51436 21532 51492
rect 21588 51436 21598 51492
rect 33954 51436 33964 51492
rect 34020 51436 35756 51492
rect 35812 51436 35822 51492
rect 38612 51436 41692 51492
rect 41748 51436 41758 51492
rect 15474 51324 15484 51380
rect 15540 51324 21868 51380
rect 21924 51324 21934 51380
rect 23986 51324 23996 51380
rect 24052 51324 24780 51380
rect 24836 51324 24846 51380
rect 26786 51324 26796 51380
rect 26852 51324 32172 51380
rect 32228 51324 32238 51380
rect 32386 51324 32396 51380
rect 32452 51324 33404 51380
rect 33460 51324 33470 51380
rect 34962 51324 34972 51380
rect 35028 51324 35420 51380
rect 35476 51324 35486 51380
rect 6822 51212 6860 51268
rect 6916 51212 6926 51268
rect 11554 51212 11564 51268
rect 11620 51212 12684 51268
rect 12740 51212 12750 51268
rect 13244 51212 13356 51268
rect 13412 51212 13422 51268
rect 14690 51212 14700 51268
rect 14756 51212 15820 51268
rect 15876 51212 15886 51268
rect 19506 51212 19516 51268
rect 19572 51212 21196 51268
rect 21252 51212 21644 51268
rect 21700 51212 21710 51268
rect 35298 51212 35308 51268
rect 35364 51212 36316 51268
rect 36372 51212 36382 51268
rect 13244 51156 13300 51212
rect 38612 51156 38668 51436
rect 49532 51380 49588 51548
rect 52892 51492 52948 51548
rect 50306 51436 50316 51492
rect 50372 51436 52108 51492
rect 52164 51436 52174 51492
rect 52892 51436 57036 51492
rect 57092 51436 57102 51492
rect 57474 51436 57484 51492
rect 57540 51436 58380 51492
rect 58436 51436 60844 51492
rect 60900 51436 60910 51492
rect 49186 51324 49196 51380
rect 49252 51324 49532 51380
rect 49588 51324 49598 51380
rect 50306 51324 50316 51380
rect 50372 51268 50428 51380
rect 52994 51324 53004 51380
rect 53060 51324 54572 51380
rect 54628 51324 58828 51380
rect 58884 51324 58894 51380
rect 48962 51212 48972 51268
rect 49028 51212 49868 51268
rect 49924 51212 49934 51268
rect 50372 51212 51828 51268
rect 57810 51212 57820 51268
rect 57876 51212 59164 51268
rect 59220 51212 59230 51268
rect 60050 51212 60060 51268
rect 60116 51212 60396 51268
rect 60452 51212 60462 51268
rect 6402 51100 6412 51156
rect 6468 51100 8204 51156
rect 8260 51100 12796 51156
rect 12852 51100 13300 51156
rect 16370 51100 16380 51156
rect 16436 51100 22316 51156
rect 22372 51100 22382 51156
rect 34524 51100 38668 51156
rect 43782 51100 43820 51156
rect 43876 51100 43886 51156
rect 34524 51044 34580 51100
rect 51772 51044 51828 51212
rect 52098 51100 52108 51156
rect 52164 51100 57708 51156
rect 57764 51100 57774 51156
rect 57922 51100 57932 51156
rect 57988 51100 61404 51156
rect 61460 51100 61740 51156
rect 61796 51100 61806 51156
rect 57708 51044 57764 51100
rect 9090 50988 9100 51044
rect 9156 50988 25788 51044
rect 25844 50988 25854 51044
rect 26852 50988 34524 51044
rect 34580 50988 34590 51044
rect 47954 50988 47964 51044
rect 48020 50988 48748 51044
rect 48804 50988 48814 51044
rect 51762 50988 51772 51044
rect 51828 50988 51838 51044
rect 53554 50988 53564 51044
rect 53620 50988 54124 51044
rect 54180 50988 54190 51044
rect 57708 50988 58716 51044
rect 58772 50988 58782 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 26852 50932 26908 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 11218 50876 11228 50932
rect 11284 50876 12348 50932
rect 12404 50876 12414 50932
rect 13682 50876 13692 50932
rect 13748 50876 26908 50932
rect 30482 50876 30492 50932
rect 30548 50876 32508 50932
rect 32564 50876 32574 50932
rect 35532 50876 43932 50932
rect 43988 50876 44492 50932
rect 44548 50876 46396 50932
rect 46452 50876 46462 50932
rect 48626 50876 48636 50932
rect 48692 50876 53284 50932
rect 57026 50876 57036 50932
rect 57092 50876 60620 50932
rect 60676 50876 61516 50932
rect 61572 50876 61740 50932
rect 61796 50876 61806 50932
rect 35532 50820 35588 50876
rect 9538 50764 9548 50820
rect 9604 50764 10220 50820
rect 10276 50764 10286 50820
rect 11778 50764 11788 50820
rect 11844 50764 12460 50820
rect 12516 50764 12526 50820
rect 13346 50764 13356 50820
rect 13412 50764 16044 50820
rect 16100 50764 16110 50820
rect 32050 50764 32060 50820
rect 32116 50764 35588 50820
rect 36306 50764 36316 50820
rect 36372 50764 39116 50820
rect 39172 50764 39788 50820
rect 39844 50764 40124 50820
rect 40180 50764 40190 50820
rect 49410 50764 49420 50820
rect 49476 50764 50764 50820
rect 50820 50764 50830 50820
rect 51538 50764 51548 50820
rect 51604 50764 51660 50820
rect 51716 50764 51726 50820
rect 53228 50708 53284 50876
rect 57250 50764 57260 50820
rect 57316 50764 59948 50820
rect 60004 50764 60014 50820
rect 4162 50652 4172 50708
rect 4228 50652 7868 50708
rect 7924 50652 8092 50708
rect 8148 50652 8158 50708
rect 9314 50652 9324 50708
rect 9380 50652 9996 50708
rect 10052 50652 10062 50708
rect 12562 50652 12572 50708
rect 12628 50652 13804 50708
rect 13860 50652 13870 50708
rect 15250 50652 15260 50708
rect 15316 50652 16268 50708
rect 16324 50652 16334 50708
rect 30146 50652 30156 50708
rect 30212 50652 33516 50708
rect 33572 50652 37436 50708
rect 37492 50652 37502 50708
rect 39218 50652 39228 50708
rect 39284 50652 41692 50708
rect 41748 50652 41758 50708
rect 49746 50652 49756 50708
rect 49812 50652 49980 50708
rect 50036 50652 50046 50708
rect 50306 50652 50316 50708
rect 50372 50652 51212 50708
rect 51268 50652 51436 50708
rect 51492 50652 51502 50708
rect 53218 50652 53228 50708
rect 53284 50652 53294 50708
rect 57026 50652 57036 50708
rect 57092 50652 60620 50708
rect 60676 50652 60686 50708
rect 2818 50540 2828 50596
rect 2884 50540 5180 50596
rect 5236 50540 6860 50596
rect 6916 50540 6926 50596
rect 7074 50540 7084 50596
rect 7140 50540 9436 50596
rect 9492 50540 9502 50596
rect 10098 50540 10108 50596
rect 10164 50540 10668 50596
rect 10724 50540 11564 50596
rect 11620 50540 11630 50596
rect 12674 50540 12684 50596
rect 12740 50540 13020 50596
rect 13076 50540 14364 50596
rect 14420 50540 14430 50596
rect 20514 50540 20524 50596
rect 20580 50540 22764 50596
rect 22820 50540 22830 50596
rect 28018 50540 28028 50596
rect 28084 50540 29932 50596
rect 29988 50540 30940 50596
rect 30996 50540 31500 50596
rect 31556 50540 31566 50596
rect 32610 50540 32620 50596
rect 32676 50540 32686 50596
rect 34486 50540 34524 50596
rect 34580 50540 34590 50596
rect 35074 50540 35084 50596
rect 35140 50540 35868 50596
rect 35924 50540 35934 50596
rect 38994 50540 39004 50596
rect 39060 50540 41244 50596
rect 41300 50540 41310 50596
rect 42774 50540 42812 50596
rect 42868 50540 42878 50596
rect 50978 50540 50988 50596
rect 51044 50540 53564 50596
rect 53620 50540 53630 50596
rect 55682 50540 55692 50596
rect 55748 50540 58044 50596
rect 58100 50540 58110 50596
rect 32620 50484 32676 50540
rect 4274 50428 4284 50484
rect 4340 50428 4396 50484
rect 4452 50428 4462 50484
rect 8978 50428 8988 50484
rect 9044 50428 15708 50484
rect 15764 50428 15774 50484
rect 20626 50428 20636 50484
rect 20692 50428 21756 50484
rect 21812 50428 21822 50484
rect 29810 50428 29820 50484
rect 29876 50428 31724 50484
rect 31780 50428 36316 50484
rect 36372 50428 36382 50484
rect 39554 50428 39564 50484
rect 39620 50428 41020 50484
rect 41076 50428 41086 50484
rect 44370 50428 44380 50484
rect 44436 50428 45724 50484
rect 45780 50428 47404 50484
rect 47460 50428 47470 50484
rect 49970 50428 49980 50484
rect 50036 50428 51492 50484
rect 51846 50428 51884 50484
rect 51940 50428 51950 50484
rect 56914 50428 56924 50484
rect 56980 50428 58492 50484
rect 58548 50428 58558 50484
rect 51436 50372 51492 50428
rect 6738 50316 6748 50372
rect 6804 50316 8316 50372
rect 8372 50316 8382 50372
rect 10434 50316 10444 50372
rect 10500 50316 12012 50372
rect 12068 50316 12078 50372
rect 12338 50316 12348 50372
rect 12404 50316 16604 50372
rect 16660 50316 16670 50372
rect 20290 50316 20300 50372
rect 20356 50316 20366 50372
rect 20738 50316 20748 50372
rect 20804 50316 24164 50372
rect 40338 50316 40348 50372
rect 40404 50316 40796 50372
rect 40852 50316 40862 50372
rect 44258 50316 44268 50372
rect 44324 50316 45052 50372
rect 45108 50316 45118 50372
rect 47282 50316 47292 50372
rect 47348 50316 48524 50372
rect 48580 50316 48590 50372
rect 49186 50316 49196 50372
rect 49252 50316 50428 50372
rect 50484 50316 50494 50372
rect 51426 50316 51436 50372
rect 51492 50316 51502 50372
rect 61170 50316 61180 50372
rect 61236 50316 61516 50372
rect 61572 50316 61582 50372
rect 20300 50260 20356 50316
rect 24108 50260 24164 50316
rect 48524 50260 48580 50316
rect 20300 50204 21308 50260
rect 21364 50204 21374 50260
rect 24098 50204 24108 50260
rect 24164 50204 24174 50260
rect 48524 50204 49644 50260
rect 49700 50204 49710 50260
rect 49942 50204 49980 50260
rect 50036 50204 50046 50260
rect 51734 50204 51772 50260
rect 51828 50204 51838 50260
rect 56690 50204 56700 50260
rect 56756 50204 61852 50260
rect 61908 50204 61918 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 8642 50092 8652 50148
rect 8708 50092 15148 50148
rect 20290 50092 20300 50148
rect 20356 50092 21644 50148
rect 21700 50092 29932 50148
rect 29988 50092 29998 50148
rect 30818 50092 30828 50148
rect 30884 50092 31164 50148
rect 31220 50092 32732 50148
rect 32788 50092 36652 50148
rect 36708 50092 36718 50148
rect 50166 50092 50204 50148
rect 50260 50092 50270 50148
rect 50978 50092 50988 50148
rect 51044 50092 51660 50148
rect 51716 50092 53676 50148
rect 53732 50092 53742 50148
rect 55794 50092 55804 50148
rect 55860 50092 57484 50148
rect 57540 50092 57550 50148
rect 15092 50036 15148 50092
rect 5954 49980 5964 50036
rect 6020 49980 6636 50036
rect 6692 49980 7084 50036
rect 7140 49980 7150 50036
rect 7298 49980 7308 50036
rect 7364 49980 9100 50036
rect 9156 49980 9166 50036
rect 15092 49980 16716 50036
rect 16772 49980 16782 50036
rect 24546 49980 24556 50036
rect 24612 49980 25676 50036
rect 25732 49980 25742 50036
rect 43474 49980 43484 50036
rect 43540 49980 45500 50036
rect 45556 49980 45566 50036
rect 53218 49980 53228 50036
rect 53284 49980 54908 50036
rect 54964 49980 54974 50036
rect 55234 49980 55244 50036
rect 55300 49980 56588 50036
rect 56644 49980 56654 50036
rect 8530 49868 8540 49924
rect 8596 49868 9660 49924
rect 9716 49868 9726 49924
rect 13794 49868 13804 49924
rect 13860 49868 14140 49924
rect 14196 49868 14206 49924
rect 15474 49868 15484 49924
rect 15540 49868 16380 49924
rect 16436 49868 17612 49924
rect 17668 49868 17678 49924
rect 18946 49868 18956 49924
rect 19012 49868 30380 49924
rect 30436 49868 30446 49924
rect 31490 49868 31500 49924
rect 31556 49868 33180 49924
rect 33236 49868 33246 49924
rect 37538 49868 37548 49924
rect 37604 49868 40348 49924
rect 40404 49868 40414 49924
rect 40562 49868 40572 49924
rect 40628 49868 42140 49924
rect 42196 49868 42206 49924
rect 2706 49756 2716 49812
rect 2772 49756 3388 49812
rect 3444 49756 14196 49812
rect 15698 49756 15708 49812
rect 15764 49756 19516 49812
rect 19572 49756 20076 49812
rect 20132 49756 20142 49812
rect 27122 49756 27132 49812
rect 27188 49756 27804 49812
rect 27860 49756 37884 49812
rect 37940 49756 37950 49812
rect 40786 49756 40796 49812
rect 40852 49756 42812 49812
rect 42868 49756 42878 49812
rect 14140 49700 14196 49756
rect 3332 49644 7756 49700
rect 7812 49644 7822 49700
rect 8866 49644 8876 49700
rect 8932 49644 12124 49700
rect 12180 49644 12190 49700
rect 14130 49644 14140 49700
rect 14196 49644 14206 49700
rect 14466 49644 14476 49700
rect 14532 49644 14812 49700
rect 14868 49644 14878 49700
rect 16034 49644 16044 49700
rect 16100 49644 16380 49700
rect 16436 49644 16446 49700
rect 18050 49644 18060 49700
rect 18116 49644 21308 49700
rect 21364 49644 21374 49700
rect 27682 49644 27692 49700
rect 27748 49644 29820 49700
rect 29876 49644 29886 49700
rect 31938 49644 31948 49700
rect 32004 49644 41356 49700
rect 41412 49644 41422 49700
rect 3332 49588 3388 49644
rect 43484 49588 43540 49980
rect 54908 49924 54964 49980
rect 49746 49868 49756 49924
rect 49812 49868 50204 49924
rect 50260 49868 53116 49924
rect 53172 49868 53182 49924
rect 54908 49868 57148 49924
rect 57204 49868 57214 49924
rect 46946 49756 46956 49812
rect 47012 49756 47740 49812
rect 47796 49756 47806 49812
rect 53778 49756 53788 49812
rect 53844 49756 54236 49812
rect 54292 49756 56924 49812
rect 56980 49756 59052 49812
rect 59108 49756 59118 49812
rect 47058 49644 47068 49700
rect 47124 49644 47516 49700
rect 47572 49644 48972 49700
rect 49028 49644 52556 49700
rect 52612 49644 52622 49700
rect 55346 49644 55356 49700
rect 55412 49644 57932 49700
rect 57988 49644 57998 49700
rect 60274 49644 60284 49700
rect 60340 49644 61516 49700
rect 61572 49644 61582 49700
rect 1586 49532 1596 49588
rect 1652 49532 3388 49588
rect 3938 49532 3948 49588
rect 4004 49532 5516 49588
rect 5572 49532 5582 49588
rect 13906 49532 13916 49588
rect 13972 49532 15372 49588
rect 15428 49532 15438 49588
rect 18498 49532 18508 49588
rect 18564 49532 19964 49588
rect 20020 49532 20030 49588
rect 29026 49532 29036 49588
rect 29092 49532 29708 49588
rect 29764 49532 29774 49588
rect 31826 49532 31836 49588
rect 31892 49532 35756 49588
rect 35812 49532 35822 49588
rect 38612 49532 38780 49588
rect 38836 49532 38846 49588
rect 43362 49532 43372 49588
rect 43428 49532 43540 49588
rect 46050 49532 46060 49588
rect 46116 49532 51660 49588
rect 51716 49532 51726 49588
rect 53778 49532 53788 49588
rect 53844 49532 57820 49588
rect 57876 49532 57886 49588
rect 15250 49420 15260 49476
rect 15316 49420 15484 49476
rect 15540 49420 16044 49476
rect 16100 49420 19740 49476
rect 19796 49420 33740 49476
rect 33796 49420 33806 49476
rect 34150 49420 34188 49476
rect 34244 49420 34254 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 38612 49364 38668 49532
rect 46610 49420 46620 49476
rect 46676 49420 55804 49476
rect 55860 49420 55870 49476
rect 8306 49308 8316 49364
rect 8372 49308 16828 49364
rect 16884 49308 17388 49364
rect 17444 49308 17454 49364
rect 18274 49308 18284 49364
rect 18340 49308 21532 49364
rect 21588 49308 21598 49364
rect 35970 49308 35980 49364
rect 36036 49308 37436 49364
rect 37492 49308 38668 49364
rect 45826 49308 45836 49364
rect 45892 49308 47964 49364
rect 48020 49308 48860 49364
rect 48916 49308 48926 49364
rect 58034 49308 58044 49364
rect 58100 49308 59948 49364
rect 60004 49308 60014 49364
rect 1922 49196 1932 49252
rect 1988 49196 2492 49252
rect 2548 49196 8428 49252
rect 8484 49196 8494 49252
rect 10994 49196 11004 49252
rect 11060 49196 13916 49252
rect 13972 49196 13982 49252
rect 14130 49196 14140 49252
rect 14196 49196 27020 49252
rect 27076 49196 27086 49252
rect 29586 49196 29596 49252
rect 29652 49196 30940 49252
rect 30996 49196 31836 49252
rect 31892 49196 31902 49252
rect 34962 49196 34972 49252
rect 35028 49196 37660 49252
rect 37716 49196 37726 49252
rect 37874 49196 37884 49252
rect 37940 49196 40964 49252
rect 41122 49196 41132 49252
rect 41188 49196 42700 49252
rect 42756 49196 42766 49252
rect 47170 49196 47180 49252
rect 47236 49196 47740 49252
rect 47796 49196 47806 49252
rect 50418 49196 50428 49252
rect 50484 49196 52052 49252
rect 52882 49196 52892 49252
rect 52948 49196 54572 49252
rect 54628 49196 55692 49252
rect 55748 49196 55758 49252
rect 57474 49196 57484 49252
rect 57540 49196 58156 49252
rect 58212 49196 58716 49252
rect 58772 49196 58782 49252
rect 40908 49140 40964 49196
rect 51996 49140 52052 49196
rect 3826 49084 3836 49140
rect 3892 49084 4508 49140
rect 4564 49084 5628 49140
rect 5684 49084 5694 49140
rect 9874 49084 9884 49140
rect 9940 49084 10444 49140
rect 10500 49084 12236 49140
rect 12292 49084 12302 49140
rect 18386 49084 18396 49140
rect 18452 49084 21420 49140
rect 21476 49084 21486 49140
rect 25330 49084 25340 49140
rect 25396 49084 39508 49140
rect 40908 49084 44044 49140
rect 44100 49084 44110 49140
rect 45490 49084 45500 49140
rect 45556 49084 49028 49140
rect 49298 49084 49308 49140
rect 49364 49084 50876 49140
rect 50932 49084 50942 49140
rect 51986 49084 51996 49140
rect 52052 49084 52780 49140
rect 52836 49084 52846 49140
rect 57138 49084 57148 49140
rect 57204 49084 58380 49140
rect 58436 49084 59276 49140
rect 59332 49084 59342 49140
rect 4050 48972 4060 49028
rect 4116 48972 4732 49028
rect 4788 48972 5852 49028
rect 5908 48972 5918 49028
rect 16594 48972 16604 49028
rect 16660 48972 16670 49028
rect 17602 48972 17612 49028
rect 17668 48972 18284 49028
rect 18340 48972 18350 49028
rect 30034 48972 30044 49028
rect 30100 48972 30604 49028
rect 30660 48972 32172 49028
rect 32228 48972 32238 49028
rect 35644 48972 36876 49028
rect 36932 48972 36942 49028
rect 37202 48972 37212 49028
rect 37268 48972 38108 49028
rect 38164 48972 38556 49028
rect 38612 48972 38622 49028
rect 16604 48916 16660 48972
rect 35644 48916 35700 48972
rect 39452 48916 39508 49084
rect 42354 48972 42364 49028
rect 42420 48972 45948 49028
rect 46004 48972 46014 49028
rect 46274 48972 46284 49028
rect 46340 48972 47180 49028
rect 47236 48972 47246 49028
rect 48972 48916 49028 49084
rect 49858 48972 49868 49028
rect 49924 48972 50764 49028
rect 50820 48972 50830 49028
rect 55458 48972 55468 49028
rect 55524 48972 58156 49028
rect 58212 48972 59052 49028
rect 59108 48972 59612 49028
rect 59668 48972 59678 49028
rect 2034 48860 2044 48916
rect 2100 48860 2716 48916
rect 2772 48860 2782 48916
rect 3490 48860 3500 48916
rect 3556 48860 4956 48916
rect 5012 48860 5022 48916
rect 11302 48860 11340 48916
rect 11396 48860 11406 48916
rect 12898 48860 12908 48916
rect 12964 48860 14364 48916
rect 14420 48860 14430 48916
rect 16604 48860 21756 48916
rect 21812 48860 21822 48916
rect 26674 48860 26684 48916
rect 26740 48860 27244 48916
rect 27300 48860 27310 48916
rect 33618 48860 33628 48916
rect 33684 48860 35644 48916
rect 35700 48860 35710 48916
rect 36082 48860 36092 48916
rect 36148 48860 37380 48916
rect 39442 48860 39452 48916
rect 39508 48860 39518 48916
rect 43250 48860 43260 48916
rect 43316 48860 43326 48916
rect 43474 48860 43484 48916
rect 43540 48860 45052 48916
rect 45108 48860 47068 48916
rect 47124 48860 47134 48916
rect 47730 48860 47740 48916
rect 47796 48860 48748 48916
rect 48804 48860 48814 48916
rect 48972 48860 52556 48916
rect 52612 48860 56700 48916
rect 56756 48860 56766 48916
rect 58482 48860 58492 48916
rect 58548 48860 60508 48916
rect 60564 48860 60574 48916
rect 60722 48860 60732 48916
rect 60788 48860 61740 48916
rect 61796 48860 61806 48916
rect 37324 48804 37380 48860
rect 43260 48804 43316 48860
rect 1670 48748 1708 48804
rect 1764 48748 1774 48804
rect 3910 48748 3948 48804
rect 4004 48748 4014 48804
rect 12562 48748 12572 48804
rect 12628 48748 15260 48804
rect 15316 48748 16604 48804
rect 16660 48748 18508 48804
rect 18564 48748 18574 48804
rect 23874 48748 23884 48804
rect 23940 48748 24780 48804
rect 24836 48748 25452 48804
rect 25508 48748 25518 48804
rect 29586 48748 29596 48804
rect 29652 48748 31052 48804
rect 31108 48748 31118 48804
rect 35298 48748 35308 48804
rect 35364 48748 36652 48804
rect 36708 48748 36718 48804
rect 37314 48748 37324 48804
rect 37380 48748 41468 48804
rect 41524 48748 41534 48804
rect 43260 48748 43820 48804
rect 43876 48748 43886 48804
rect 46050 48748 46060 48804
rect 46116 48748 47628 48804
rect 47684 48748 48188 48804
rect 48244 48748 49196 48804
rect 49252 48748 49262 48804
rect 51090 48748 51100 48804
rect 51156 48748 51772 48804
rect 51828 48748 51838 48804
rect 56354 48748 56364 48804
rect 56420 48748 58716 48804
rect 58772 48748 58782 48804
rect 59154 48748 59164 48804
rect 59220 48748 59836 48804
rect 59892 48748 60732 48804
rect 60788 48748 61628 48804
rect 61684 48748 61694 48804
rect 4162 48636 4172 48692
rect 4228 48636 6076 48692
rect 6132 48636 6142 48692
rect 8754 48636 8764 48692
rect 8820 48636 15148 48692
rect 29922 48636 29932 48692
rect 29988 48636 33180 48692
rect 33236 48636 33246 48692
rect 33730 48636 33740 48692
rect 33796 48636 35084 48692
rect 35140 48636 35644 48692
rect 35700 48636 35710 48692
rect 39666 48636 39676 48692
rect 39732 48636 41132 48692
rect 41188 48636 41198 48692
rect 42802 48636 42812 48692
rect 42868 48636 43260 48692
rect 43316 48636 43326 48692
rect 50988 48636 57036 48692
rect 57092 48636 57102 48692
rect 15092 48580 15148 48636
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 33180 48580 33236 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 13570 48524 13580 48580
rect 13636 48524 14588 48580
rect 14644 48524 14654 48580
rect 15092 48524 16156 48580
rect 16212 48524 16222 48580
rect 33180 48524 37772 48580
rect 37828 48524 37838 48580
rect 38098 48524 38108 48580
rect 38164 48524 40236 48580
rect 40292 48524 40302 48580
rect 42354 48524 42364 48580
rect 42420 48524 43148 48580
rect 43204 48524 43214 48580
rect 49158 48524 49196 48580
rect 49252 48524 49262 48580
rect 37772 48468 37828 48524
rect 50988 48468 51044 48636
rect 22082 48412 22092 48468
rect 22148 48412 23324 48468
rect 23380 48412 23996 48468
rect 24052 48412 24062 48468
rect 29810 48412 29820 48468
rect 29876 48412 35308 48468
rect 35364 48412 35374 48468
rect 36540 48412 37436 48468
rect 37492 48412 37502 48468
rect 37772 48412 39228 48468
rect 39284 48412 39294 48468
rect 40114 48412 40124 48468
rect 40180 48412 42028 48468
rect 42084 48412 42094 48468
rect 45266 48412 45276 48468
rect 45332 48412 48748 48468
rect 48804 48412 51044 48468
rect 56690 48412 56700 48468
rect 56756 48412 57036 48468
rect 57092 48412 59724 48468
rect 59780 48412 59790 48468
rect 36540 48356 36596 48412
rect 7522 48300 7532 48356
rect 7588 48300 11396 48356
rect 11890 48300 11900 48356
rect 11956 48300 13132 48356
rect 13188 48300 14252 48356
rect 14308 48300 14318 48356
rect 16482 48300 16492 48356
rect 16548 48300 18508 48356
rect 18564 48300 18574 48356
rect 22306 48300 22316 48356
rect 22372 48300 23772 48356
rect 23828 48300 28028 48356
rect 28084 48300 28094 48356
rect 29586 48300 29596 48356
rect 29652 48300 30604 48356
rect 30660 48300 30670 48356
rect 33058 48300 33068 48356
rect 33124 48300 36596 48356
rect 36652 48300 38668 48356
rect 40002 48300 40012 48356
rect 40068 48300 41580 48356
rect 41636 48300 45164 48356
rect 45220 48300 45230 48356
rect 49858 48300 49868 48356
rect 49924 48300 50316 48356
rect 50372 48300 50382 48356
rect 50866 48300 50876 48356
rect 50932 48300 51884 48356
rect 51940 48300 51950 48356
rect 57026 48300 57036 48356
rect 57092 48300 57820 48356
rect 57876 48300 58940 48356
rect 58996 48300 59006 48356
rect 62038 48300 62076 48356
rect 62132 48300 62142 48356
rect 1250 48188 1260 48244
rect 1316 48188 1932 48244
rect 1988 48188 2380 48244
rect 2436 48188 2446 48244
rect 8306 48188 8316 48244
rect 8372 48188 10556 48244
rect 10612 48188 10622 48244
rect 11340 48132 11396 48300
rect 36652 48244 36708 48300
rect 38612 48244 38668 48300
rect 12786 48188 12796 48244
rect 12852 48188 14700 48244
rect 14756 48188 14766 48244
rect 15922 48188 15932 48244
rect 15988 48188 18060 48244
rect 18116 48188 18126 48244
rect 19170 48188 19180 48244
rect 19236 48188 20524 48244
rect 20580 48188 20590 48244
rect 28242 48188 28252 48244
rect 28308 48188 29036 48244
rect 29092 48188 34860 48244
rect 34916 48188 34926 48244
rect 36642 48188 36652 48244
rect 36708 48188 36718 48244
rect 37202 48188 37212 48244
rect 37268 48188 37278 48244
rect 38612 48188 39564 48244
rect 39620 48188 39630 48244
rect 40338 48188 40348 48244
rect 40404 48188 42588 48244
rect 42644 48188 43372 48244
rect 43428 48188 43438 48244
rect 44594 48188 44604 48244
rect 44660 48188 45388 48244
rect 45444 48188 45454 48244
rect 46610 48188 46620 48244
rect 46676 48188 51772 48244
rect 51828 48188 51838 48244
rect 57894 48188 57932 48244
rect 57988 48188 60956 48244
rect 61012 48188 61964 48244
rect 62020 48188 62030 48244
rect 37212 48132 37268 48188
rect 1670 48076 1708 48132
rect 1764 48076 7084 48132
rect 7140 48076 7150 48132
rect 11340 48076 15820 48132
rect 15876 48076 15886 48132
rect 30370 48076 30380 48132
rect 30436 48076 33852 48132
rect 33908 48076 33918 48132
rect 34402 48076 34412 48132
rect 34468 48076 35084 48132
rect 35140 48076 35150 48132
rect 37212 48076 40012 48132
rect 40068 48076 40078 48132
rect 42130 48076 42140 48132
rect 42196 48076 43036 48132
rect 43092 48076 43102 48132
rect 43586 48076 43596 48132
rect 43652 48076 45500 48132
rect 45556 48076 45566 48132
rect 46722 48076 46732 48132
rect 46788 48076 51324 48132
rect 51380 48076 51390 48132
rect 55010 48076 55020 48132
rect 55076 48076 58044 48132
rect 58100 48076 58492 48132
rect 58548 48076 58558 48132
rect 33852 48020 33908 48076
rect 12338 47964 12348 48020
rect 12404 47964 18284 48020
rect 18340 47964 18350 48020
rect 23650 47964 23660 48020
rect 23716 47964 25900 48020
rect 25956 47964 28476 48020
rect 28532 47964 28542 48020
rect 33852 47964 38108 48020
rect 38164 47964 38174 48020
rect 46274 47964 46284 48020
rect 46340 47964 47740 48020
rect 47796 47964 47806 48020
rect 49410 47964 49420 48020
rect 49476 47964 51660 48020
rect 51716 47964 51726 48020
rect 14130 47852 14140 47908
rect 14196 47852 15484 47908
rect 15540 47852 21084 47908
rect 21140 47852 26908 47908
rect 28354 47852 28364 47908
rect 28420 47852 29820 47908
rect 29876 47852 29886 47908
rect 37874 47852 37884 47908
rect 37940 47852 38444 47908
rect 38500 47852 38510 47908
rect 40226 47852 40236 47908
rect 40292 47852 50876 47908
rect 50932 47852 50942 47908
rect 56914 47852 56924 47908
rect 56980 47852 62076 47908
rect 62132 47852 62142 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 26852 47796 26908 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 4946 47740 4956 47796
rect 5012 47740 5022 47796
rect 9202 47740 9212 47796
rect 9268 47740 9884 47796
rect 9940 47740 9950 47796
rect 16258 47740 16268 47796
rect 16324 47740 16604 47796
rect 16660 47740 19292 47796
rect 19348 47740 19964 47796
rect 20020 47740 20524 47796
rect 20580 47740 20590 47796
rect 23538 47740 23548 47796
rect 23604 47740 23996 47796
rect 24052 47740 24062 47796
rect 26852 47740 33068 47796
rect 33124 47740 33134 47796
rect 43698 47740 43708 47796
rect 43764 47740 47516 47796
rect 47572 47740 47582 47796
rect 50642 47740 50652 47796
rect 50708 47740 51436 47796
rect 51492 47740 51502 47796
rect 53218 47740 53228 47796
rect 53284 47740 55468 47796
rect 55524 47740 55534 47796
rect 56018 47740 56028 47796
rect 56084 47740 58492 47796
rect 58548 47740 58558 47796
rect 60946 47740 60956 47796
rect 61012 47740 61348 47796
rect 4956 47684 5012 47740
rect 61292 47684 61348 47740
rect 4722 47628 4732 47684
rect 4788 47628 5012 47684
rect 8306 47628 8316 47684
rect 8372 47628 11228 47684
rect 11284 47628 11294 47684
rect 18610 47628 18620 47684
rect 18676 47628 19852 47684
rect 19908 47628 19918 47684
rect 22194 47628 22204 47684
rect 22260 47628 25004 47684
rect 25060 47628 26572 47684
rect 26628 47628 26638 47684
rect 26852 47628 32060 47684
rect 32116 47628 32126 47684
rect 34290 47628 34300 47684
rect 34356 47628 35308 47684
rect 35364 47628 35374 47684
rect 37202 47628 37212 47684
rect 37268 47628 40684 47684
rect 40740 47628 41580 47684
rect 41636 47628 41646 47684
rect 43810 47628 43820 47684
rect 43876 47628 45612 47684
rect 45668 47628 45678 47684
rect 48066 47628 48076 47684
rect 48132 47628 51212 47684
rect 51268 47628 51278 47684
rect 54786 47628 54796 47684
rect 54852 47628 55356 47684
rect 55412 47628 59276 47684
rect 59332 47628 59342 47684
rect 61282 47628 61292 47684
rect 61348 47628 61358 47684
rect 61506 47628 61516 47684
rect 61572 47628 61582 47684
rect 26852 47572 26908 47628
rect 61516 47572 61572 47628
rect 8418 47516 8428 47572
rect 8484 47516 10556 47572
rect 10612 47516 10622 47572
rect 10882 47516 10892 47572
rect 10948 47516 13020 47572
rect 13076 47516 13086 47572
rect 18050 47516 18060 47572
rect 18116 47516 21308 47572
rect 21364 47516 21374 47572
rect 22530 47516 22540 47572
rect 22596 47516 26908 47572
rect 28130 47516 28140 47572
rect 28196 47516 30604 47572
rect 30660 47516 30670 47572
rect 33058 47516 33068 47572
rect 33124 47516 39228 47572
rect 39284 47516 39294 47572
rect 42690 47516 42700 47572
rect 42756 47516 44828 47572
rect 44884 47516 44894 47572
rect 51314 47516 51324 47572
rect 51380 47516 52444 47572
rect 52500 47516 52510 47572
rect 54226 47516 54236 47572
rect 54292 47516 58380 47572
rect 58436 47516 58446 47572
rect 61058 47516 61068 47572
rect 61124 47516 61572 47572
rect 7410 47404 7420 47460
rect 7476 47404 11900 47460
rect 11956 47404 11966 47460
rect 12674 47404 12684 47460
rect 12740 47404 13468 47460
rect 13524 47404 13534 47460
rect 18162 47404 18172 47460
rect 18228 47404 20300 47460
rect 20356 47404 20366 47460
rect 24434 47404 24444 47460
rect 24500 47404 26012 47460
rect 26068 47404 26078 47460
rect 28690 47404 28700 47460
rect 28756 47404 30044 47460
rect 30100 47404 30110 47460
rect 31042 47404 31052 47460
rect 31108 47404 31500 47460
rect 31556 47404 32284 47460
rect 32340 47404 32350 47460
rect 34290 47404 34300 47460
rect 34356 47404 36652 47460
rect 36708 47404 36718 47460
rect 40002 47404 40012 47460
rect 40068 47404 41804 47460
rect 41860 47404 41870 47460
rect 43474 47404 43484 47460
rect 43540 47404 44156 47460
rect 44212 47404 44222 47460
rect 45714 47404 45724 47460
rect 45780 47404 46844 47460
rect 46900 47404 47516 47460
rect 47572 47404 48300 47460
rect 48356 47404 48366 47460
rect 54898 47404 54908 47460
rect 54964 47404 55468 47460
rect 55524 47404 58268 47460
rect 58324 47404 58334 47460
rect 60582 47404 60620 47460
rect 60676 47404 60686 47460
rect 4946 47292 4956 47348
rect 5012 47292 5404 47348
rect 5460 47292 6524 47348
rect 6580 47292 6590 47348
rect 8642 47292 8652 47348
rect 8708 47292 9212 47348
rect 9268 47292 9548 47348
rect 9604 47292 9614 47348
rect 13794 47292 13804 47348
rect 13860 47292 14364 47348
rect 14420 47292 15372 47348
rect 15428 47292 16268 47348
rect 16324 47292 16334 47348
rect 26898 47292 26908 47348
rect 26964 47292 29372 47348
rect 29428 47292 29708 47348
rect 29764 47292 29774 47348
rect 36978 47292 36988 47348
rect 37044 47292 37212 47348
rect 37268 47292 37278 47348
rect 39106 47292 39116 47348
rect 39172 47292 42588 47348
rect 42644 47292 42654 47348
rect 43362 47292 43372 47348
rect 43428 47292 45836 47348
rect 45892 47292 45902 47348
rect 50194 47292 50204 47348
rect 50260 47292 56700 47348
rect 56756 47292 56766 47348
rect 58034 47292 58044 47348
rect 58100 47292 60732 47348
rect 60788 47292 60798 47348
rect 5058 47180 5068 47236
rect 5124 47180 5628 47236
rect 5684 47180 8316 47236
rect 8372 47180 8382 47236
rect 9650 47180 9660 47236
rect 9716 47180 10332 47236
rect 10388 47180 10398 47236
rect 10658 47180 10668 47236
rect 10724 47180 13468 47236
rect 13524 47180 13534 47236
rect 15484 47180 25900 47236
rect 25956 47180 25966 47236
rect 29138 47180 29148 47236
rect 29204 47180 31948 47236
rect 32004 47180 32014 47236
rect 32162 47180 32172 47236
rect 32228 47180 44268 47236
rect 44324 47180 49420 47236
rect 49476 47180 49486 47236
rect 53890 47180 53900 47236
rect 53956 47180 60620 47236
rect 60676 47180 60686 47236
rect 15484 47124 15540 47180
rect 62132 47124 62188 47348
rect 62244 47292 62254 47348
rect 8978 47068 8988 47124
rect 9044 47068 9884 47124
rect 9940 47068 14700 47124
rect 14756 47068 14766 47124
rect 15474 47068 15484 47124
rect 15540 47068 15550 47124
rect 27468 47068 28028 47124
rect 28084 47068 28094 47124
rect 43138 47068 43148 47124
rect 43204 47068 45836 47124
rect 45892 47068 45902 47124
rect 48710 47068 48748 47124
rect 48804 47068 48814 47124
rect 55234 47068 55244 47124
rect 55300 47068 56252 47124
rect 56308 47068 56318 47124
rect 57698 47068 57708 47124
rect 57764 47068 59276 47124
rect 59332 47068 60284 47124
rect 60340 47068 62188 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 27468 47012 27524 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 1474 46956 1484 47012
rect 1540 46956 3948 47012
rect 4004 46956 4014 47012
rect 9650 46956 9660 47012
rect 9716 46956 10108 47012
rect 10164 46956 10174 47012
rect 11666 46956 11676 47012
rect 11732 46956 13132 47012
rect 13188 46956 13198 47012
rect 16146 46956 16156 47012
rect 16212 46956 17948 47012
rect 18004 46956 18014 47012
rect 24630 46956 24668 47012
rect 24724 46956 24734 47012
rect 27458 46956 27468 47012
rect 27524 46956 27534 47012
rect 30930 46956 30940 47012
rect 30996 46956 34076 47012
rect 34132 46956 34142 47012
rect 36306 46956 36316 47012
rect 36372 46956 41916 47012
rect 41972 46956 42812 47012
rect 42868 46956 42878 47012
rect 45938 46956 45948 47012
rect 46004 46956 47516 47012
rect 47572 46956 48636 47012
rect 48692 46956 48702 47012
rect 48962 46956 48972 47012
rect 49028 46956 50316 47012
rect 50372 46956 50382 47012
rect 60694 46956 60732 47012
rect 60788 46956 60798 47012
rect 61282 46956 61292 47012
rect 61348 46956 61516 47012
rect 61572 46956 61582 47012
rect 61954 46956 61964 47012
rect 62020 46956 62058 47012
rect 2482 46844 2492 46900
rect 2548 46844 3612 46900
rect 3668 46844 3678 46900
rect 5282 46844 5292 46900
rect 5348 46844 7308 46900
rect 7364 46844 9772 46900
rect 9828 46844 9838 46900
rect 10210 46844 10220 46900
rect 10276 46844 11116 46900
rect 11172 46844 11182 46900
rect 13010 46844 13020 46900
rect 13076 46844 14028 46900
rect 14084 46844 14094 46900
rect 14466 46844 14476 46900
rect 14532 46844 15372 46900
rect 15428 46844 15438 46900
rect 18498 46844 18508 46900
rect 18564 46844 19740 46900
rect 19796 46844 20188 46900
rect 20244 46844 20254 46900
rect 22950 46844 22988 46900
rect 23044 46844 23054 46900
rect 23314 46844 23324 46900
rect 23380 46844 26908 46900
rect 31266 46844 31276 46900
rect 31332 46844 36428 46900
rect 36484 46844 36494 46900
rect 38612 46844 40236 46900
rect 40292 46844 40302 46900
rect 43250 46844 43260 46900
rect 43316 46844 44044 46900
rect 44100 46844 44110 46900
rect 49410 46844 49420 46900
rect 49476 46844 50204 46900
rect 50260 46844 52892 46900
rect 52948 46844 52958 46900
rect 53666 46844 53676 46900
rect 53732 46844 57820 46900
rect 57876 46844 57886 46900
rect 61730 46844 61740 46900
rect 61796 46844 62188 46900
rect 62244 46844 62254 46900
rect 2258 46732 2268 46788
rect 2324 46732 6188 46788
rect 6244 46732 6860 46788
rect 6916 46732 6926 46788
rect 8866 46732 8876 46788
rect 8932 46732 10444 46788
rect 10500 46732 10510 46788
rect 10854 46732 10892 46788
rect 10948 46732 10958 46788
rect 15922 46732 15932 46788
rect 15988 46732 17276 46788
rect 17332 46732 17342 46788
rect 17714 46732 17724 46788
rect 17780 46732 22876 46788
rect 22932 46732 22942 46788
rect 24546 46732 24556 46788
rect 24612 46732 25564 46788
rect 25620 46732 25630 46788
rect 26852 46676 26908 46844
rect 38612 46788 38668 46844
rect 32498 46732 32508 46788
rect 32564 46732 38668 46788
rect 38770 46732 38780 46788
rect 38836 46732 40460 46788
rect 40516 46732 40908 46788
rect 40964 46732 40974 46788
rect 45602 46732 45612 46788
rect 45668 46732 46060 46788
rect 46116 46732 46126 46788
rect 48178 46732 48188 46788
rect 48244 46732 49532 46788
rect 49588 46732 51436 46788
rect 51492 46732 51502 46788
rect 55570 46732 55580 46788
rect 55636 46732 57260 46788
rect 57316 46732 57326 46788
rect 57586 46732 57596 46788
rect 57652 46732 61740 46788
rect 61796 46732 61806 46788
rect 3826 46620 3836 46676
rect 3892 46620 3902 46676
rect 4050 46620 4060 46676
rect 4116 46620 4154 46676
rect 9538 46620 9548 46676
rect 9604 46620 11788 46676
rect 11844 46620 11854 46676
rect 14690 46620 14700 46676
rect 14756 46620 16156 46676
rect 16212 46620 16222 46676
rect 17378 46620 17388 46676
rect 17444 46620 18340 46676
rect 21746 46620 21756 46676
rect 21812 46620 23324 46676
rect 23380 46620 23390 46676
rect 24322 46620 24332 46676
rect 24388 46620 26236 46676
rect 26292 46620 26302 46676
rect 26852 46620 27804 46676
rect 27860 46620 29932 46676
rect 29988 46620 29998 46676
rect 41682 46620 41692 46676
rect 41748 46620 44828 46676
rect 44884 46620 44894 46676
rect 48038 46620 48076 46676
rect 48132 46620 48748 46676
rect 48804 46620 48814 46676
rect 61366 46620 61404 46676
rect 61460 46620 61470 46676
rect 3836 46564 3892 46620
rect 18284 46564 18340 46620
rect 3836 46508 14252 46564
rect 14308 46508 15036 46564
rect 15092 46508 15102 46564
rect 16258 46508 16268 46564
rect 16324 46508 17724 46564
rect 17780 46508 17790 46564
rect 18274 46508 18284 46564
rect 18340 46508 21308 46564
rect 21364 46508 32788 46564
rect 34962 46508 34972 46564
rect 35028 46508 40796 46564
rect 40852 46508 40862 46564
rect 43362 46508 43372 46564
rect 43428 46508 44940 46564
rect 44996 46508 45724 46564
rect 45780 46508 45790 46564
rect 53778 46508 53788 46564
rect 53844 46508 54796 46564
rect 54852 46508 57540 46564
rect 61282 46508 61292 46564
rect 61348 46508 62860 46564
rect 62916 46508 62926 46564
rect 32732 46452 32788 46508
rect 57484 46452 57540 46508
rect 4498 46396 4508 46452
rect 4564 46396 11452 46452
rect 11508 46396 11518 46452
rect 15362 46396 15372 46452
rect 15428 46396 21420 46452
rect 21476 46396 21486 46452
rect 32732 46396 35756 46452
rect 35812 46396 35822 46452
rect 38994 46396 39004 46452
rect 39060 46396 41132 46452
rect 41188 46396 41198 46452
rect 50418 46396 50428 46452
rect 50484 46396 50988 46452
rect 51044 46396 51054 46452
rect 54338 46396 54348 46452
rect 54404 46396 55020 46452
rect 55076 46396 55086 46452
rect 55234 46396 55244 46452
rect 55300 46396 57260 46452
rect 57316 46396 57326 46452
rect 57484 46396 62636 46452
rect 62692 46396 62702 46452
rect 16706 46284 16716 46340
rect 16772 46284 19404 46340
rect 19460 46284 26908 46340
rect 42018 46284 42028 46340
rect 42084 46284 44940 46340
rect 44996 46284 45006 46340
rect 51874 46284 51884 46340
rect 51940 46284 52668 46340
rect 52724 46284 52734 46340
rect 58370 46284 58380 46340
rect 58436 46284 61516 46340
rect 61572 46284 61582 46340
rect 61730 46284 61740 46340
rect 61796 46284 61834 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 22082 46172 22092 46228
rect 22148 46172 23884 46228
rect 23940 46172 23950 46228
rect 26852 46116 26908 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 27878 46172 27916 46228
rect 27972 46172 27982 46228
rect 30370 46172 30380 46228
rect 30436 46172 34636 46228
rect 34692 46172 34702 46228
rect 51202 46172 51212 46228
rect 51268 46172 53340 46228
rect 53396 46172 55580 46228
rect 55636 46172 55646 46228
rect 58706 46172 58716 46228
rect 58772 46172 62076 46228
rect 62132 46172 62142 46228
rect 2706 46060 2716 46116
rect 2772 46060 3612 46116
rect 3668 46060 3678 46116
rect 10994 46060 11004 46116
rect 11060 46060 11452 46116
rect 11508 46060 11518 46116
rect 13906 46060 13916 46116
rect 13972 46060 14252 46116
rect 14308 46060 14318 46116
rect 16818 46060 16828 46116
rect 16884 46060 18172 46116
rect 18228 46060 18844 46116
rect 18900 46060 18910 46116
rect 23762 46060 23772 46116
rect 23828 46060 24780 46116
rect 24836 46060 24846 46116
rect 26852 46060 27468 46116
rect 27524 46060 27534 46116
rect 33478 46060 33516 46116
rect 33572 46060 33582 46116
rect 33730 46060 33740 46116
rect 33796 46060 39676 46116
rect 39732 46060 39742 46116
rect 45154 46060 45164 46116
rect 45220 46060 46732 46116
rect 46788 46060 50036 46116
rect 50306 46060 50316 46116
rect 50372 46060 50764 46116
rect 50820 46060 51436 46116
rect 51492 46060 51502 46116
rect 49980 46004 50036 46060
rect 2370 45948 2380 46004
rect 2436 45948 5740 46004
rect 5796 45948 6748 46004
rect 6804 45948 6814 46004
rect 8754 45948 8764 46004
rect 8820 45948 11340 46004
rect 11396 45948 11406 46004
rect 11666 45948 11676 46004
rect 11732 45948 12572 46004
rect 12628 45948 13020 46004
rect 13076 45948 13086 46004
rect 17602 45948 17612 46004
rect 17668 45948 18956 46004
rect 19012 45948 19022 46004
rect 20066 45948 20076 46004
rect 20132 45948 40068 46004
rect 42102 45948 42140 46004
rect 42196 45948 42206 46004
rect 44930 45948 44940 46004
rect 44996 45948 47516 46004
rect 47572 45948 47582 46004
rect 49186 45948 49196 46004
rect 49252 45948 49756 46004
rect 49812 45948 49822 46004
rect 49980 45948 50428 46004
rect 50484 45948 51548 46004
rect 51604 45948 51614 46004
rect 59602 45948 59612 46004
rect 59668 45948 60620 46004
rect 60676 45948 60686 46004
rect 3602 45836 3612 45892
rect 3668 45836 4172 45892
rect 4228 45836 6300 45892
rect 6356 45836 6366 45892
rect 10098 45836 10108 45892
rect 10164 45836 13468 45892
rect 13524 45836 13534 45892
rect 15092 45780 15148 45892
rect 15204 45836 15214 45892
rect 17714 45836 17724 45892
rect 17780 45836 18620 45892
rect 18676 45836 18686 45892
rect 20402 45836 20412 45892
rect 20468 45836 20860 45892
rect 20916 45836 20926 45892
rect 23986 45836 23996 45892
rect 24052 45836 24556 45892
rect 24612 45836 24622 45892
rect 26002 45836 26012 45892
rect 26068 45836 26796 45892
rect 26852 45836 28924 45892
rect 28980 45836 28990 45892
rect 29474 45836 29484 45892
rect 29540 45836 29932 45892
rect 29988 45836 29998 45892
rect 31154 45836 31164 45892
rect 31220 45836 33292 45892
rect 33348 45836 33358 45892
rect 33618 45836 33628 45892
rect 33684 45836 35196 45892
rect 35252 45836 36316 45892
rect 36372 45836 36382 45892
rect 24556 45780 24612 45836
rect 40012 45780 40068 45948
rect 46946 45836 46956 45892
rect 47012 45836 47852 45892
rect 47908 45836 47918 45892
rect 50082 45836 50092 45892
rect 50148 45836 51212 45892
rect 51268 45836 51278 45892
rect 53330 45836 53340 45892
rect 53396 45836 53452 45892
rect 53508 45836 53518 45892
rect 57922 45836 57932 45892
rect 57988 45836 60844 45892
rect 60900 45836 60910 45892
rect 61254 45836 61292 45892
rect 61348 45836 61358 45892
rect 62150 45836 62188 45892
rect 62244 45836 62254 45892
rect 47852 45780 47908 45836
rect 2594 45724 2604 45780
rect 2660 45724 6748 45780
rect 6804 45724 6814 45780
rect 10770 45724 10780 45780
rect 10836 45724 11228 45780
rect 11284 45724 11294 45780
rect 12898 45724 12908 45780
rect 12964 45724 15148 45780
rect 17266 45724 17276 45780
rect 17332 45724 17612 45780
rect 17668 45724 19740 45780
rect 19796 45724 19806 45780
rect 24556 45724 25788 45780
rect 25844 45724 26908 45780
rect 26964 45724 26974 45780
rect 30930 45724 30940 45780
rect 30996 45724 31006 45780
rect 32162 45724 32172 45780
rect 32228 45724 33068 45780
rect 33124 45724 33964 45780
rect 34020 45724 34030 45780
rect 38210 45724 38220 45780
rect 38276 45724 39004 45780
rect 39060 45724 39070 45780
rect 40012 45724 41692 45780
rect 41748 45724 43820 45780
rect 43876 45724 43886 45780
rect 45378 45724 45388 45780
rect 45444 45724 47068 45780
rect 47124 45724 47134 45780
rect 47852 45724 50988 45780
rect 51044 45724 51054 45780
rect 51986 45724 51996 45780
rect 52052 45724 54684 45780
rect 54740 45724 54750 45780
rect 30940 45668 30996 45724
rect 3332 45612 4844 45668
rect 4900 45612 4910 45668
rect 8978 45612 8988 45668
rect 9044 45612 9660 45668
rect 9716 45612 9726 45668
rect 11442 45612 11452 45668
rect 11508 45612 11788 45668
rect 11844 45612 12012 45668
rect 12068 45612 12796 45668
rect 12852 45612 12862 45668
rect 17388 45612 18060 45668
rect 18116 45612 20076 45668
rect 20132 45612 20142 45668
rect 20822 45612 20860 45668
rect 20916 45612 20926 45668
rect 23202 45612 23212 45668
rect 23268 45612 26012 45668
rect 26068 45612 26078 45668
rect 26786 45612 26796 45668
rect 26852 45612 30996 45668
rect 32386 45612 32396 45668
rect 32452 45612 34300 45668
rect 34356 45612 34860 45668
rect 34916 45612 34926 45668
rect 44258 45612 44268 45668
rect 44324 45612 44828 45668
rect 44884 45612 44894 45668
rect 48290 45612 48300 45668
rect 48356 45612 51884 45668
rect 51940 45612 51950 45668
rect 58930 45612 58940 45668
rect 58996 45612 61628 45668
rect 61684 45612 61694 45668
rect 3332 45556 3388 45612
rect 17388 45556 17444 45612
rect 1138 45500 1148 45556
rect 1204 45500 3388 45556
rect 4274 45500 4284 45556
rect 4340 45500 4788 45556
rect 9762 45500 9772 45556
rect 9828 45500 13020 45556
rect 13076 45500 13086 45556
rect 17378 45500 17388 45556
rect 17444 45500 17454 45556
rect 23874 45500 23884 45556
rect 23940 45500 25340 45556
rect 25396 45500 25406 45556
rect 26226 45500 26236 45556
rect 26292 45500 26684 45556
rect 26740 45500 26750 45556
rect 30258 45500 30268 45556
rect 30324 45500 31388 45556
rect 31444 45500 32844 45556
rect 32900 45500 32910 45556
rect 34626 45500 34636 45556
rect 34692 45500 37548 45556
rect 37604 45500 37614 45556
rect 42130 45500 42140 45556
rect 42196 45500 43260 45556
rect 43316 45500 43326 45556
rect 44370 45500 44380 45556
rect 44436 45500 44446 45556
rect 50082 45500 50092 45556
rect 50148 45500 50204 45556
rect 50260 45500 50270 45556
rect 53302 45500 53340 45556
rect 53396 45500 53406 45556
rect 53554 45500 53564 45556
rect 53620 45500 53630 45556
rect 4732 45444 4788 45500
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 2706 45388 2716 45444
rect 2772 45388 4508 45444
rect 4564 45388 4574 45444
rect 4732 45388 14028 45444
rect 14084 45388 14924 45444
rect 14980 45388 14990 45444
rect 21410 45388 21420 45444
rect 21476 45388 27132 45444
rect 27188 45388 29260 45444
rect 29316 45388 29326 45444
rect 29474 45388 29484 45444
rect 29540 45388 30380 45444
rect 30436 45388 30446 45444
rect 35522 45388 35532 45444
rect 35588 45388 40236 45444
rect 40292 45388 40302 45444
rect 42140 45332 42196 45500
rect 43894 45388 43932 45444
rect 43988 45388 43998 45444
rect 44380 45332 44436 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 51538 45388 51548 45444
rect 51604 45388 51884 45444
rect 51940 45388 51950 45444
rect 5964 45276 7308 45332
rect 7364 45276 8204 45332
rect 8260 45276 8270 45332
rect 8418 45276 8428 45332
rect 8484 45276 13804 45332
rect 13860 45276 13870 45332
rect 20514 45276 20524 45332
rect 20580 45276 23324 45332
rect 23380 45276 23390 45332
rect 24098 45276 24108 45332
rect 24164 45276 24780 45332
rect 24836 45276 25116 45332
rect 25172 45276 25182 45332
rect 25414 45276 25452 45332
rect 25508 45276 25518 45332
rect 25666 45276 25676 45332
rect 25732 45276 25770 45332
rect 33394 45276 33404 45332
rect 33460 45276 35196 45332
rect 35252 45276 35262 45332
rect 35410 45276 35420 45332
rect 35476 45276 42196 45332
rect 43250 45276 43260 45332
rect 43316 45276 44436 45332
rect 53564 45332 53620 45500
rect 53564 45276 56924 45332
rect 56980 45276 56990 45332
rect 3154 45164 3164 45220
rect 3220 45164 3388 45220
rect 3444 45164 4060 45220
rect 4116 45164 4126 45220
rect 5964 45108 6020 45276
rect 6626 45164 6636 45220
rect 6692 45164 7420 45220
rect 7476 45164 7486 45220
rect 10546 45164 10556 45220
rect 10612 45164 12348 45220
rect 12404 45164 14700 45220
rect 14756 45164 14766 45220
rect 21970 45164 21980 45220
rect 22036 45164 25900 45220
rect 25956 45164 25966 45220
rect 26562 45164 26572 45220
rect 26628 45164 28252 45220
rect 28308 45164 28318 45220
rect 32620 45164 35644 45220
rect 35700 45164 35710 45220
rect 35858 45164 35868 45220
rect 35924 45164 41132 45220
rect 41188 45164 41198 45220
rect 43362 45164 43372 45220
rect 43428 45164 43820 45220
rect 43876 45164 43886 45220
rect 45154 45164 45164 45220
rect 45220 45164 47628 45220
rect 47684 45164 48188 45220
rect 48244 45164 48254 45220
rect 48738 45164 48748 45220
rect 48804 45164 48860 45220
rect 48916 45164 48926 45220
rect 49522 45164 49532 45220
rect 49588 45164 49868 45220
rect 49924 45164 49934 45220
rect 55906 45164 55916 45220
rect 55972 45164 57708 45220
rect 57764 45164 57774 45220
rect 61618 45164 61628 45220
rect 61684 45164 62636 45220
rect 62692 45164 62702 45220
rect 1698 45052 1708 45108
rect 1764 45052 3052 45108
rect 3108 45052 3118 45108
rect 3378 45052 3388 45108
rect 3444 45052 4172 45108
rect 4228 45052 4238 45108
rect 4610 45052 4620 45108
rect 4676 45052 5964 45108
rect 6020 45052 6030 45108
rect 6514 45052 6524 45108
rect 6580 45052 8764 45108
rect 8820 45052 9548 45108
rect 9604 45052 9614 45108
rect 10770 45052 10780 45108
rect 10836 45052 11564 45108
rect 11620 45052 11630 45108
rect 14130 45052 14140 45108
rect 14196 45052 15372 45108
rect 15428 45052 15438 45108
rect 15586 45052 15596 45108
rect 15652 45052 15764 45108
rect 18050 45052 18060 45108
rect 18116 45052 20188 45108
rect 20244 45052 20254 45108
rect 20626 45052 20636 45108
rect 20692 45052 23100 45108
rect 23156 45052 23166 45108
rect 23426 45052 23436 45108
rect 23492 45052 23996 45108
rect 24052 45052 24062 45108
rect 24658 45052 24668 45108
rect 24724 45052 27020 45108
rect 27076 45052 27086 45108
rect 15708 44996 15764 45052
rect 4834 44940 4844 44996
rect 4900 44940 15484 44996
rect 15540 44940 15550 44996
rect 15708 44940 22652 44996
rect 22708 44940 22718 44996
rect 26002 44940 26012 44996
rect 26068 44940 30156 44996
rect 30212 44940 30222 44996
rect 32620 44884 32676 45164
rect 35644 45108 35700 45164
rect 32834 45052 32844 45108
rect 32900 45052 33740 45108
rect 33796 45052 34636 45108
rect 34692 45052 34702 45108
rect 35410 45052 35420 45108
rect 35476 45052 35486 45108
rect 35644 45052 36316 45108
rect 36372 45052 36876 45108
rect 36932 45052 36942 45108
rect 37202 45052 37212 45108
rect 37268 45052 38780 45108
rect 38836 45052 38846 45108
rect 39218 45052 39228 45108
rect 39284 45052 40348 45108
rect 40404 45052 40414 45108
rect 44482 45052 44492 45108
rect 44548 45052 47740 45108
rect 47796 45052 47806 45108
rect 48962 45052 48972 45108
rect 49028 45052 50316 45108
rect 33394 44940 33404 44996
rect 33460 44940 33964 44996
rect 34020 44940 34860 44996
rect 34916 44940 34926 44996
rect 35420 44884 35476 45052
rect 39228 44996 39284 45052
rect 50372 44996 50428 45108
rect 51090 45052 51100 45108
rect 51156 45052 53228 45108
rect 53284 45052 53294 45108
rect 53666 45052 53676 45108
rect 53732 45052 54684 45108
rect 54740 45052 55132 45108
rect 55188 45052 55198 45108
rect 59826 45052 59836 45108
rect 59892 45052 61404 45108
rect 61460 45052 61470 45108
rect 37090 44940 37100 44996
rect 37156 44940 39284 44996
rect 40226 44940 40236 44996
rect 40292 44940 41468 44996
rect 41524 44940 41534 44996
rect 43138 44940 43148 44996
rect 43204 44940 44716 44996
rect 44772 44940 47180 44996
rect 47236 44940 47246 44996
rect 50372 44940 52668 44996
rect 52724 44940 52734 44996
rect 55542 44940 55580 44996
rect 55636 44940 55646 44996
rect 55906 44940 55916 44996
rect 55972 44940 60284 44996
rect 60340 44940 60350 44996
rect 55580 44884 55636 44940
rect 5730 44828 5740 44884
rect 5796 44828 7084 44884
rect 7140 44828 7150 44884
rect 11554 44828 11564 44884
rect 11620 44828 16492 44884
rect 16548 44828 16558 44884
rect 16706 44828 16716 44884
rect 16772 44828 32676 44884
rect 32732 44828 35476 44884
rect 37986 44828 37996 44884
rect 38052 44828 39900 44884
rect 39956 44828 39966 44884
rect 55580 44828 57932 44884
rect 57988 44828 57998 44884
rect 58818 44828 58828 44884
rect 58884 44828 62076 44884
rect 62132 44828 62142 44884
rect 32732 44772 32788 44828
rect 15026 44716 15036 44772
rect 15092 44716 22876 44772
rect 22932 44716 25676 44772
rect 25732 44716 25742 44772
rect 25890 44716 25900 44772
rect 25956 44716 32788 44772
rect 38098 44716 38108 44772
rect 38164 44716 43988 44772
rect 46050 44716 46060 44772
rect 46116 44716 47404 44772
rect 47460 44716 47964 44772
rect 48020 44716 48030 44772
rect 54562 44716 54572 44772
rect 54628 44716 58156 44772
rect 58212 44716 60620 44772
rect 60676 44716 60686 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 18610 44604 18620 44660
rect 18676 44604 23548 44660
rect 23604 44604 24780 44660
rect 24836 44604 24846 44660
rect 25414 44604 25452 44660
rect 25508 44604 25518 44660
rect 26226 44604 26236 44660
rect 26292 44604 31164 44660
rect 31220 44604 31230 44660
rect 40114 44604 40124 44660
rect 40180 44604 43764 44660
rect 43708 44548 43764 44604
rect 43932 44548 43988 44716
rect 53330 44604 53340 44660
rect 53396 44604 56588 44660
rect 56644 44604 56654 44660
rect 5506 44492 5516 44548
rect 5572 44492 6076 44548
rect 6132 44492 9324 44548
rect 9380 44492 10332 44548
rect 10388 44492 10398 44548
rect 16258 44492 16268 44548
rect 16324 44492 35812 44548
rect 36530 44492 36540 44548
rect 36596 44492 37436 44548
rect 37492 44492 37502 44548
rect 37874 44492 37884 44548
rect 37940 44492 39676 44548
rect 39732 44492 39742 44548
rect 40338 44492 40348 44548
rect 40404 44492 41300 44548
rect 43670 44492 43708 44548
rect 43764 44492 43774 44548
rect 43922 44492 43932 44548
rect 43988 44492 43998 44548
rect 48850 44492 48860 44548
rect 48916 44492 49756 44548
rect 49812 44492 49822 44548
rect 53106 44492 53116 44548
rect 53172 44492 54460 44548
rect 54516 44492 54526 44548
rect 0 44436 800 44464
rect 0 44380 1876 44436
rect 3490 44380 3500 44436
rect 3556 44380 4620 44436
rect 4676 44380 5740 44436
rect 5796 44380 5806 44436
rect 6290 44380 6300 44436
rect 6356 44380 7868 44436
rect 7924 44380 8316 44436
rect 8372 44380 10220 44436
rect 10276 44380 10286 44436
rect 11330 44380 11340 44436
rect 11396 44380 12236 44436
rect 12292 44380 12302 44436
rect 21746 44380 21756 44436
rect 21812 44380 24556 44436
rect 24612 44380 25116 44436
rect 25172 44380 25182 44436
rect 27794 44380 27804 44436
rect 27860 44380 29036 44436
rect 29092 44380 29102 44436
rect 34402 44380 34412 44436
rect 34468 44380 34860 44436
rect 34916 44380 34926 44436
rect 0 44352 800 44380
rect 1820 44324 1876 44380
rect 1810 44268 1820 44324
rect 1876 44268 2268 44324
rect 2324 44268 2334 44324
rect 2594 44268 2604 44324
rect 2660 44268 3388 44324
rect 3444 44268 4396 44324
rect 4452 44268 4462 44324
rect 7186 44268 7196 44324
rect 7252 44268 8540 44324
rect 8596 44268 8606 44324
rect 10854 44268 10892 44324
rect 10948 44268 10958 44324
rect 16370 44268 16380 44324
rect 16436 44268 17388 44324
rect 17444 44268 20524 44324
rect 20580 44268 20590 44324
rect 22306 44268 22316 44324
rect 22372 44268 23212 44324
rect 23268 44268 23660 44324
rect 23716 44268 23726 44324
rect 24098 44268 24108 44324
rect 24164 44268 24444 44324
rect 24500 44268 24510 44324
rect 24882 44268 24892 44324
rect 24948 44268 25340 44324
rect 25396 44268 25406 44324
rect 33282 44268 33292 44324
rect 33348 44268 33628 44324
rect 33684 44268 34300 44324
rect 34356 44268 34366 44324
rect 35756 44212 35812 44492
rect 41244 44436 41300 44492
rect 39554 44380 39564 44436
rect 39620 44380 40124 44436
rect 40180 44380 41020 44436
rect 41076 44380 41086 44436
rect 41244 44380 46172 44436
rect 46228 44380 46238 44436
rect 50642 44380 50652 44436
rect 50708 44380 50718 44436
rect 53974 44380 54012 44436
rect 54068 44380 54078 44436
rect 55906 44380 55916 44436
rect 55972 44380 56476 44436
rect 56532 44380 56542 44436
rect 36194 44268 36204 44324
rect 36260 44268 37324 44324
rect 37380 44268 38108 44324
rect 38164 44268 38174 44324
rect 43138 44268 43148 44324
rect 43204 44268 44940 44324
rect 44996 44268 45006 44324
rect 48066 44268 48076 44324
rect 48132 44268 50428 44324
rect 50484 44268 50494 44324
rect 50652 44212 50708 44380
rect 54898 44268 54908 44324
rect 54964 44268 57036 44324
rect 57092 44268 60844 44324
rect 60900 44268 60910 44324
rect 2034 44156 2044 44212
rect 2100 44156 2380 44212
rect 2436 44156 3052 44212
rect 3108 44156 4172 44212
rect 4228 44156 4238 44212
rect 26450 44156 26460 44212
rect 26516 44156 27804 44212
rect 27860 44156 27870 44212
rect 35756 44156 36988 44212
rect 37044 44156 37884 44212
rect 37940 44156 37950 44212
rect 38612 44156 42812 44212
rect 42868 44156 42878 44212
rect 44370 44156 44380 44212
rect 44436 44156 45388 44212
rect 45444 44156 45454 44212
rect 49634 44156 49644 44212
rect 49700 44156 54012 44212
rect 54068 44156 54078 44212
rect 56242 44156 56252 44212
rect 56308 44156 56812 44212
rect 56868 44156 57596 44212
rect 57652 44156 57662 44212
rect 38612 44100 38668 44156
rect 3266 44044 3276 44100
rect 3332 44044 4060 44100
rect 4116 44044 4126 44100
rect 10210 44044 10220 44100
rect 10276 44044 19516 44100
rect 19572 44044 20524 44100
rect 20580 44044 20590 44100
rect 28662 44044 28700 44100
rect 28756 44044 28766 44100
rect 29026 44044 29036 44100
rect 29092 44044 30156 44100
rect 30212 44044 30222 44100
rect 37538 44044 37548 44100
rect 37604 44044 38668 44100
rect 47954 44044 47964 44100
rect 48020 44044 48748 44100
rect 48804 44044 48814 44100
rect 50642 44044 50652 44100
rect 50708 44044 52948 44100
rect 53890 44044 53900 44100
rect 53956 44044 55580 44100
rect 55636 44044 55646 44100
rect 52892 43988 52948 44044
rect 26852 43932 41356 43988
rect 41412 43932 41422 43988
rect 52882 43932 52892 43988
rect 52948 43932 53564 43988
rect 53620 43932 53630 43988
rect 53778 43932 53788 43988
rect 53844 43932 55356 43988
rect 55412 43932 55422 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 3798 43820 3836 43876
rect 3892 43820 3902 43876
rect 20290 43820 20300 43876
rect 20356 43820 20636 43876
rect 20692 43820 20702 43876
rect 26852 43764 26908 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 12450 43708 12460 43764
rect 12516 43708 14140 43764
rect 14196 43708 14206 43764
rect 15092 43708 26908 43764
rect 27132 43820 30268 43876
rect 30324 43820 30334 43876
rect 40114 43820 40124 43876
rect 40180 43820 41580 43876
rect 41636 43820 41646 43876
rect 44818 43820 44828 43876
rect 44884 43820 44894 43876
rect 48710 43820 48748 43876
rect 48804 43820 48814 43876
rect 53218 43820 53228 43876
rect 53284 43820 54236 43876
rect 54292 43820 54796 43876
rect 54852 43820 54862 43876
rect 56662 43820 56700 43876
rect 56756 43820 56766 43876
rect 15092 43652 15148 43708
rect 6402 43596 6412 43652
rect 6468 43596 7084 43652
rect 7140 43596 7150 43652
rect 8866 43596 8876 43652
rect 8932 43596 9100 43652
rect 9156 43596 9660 43652
rect 9716 43596 9726 43652
rect 9874 43596 9884 43652
rect 9940 43596 12796 43652
rect 12852 43596 12862 43652
rect 14690 43596 14700 43652
rect 14756 43596 15148 43652
rect 16146 43596 16156 43652
rect 16212 43596 19068 43652
rect 19124 43596 19134 43652
rect 19842 43596 19852 43652
rect 19908 43596 21756 43652
rect 21812 43596 21822 43652
rect 22978 43596 22988 43652
rect 23044 43596 23212 43652
rect 23268 43596 26908 43652
rect 26852 43540 26908 43596
rect 27132 43540 27188 43820
rect 29810 43708 29820 43764
rect 29876 43708 30380 43764
rect 30436 43708 30446 43764
rect 34402 43708 34412 43764
rect 34468 43708 35308 43764
rect 35364 43708 35374 43764
rect 42242 43708 42252 43764
rect 42308 43708 44268 43764
rect 44324 43708 44334 43764
rect 44828 43652 44884 43820
rect 48178 43708 48188 43764
rect 48244 43708 49196 43764
rect 49252 43708 49262 43764
rect 51986 43708 51996 43764
rect 52052 43708 52780 43764
rect 52836 43708 52846 43764
rect 54338 43708 54348 43764
rect 54404 43708 60620 43764
rect 60676 43708 60686 43764
rect 30594 43596 30604 43652
rect 30660 43596 33068 43652
rect 33124 43596 33134 43652
rect 36866 43596 36876 43652
rect 36932 43596 37772 43652
rect 37828 43596 37838 43652
rect 38434 43596 38444 43652
rect 38500 43596 40908 43652
rect 40964 43596 40974 43652
rect 43474 43596 43484 43652
rect 43540 43596 43820 43652
rect 43876 43596 43886 43652
rect 44828 43596 46732 43652
rect 46788 43596 46798 43652
rect 47842 43596 47852 43652
rect 47908 43596 48524 43652
rect 48580 43596 49308 43652
rect 49364 43596 50204 43652
rect 50260 43596 50270 43652
rect 54002 43596 54012 43652
rect 54068 43596 55804 43652
rect 55860 43596 55870 43652
rect 57810 43596 57820 43652
rect 57876 43596 58716 43652
rect 58772 43596 61516 43652
rect 61572 43596 61582 43652
rect 6626 43484 6636 43540
rect 6692 43484 8988 43540
rect 9044 43484 9548 43540
rect 9604 43484 9996 43540
rect 10052 43484 10062 43540
rect 10994 43484 11004 43540
rect 11060 43484 11676 43540
rect 11732 43484 11742 43540
rect 15092 43484 18508 43540
rect 18564 43484 18574 43540
rect 18722 43484 18732 43540
rect 18788 43484 19516 43540
rect 19572 43484 19582 43540
rect 20290 43484 20300 43540
rect 20356 43484 21868 43540
rect 21924 43484 21934 43540
rect 22082 43484 22092 43540
rect 22148 43484 26124 43540
rect 26180 43484 26190 43540
rect 26852 43484 27188 43540
rect 27794 43484 27804 43540
rect 27860 43484 29372 43540
rect 29428 43484 29438 43540
rect 29586 43484 29596 43540
rect 29652 43484 30044 43540
rect 30100 43484 30110 43540
rect 31042 43484 31052 43540
rect 31108 43484 32060 43540
rect 32116 43484 32126 43540
rect 34290 43484 34300 43540
rect 34356 43484 36652 43540
rect 36708 43484 36718 43540
rect 37650 43484 37660 43540
rect 37716 43484 38556 43540
rect 38612 43484 38622 43540
rect 39106 43484 39116 43540
rect 39172 43484 40796 43540
rect 40852 43484 41692 43540
rect 41748 43484 42252 43540
rect 42308 43484 42318 43540
rect 42914 43484 42924 43540
rect 42980 43484 43596 43540
rect 43652 43484 44156 43540
rect 44212 43484 44222 43540
rect 50754 43484 50764 43540
rect 50820 43484 51772 43540
rect 51828 43484 52892 43540
rect 52948 43484 52958 43540
rect 55010 43484 55020 43540
rect 55076 43484 57260 43540
rect 57316 43484 57326 43540
rect 61926 43484 61964 43540
rect 62020 43484 62030 43540
rect 15092 43428 15148 43484
rect 29372 43428 29428 43484
rect 4134 43372 4172 43428
rect 4228 43372 4238 43428
rect 7074 43372 7084 43428
rect 7140 43372 10108 43428
rect 10164 43372 15148 43428
rect 17938 43372 17948 43428
rect 18004 43372 20636 43428
rect 20692 43372 20702 43428
rect 21196 43372 24556 43428
rect 24612 43372 24622 43428
rect 25442 43372 25452 43428
rect 25508 43372 26236 43428
rect 26292 43372 26302 43428
rect 27906 43372 27916 43428
rect 27972 43372 28028 43428
rect 28084 43372 28364 43428
rect 28420 43372 28430 43428
rect 29372 43372 31500 43428
rect 31556 43372 31566 43428
rect 46946 43372 46956 43428
rect 47012 43372 47180 43428
rect 47236 43372 49308 43428
rect 49364 43372 51324 43428
rect 51380 43372 51390 43428
rect 3714 43260 3724 43316
rect 3780 43260 4508 43316
rect 4564 43260 4574 43316
rect 6290 43260 6300 43316
rect 6356 43260 8876 43316
rect 8932 43260 8942 43316
rect 18386 43260 18396 43316
rect 18452 43260 19292 43316
rect 19348 43260 19358 43316
rect 21196 43204 21252 43372
rect 23492 43260 24108 43316
rect 24164 43260 24668 43316
rect 24724 43260 26796 43316
rect 26852 43260 26862 43316
rect 27570 43260 27580 43316
rect 27636 43260 27916 43316
rect 27972 43260 27982 43316
rect 29922 43260 29932 43316
rect 29988 43260 31164 43316
rect 31220 43260 31230 43316
rect 53554 43260 53564 43316
rect 53620 43260 53900 43316
rect 53956 43260 59276 43316
rect 59332 43260 59342 43316
rect 61954 43260 61964 43316
rect 62020 43260 62030 43316
rect 23492 43204 23548 43260
rect 7186 43148 7196 43204
rect 7252 43148 7532 43204
rect 7588 43148 21252 43204
rect 21308 43148 23548 43204
rect 38098 43148 38108 43204
rect 38164 43148 40236 43204
rect 40292 43148 40302 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 21308 43092 21364 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 61964 43092 62020 43260
rect 63200 43092 64000 43120
rect 13010 43036 13020 43092
rect 13076 43036 15148 43092
rect 18498 43036 18508 43092
rect 18564 43036 21364 43092
rect 21522 43036 21532 43092
rect 21588 43036 23772 43092
rect 23828 43036 23838 43092
rect 30594 43036 30604 43092
rect 30660 43036 34076 43092
rect 34132 43036 34142 43092
rect 39890 43036 39900 43092
rect 39956 43036 41132 43092
rect 41188 43036 41198 43092
rect 49074 43036 49084 43092
rect 49140 43036 52780 43092
rect 52836 43036 53900 43092
rect 53956 43036 55916 43092
rect 55972 43036 55982 43092
rect 61964 43036 64000 43092
rect 2146 42924 2156 42980
rect 2212 42924 2492 42980
rect 2548 42924 2558 42980
rect 3714 42924 3724 42980
rect 3780 42924 4172 42980
rect 4228 42924 4238 42980
rect 15092 42924 15148 43036
rect 63200 43008 64000 43036
rect 15204 42924 15242 42980
rect 15362 42924 15372 42980
rect 15428 42924 19516 42980
rect 19572 42924 19582 42980
rect 21970 42924 21980 42980
rect 22036 42924 22652 42980
rect 22708 42924 23996 42980
rect 24052 42924 24062 42980
rect 30482 42924 30492 42980
rect 30548 42924 31388 42980
rect 31444 42924 41020 42980
rect 41076 42924 41086 42980
rect 50372 42924 51212 42980
rect 51268 42924 53452 42980
rect 53508 42924 53518 42980
rect 53778 42924 53788 42980
rect 53844 42924 56364 42980
rect 56420 42924 57372 42980
rect 57428 42924 57438 42980
rect 4610 42812 4620 42868
rect 4676 42812 5740 42868
rect 5796 42812 7980 42868
rect 8036 42812 8316 42868
rect 8372 42812 8382 42868
rect 10780 42812 26908 42868
rect 26964 42812 26974 42868
rect 29698 42812 29708 42868
rect 29764 42812 31836 42868
rect 31892 42812 31902 42868
rect 32050 42812 32060 42868
rect 32116 42812 32508 42868
rect 32564 42812 32574 42868
rect 5954 42700 5964 42756
rect 6020 42700 10556 42756
rect 10612 42700 10622 42756
rect 10780 42644 10836 42812
rect 14242 42700 14252 42756
rect 14308 42700 14588 42756
rect 14644 42700 14654 42756
rect 17602 42700 17612 42756
rect 17668 42700 17948 42756
rect 18004 42700 18014 42756
rect 21186 42700 21196 42756
rect 21252 42700 21532 42756
rect 21588 42700 21598 42756
rect 23090 42700 23100 42756
rect 23156 42700 25228 42756
rect 25284 42700 25294 42756
rect 37874 42700 37884 42756
rect 37940 42700 38892 42756
rect 38948 42700 38958 42756
rect 40226 42700 40236 42756
rect 40292 42700 42140 42756
rect 42196 42700 42206 42756
rect 50372 42644 50428 42924
rect 51762 42812 51772 42868
rect 51828 42812 54572 42868
rect 54628 42812 56028 42868
rect 56084 42812 56094 42868
rect 56466 42812 56476 42868
rect 56532 42812 57036 42868
rect 57092 42812 57102 42868
rect 60946 42812 60956 42868
rect 61012 42812 61516 42868
rect 61572 42812 61582 42868
rect 51538 42700 51548 42756
rect 51604 42700 52108 42756
rect 52164 42700 52892 42756
rect 52948 42700 52958 42756
rect 53442 42700 53452 42756
rect 53508 42700 55916 42756
rect 55972 42700 60060 42756
rect 60116 42700 60126 42756
rect 61282 42700 61292 42756
rect 61348 42700 61628 42756
rect 61684 42700 61694 42756
rect 2146 42588 2156 42644
rect 2212 42588 2492 42644
rect 2548 42588 3388 42644
rect 3444 42588 4060 42644
rect 4116 42588 4844 42644
rect 4900 42588 4910 42644
rect 9874 42588 9884 42644
rect 9940 42588 10332 42644
rect 10388 42588 10836 42644
rect 12002 42588 12012 42644
rect 12068 42588 12796 42644
rect 12852 42588 13692 42644
rect 13748 42588 13758 42644
rect 15250 42588 15260 42644
rect 15316 42588 23436 42644
rect 23492 42588 23502 42644
rect 28802 42588 28812 42644
rect 28868 42588 29708 42644
rect 29764 42588 29774 42644
rect 31154 42588 31164 42644
rect 31220 42588 32172 42644
rect 32228 42588 32620 42644
rect 32676 42588 35308 42644
rect 35364 42588 35374 42644
rect 38546 42588 38556 42644
rect 38612 42588 39340 42644
rect 39396 42588 39406 42644
rect 44370 42588 44380 42644
rect 44436 42588 50428 42644
rect 3266 42476 3276 42532
rect 3332 42476 4284 42532
rect 4340 42476 4350 42532
rect 6178 42476 6188 42532
rect 6244 42476 8092 42532
rect 8148 42476 8158 42532
rect 20850 42476 20860 42532
rect 20916 42476 21980 42532
rect 22036 42476 22046 42532
rect 27458 42476 27468 42532
rect 27524 42476 27916 42532
rect 27972 42476 28476 42532
rect 28532 42476 28542 42532
rect 30706 42476 30716 42532
rect 30772 42476 31052 42532
rect 31108 42476 31118 42532
rect 31938 42476 31948 42532
rect 32004 42476 32014 42532
rect 45042 42476 45052 42532
rect 45108 42476 46508 42532
rect 46564 42476 46574 42532
rect 31948 42420 32004 42476
rect 3378 42364 3388 42420
rect 3444 42364 3482 42420
rect 5730 42364 5740 42420
rect 5796 42364 6300 42420
rect 6356 42364 8652 42420
rect 8708 42364 8718 42420
rect 20514 42364 20524 42420
rect 20580 42364 27244 42420
rect 27300 42364 27310 42420
rect 27580 42364 32004 42420
rect 57026 42364 57036 42420
rect 57092 42364 59500 42420
rect 59556 42364 61292 42420
rect 61348 42364 61964 42420
rect 62020 42364 62030 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 27580 42308 27636 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 3154 42252 3164 42308
rect 3220 42252 4172 42308
rect 4228 42252 4284 42308
rect 4340 42252 4350 42308
rect 7410 42252 7420 42308
rect 7476 42252 8316 42308
rect 8372 42252 8382 42308
rect 24546 42252 24556 42308
rect 24612 42252 27132 42308
rect 27188 42252 27636 42308
rect 27794 42252 27804 42308
rect 27860 42252 48860 42308
rect 48916 42252 48926 42308
rect 58034 42252 58044 42308
rect 58100 42252 59724 42308
rect 59780 42252 59790 42308
rect 6822 42140 6860 42196
rect 6916 42140 6926 42196
rect 7298 42140 7308 42196
rect 7364 42140 7374 42196
rect 16258 42140 16268 42196
rect 16324 42140 17948 42196
rect 18004 42140 18014 42196
rect 18386 42140 18396 42196
rect 18452 42140 21756 42196
rect 21812 42140 21822 42196
rect 24098 42140 24108 42196
rect 24164 42140 26124 42196
rect 26180 42140 26190 42196
rect 27010 42140 27020 42196
rect 27076 42140 32172 42196
rect 32228 42140 32238 42196
rect 41906 42140 41916 42196
rect 41972 42140 42924 42196
rect 42980 42140 42990 42196
rect 43670 42140 43708 42196
rect 43764 42140 43774 42196
rect 44370 42140 44380 42196
rect 44436 42140 47068 42196
rect 47124 42140 47134 42196
rect 48402 42140 48412 42196
rect 48468 42140 51548 42196
rect 51604 42140 51614 42196
rect 53414 42140 53452 42196
rect 53508 42140 53518 42196
rect 54226 42140 54236 42196
rect 54292 42140 57820 42196
rect 57876 42140 57886 42196
rect 59154 42140 59164 42196
rect 59220 42140 62412 42196
rect 62468 42140 62478 42196
rect 7308 42084 7364 42140
rect 43708 42084 43764 42140
rect 3938 42028 3948 42084
rect 4004 42028 6636 42084
rect 6692 42028 6702 42084
rect 6962 42028 6972 42084
rect 7028 42028 7364 42084
rect 7522 42028 7532 42084
rect 7588 42028 8092 42084
rect 8148 42028 8158 42084
rect 12674 42028 12684 42084
rect 12740 42028 14588 42084
rect 14644 42028 14654 42084
rect 15026 42028 15036 42084
rect 15092 42028 15148 42084
rect 15204 42028 15214 42084
rect 18162 42028 18172 42084
rect 18228 42028 21420 42084
rect 21476 42028 21486 42084
rect 27234 42028 27244 42084
rect 27300 42028 27916 42084
rect 27972 42028 27982 42084
rect 40898 42028 40908 42084
rect 40964 42028 41468 42084
rect 41524 42028 41534 42084
rect 42018 42028 42028 42084
rect 42084 42028 43764 42084
rect 44930 42028 44940 42084
rect 44996 42028 45724 42084
rect 45780 42028 45790 42084
rect 46050 42028 46060 42084
rect 46116 42028 46844 42084
rect 46900 42028 46910 42084
rect 49410 42028 49420 42084
rect 49476 42028 50316 42084
rect 50372 42028 51996 42084
rect 52052 42028 52062 42084
rect 52322 42028 52332 42084
rect 52388 42028 59612 42084
rect 59668 42028 59678 42084
rect 2034 41916 2044 41972
rect 2100 41916 2940 41972
rect 2996 41916 3006 41972
rect 3154 41916 3164 41972
rect 3220 41916 3836 41972
rect 3892 41916 3902 41972
rect 5058 41916 5068 41972
rect 5124 41916 6300 41972
rect 6356 41916 8652 41972
rect 8708 41916 8718 41972
rect 12002 41916 12012 41972
rect 12068 41916 13916 41972
rect 13972 41916 13982 41972
rect 15138 41916 15148 41972
rect 15204 41916 17500 41972
rect 17556 41916 17566 41972
rect 19282 41916 19292 41972
rect 19348 41916 20300 41972
rect 20356 41916 20748 41972
rect 20804 41916 20814 41972
rect 22418 41916 22428 41972
rect 22484 41916 23436 41972
rect 23492 41916 23502 41972
rect 24882 41916 24892 41972
rect 24948 41916 26012 41972
rect 26068 41916 26078 41972
rect 32386 41916 32396 41972
rect 32452 41916 32462 41972
rect 35522 41916 35532 41972
rect 35588 41916 36764 41972
rect 36820 41916 36830 41972
rect 37762 41916 37772 41972
rect 37828 41916 38444 41972
rect 38500 41916 38510 41972
rect 41346 41916 41356 41972
rect 41412 41916 42700 41972
rect 42756 41916 43260 41972
rect 43316 41916 43326 41972
rect 47842 41916 47852 41972
rect 47908 41916 50092 41972
rect 50148 41916 50158 41972
rect 52658 41916 52668 41972
rect 52724 41916 56700 41972
rect 56756 41916 56766 41972
rect 57026 41916 57036 41972
rect 57092 41916 58828 41972
rect 58884 41916 58894 41972
rect 61170 41916 61180 41972
rect 61236 41916 62076 41972
rect 62132 41916 62142 41972
rect 32396 41860 32452 41916
rect 2146 41804 2156 41860
rect 2212 41804 5516 41860
rect 5572 41804 5582 41860
rect 7186 41804 7196 41860
rect 7252 41804 8876 41860
rect 8932 41804 8942 41860
rect 9762 41804 9772 41860
rect 9828 41804 10780 41860
rect 10836 41804 10846 41860
rect 13234 41804 13244 41860
rect 13300 41804 14140 41860
rect 14196 41804 14206 41860
rect 16034 41804 16044 41860
rect 16100 41804 17164 41860
rect 17220 41804 17948 41860
rect 18004 41804 19404 41860
rect 19460 41804 20524 41860
rect 20580 41804 20590 41860
rect 21634 41804 21644 41860
rect 21700 41804 21868 41860
rect 21924 41804 22540 41860
rect 22596 41804 22606 41860
rect 30146 41804 30156 41860
rect 30212 41804 31836 41860
rect 31892 41804 31902 41860
rect 32396 41804 34748 41860
rect 34804 41804 35644 41860
rect 35700 41804 35710 41860
rect 47618 41804 47628 41860
rect 47684 41804 48972 41860
rect 49028 41804 49038 41860
rect 50530 41804 50540 41860
rect 50596 41804 51660 41860
rect 51716 41804 51996 41860
rect 52052 41804 52062 41860
rect 55346 41804 55356 41860
rect 55412 41804 56252 41860
rect 56308 41804 56318 41860
rect 57036 41748 57092 41916
rect 57362 41804 57372 41860
rect 57428 41804 57438 41860
rect 59490 41804 59500 41860
rect 59556 41804 61068 41860
rect 61124 41804 61134 41860
rect 61618 41804 61628 41860
rect 61684 41804 61852 41860
rect 61908 41804 61918 41860
rect 6962 41692 6972 41748
rect 7028 41692 10108 41748
rect 10164 41692 10174 41748
rect 11218 41692 11228 41748
rect 11284 41692 11900 41748
rect 11956 41692 11966 41748
rect 16930 41692 16940 41748
rect 16996 41692 19740 41748
rect 19796 41692 19806 41748
rect 22082 41692 22092 41748
rect 22148 41692 24220 41748
rect 24276 41692 24286 41748
rect 27346 41692 27356 41748
rect 27412 41692 27422 41748
rect 28130 41692 28140 41748
rect 28196 41692 33740 41748
rect 33796 41692 35084 41748
rect 35140 41692 35150 41748
rect 45266 41692 45276 41748
rect 45332 41692 46508 41748
rect 46564 41692 46574 41748
rect 53218 41692 53228 41748
rect 53284 41692 57092 41748
rect 57372 41748 57428 41804
rect 57372 41692 62300 41748
rect 62356 41692 62366 41748
rect 27356 41636 27412 41692
rect 7858 41580 7868 41636
rect 7924 41580 8764 41636
rect 8820 41580 8830 41636
rect 24434 41580 24444 41636
rect 24500 41580 25340 41636
rect 25396 41580 25406 41636
rect 27356 41580 32732 41636
rect 32788 41580 32798 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 2930 41468 2940 41524
rect 2996 41468 3388 41524
rect 23874 41468 23884 41524
rect 23940 41468 26348 41524
rect 26404 41468 26414 41524
rect 32134 41468 32172 41524
rect 32228 41468 32238 41524
rect 51202 41468 51212 41524
rect 51268 41468 61180 41524
rect 61236 41468 61246 41524
rect 3332 41412 3388 41468
rect 3332 41356 7420 41412
rect 7476 41356 9884 41412
rect 9940 41356 9950 41412
rect 15250 41356 15260 41412
rect 15316 41356 22652 41412
rect 22708 41356 22718 41412
rect 23090 41356 23100 41412
rect 23156 41356 25676 41412
rect 25732 41356 26572 41412
rect 26628 41356 26638 41412
rect 33506 41356 33516 41412
rect 33572 41356 35532 41412
rect 35588 41356 35598 41412
rect 36978 41356 36988 41412
rect 37044 41356 38108 41412
rect 38164 41356 38174 41412
rect 44146 41356 44156 41412
rect 44212 41356 52948 41412
rect 55766 41356 55804 41412
rect 55860 41356 55870 41412
rect 56466 41356 56476 41412
rect 56532 41356 56812 41412
rect 56868 41356 56878 41412
rect 60946 41356 60956 41412
rect 61012 41356 61628 41412
rect 61684 41356 61694 41412
rect 2930 41244 2940 41300
rect 2996 41244 3948 41300
rect 4004 41244 4014 41300
rect 6850 41244 6860 41300
rect 6916 41244 7644 41300
rect 7700 41244 7710 41300
rect 12562 41244 12572 41300
rect 12628 41244 12908 41300
rect 12964 41244 14476 41300
rect 14532 41244 14542 41300
rect 15362 41244 15372 41300
rect 15428 41244 15708 41300
rect 15764 41244 15774 41300
rect 34076 41244 37772 41300
rect 37828 41244 37838 41300
rect 7074 41132 7084 41188
rect 7140 41132 7532 41188
rect 7588 41132 7598 41188
rect 8306 41132 8316 41188
rect 8372 41132 11788 41188
rect 11844 41132 11854 41188
rect 12114 41132 12124 41188
rect 12180 41132 14420 41188
rect 16930 41132 16940 41188
rect 16996 41132 17612 41188
rect 17668 41132 17678 41188
rect 22530 41132 22540 41188
rect 22596 41132 24332 41188
rect 24388 41132 24398 41188
rect 28130 41132 28140 41188
rect 28196 41132 28476 41188
rect 28532 41132 29820 41188
rect 29876 41132 29886 41188
rect 8082 41020 8092 41076
rect 8148 41020 9548 41076
rect 9604 41020 9614 41076
rect 11330 41020 11340 41076
rect 11396 41020 12460 41076
rect 12516 41020 14140 41076
rect 14196 41020 14206 41076
rect 1922 40908 1932 40964
rect 1988 40908 6076 40964
rect 6132 40908 6142 40964
rect 7634 40908 7644 40964
rect 7700 40908 9772 40964
rect 9828 40908 9838 40964
rect 12674 40908 12684 40964
rect 12740 40908 13244 40964
rect 13300 40908 13580 40964
rect 13636 40908 13646 40964
rect 14364 40852 14420 41132
rect 15026 41020 15036 41076
rect 15092 41020 20636 41076
rect 20692 41020 20702 41076
rect 21746 41020 21756 41076
rect 21812 41020 22988 41076
rect 23044 41020 23054 41076
rect 25666 41020 25676 41076
rect 25732 41020 33404 41076
rect 33460 41020 33470 41076
rect 34076 40964 34132 41244
rect 52892 41188 52948 41356
rect 55346 41244 55356 41300
rect 55412 41244 55916 41300
rect 55972 41244 61740 41300
rect 61796 41244 61806 41300
rect 34290 41132 34300 41188
rect 34356 41132 34860 41188
rect 34916 41132 37884 41188
rect 37940 41132 37950 41188
rect 47730 41132 47740 41188
rect 47796 41132 52332 41188
rect 52388 41132 52398 41188
rect 52854 41132 52892 41188
rect 52948 41132 52958 41188
rect 54562 41132 54572 41188
rect 54628 41132 60508 41188
rect 60564 41132 60574 41188
rect 35074 41020 35084 41076
rect 35140 41020 37212 41076
rect 37268 41020 37278 41076
rect 40562 41020 40572 41076
rect 40628 41020 41468 41076
rect 41524 41020 41534 41076
rect 48962 41020 48972 41076
rect 49028 41020 49868 41076
rect 49924 41020 49934 41076
rect 55906 41020 55916 41076
rect 55972 41020 57036 41076
rect 57092 41020 57102 41076
rect 59714 41020 59724 41076
rect 59780 41020 61404 41076
rect 61460 41020 61470 41076
rect 15474 40908 15484 40964
rect 15540 40908 16044 40964
rect 16100 40908 16110 40964
rect 16258 40908 16268 40964
rect 16324 40908 16604 40964
rect 16660 40908 16670 40964
rect 18386 40908 18396 40964
rect 18452 40908 18844 40964
rect 18900 40908 19068 40964
rect 19124 40908 19134 40964
rect 19628 40908 20468 40964
rect 21634 40908 21644 40964
rect 21700 40908 23996 40964
rect 24052 40908 24062 40964
rect 29026 40908 29036 40964
rect 29092 40908 30828 40964
rect 30884 40908 34132 40964
rect 34486 40908 34524 40964
rect 34580 40908 34590 40964
rect 35858 40908 35868 40964
rect 35924 40908 36988 40964
rect 37044 40908 37054 40964
rect 37426 40908 37436 40964
rect 37492 40908 38444 40964
rect 38500 40908 38510 40964
rect 39666 40908 39676 40964
rect 39732 40908 40908 40964
rect 40964 40908 40974 40964
rect 46050 40908 46060 40964
rect 46116 40908 47292 40964
rect 47348 40908 47358 40964
rect 50372 40908 50764 40964
rect 50820 40908 50830 40964
rect 53106 40908 53116 40964
rect 53172 40908 55468 40964
rect 55524 40908 55534 40964
rect 56578 40908 56588 40964
rect 56644 40908 60956 40964
rect 61012 40908 61964 40964
rect 62020 40908 62030 40964
rect 19628 40852 19684 40908
rect 14364 40796 19684 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 20412 40740 20468 40908
rect 20626 40796 20636 40852
rect 20692 40796 22652 40852
rect 22708 40796 24108 40852
rect 24164 40796 24668 40852
rect 24724 40796 24734 40852
rect 28578 40796 28588 40852
rect 28644 40796 30044 40852
rect 30100 40796 31164 40852
rect 31220 40796 31230 40852
rect 32722 40796 32732 40852
rect 32788 40796 34972 40852
rect 35028 40796 36876 40852
rect 36932 40796 36942 40852
rect 39778 40796 39788 40852
rect 39844 40796 40796 40852
rect 40852 40796 40862 40852
rect 42466 40796 42476 40852
rect 42532 40796 47852 40852
rect 47908 40796 47918 40852
rect 50372 40740 50428 40908
rect 55122 40796 55132 40852
rect 55188 40796 59052 40852
rect 59108 40796 59612 40852
rect 59668 40796 59678 40852
rect 61058 40796 61068 40852
rect 61124 40796 62524 40852
rect 62580 40796 62590 40852
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 2258 40684 2268 40740
rect 2324 40684 7196 40740
rect 7252 40684 7262 40740
rect 20412 40684 24220 40740
rect 24276 40684 24612 40740
rect 24770 40684 24780 40740
rect 24836 40684 26012 40740
rect 26068 40684 26078 40740
rect 28690 40684 28700 40740
rect 28756 40684 29372 40740
rect 29428 40684 31500 40740
rect 31556 40684 31566 40740
rect 35746 40684 35756 40740
rect 35812 40684 46116 40740
rect 47058 40684 47068 40740
rect 47124 40684 47404 40740
rect 47460 40684 50428 40740
rect 54562 40684 54572 40740
rect 54628 40684 55692 40740
rect 55748 40684 61740 40740
rect 61796 40684 61806 40740
rect 24556 40628 24612 40684
rect 6178 40572 6188 40628
rect 6244 40572 7756 40628
rect 7812 40572 7822 40628
rect 10322 40572 10332 40628
rect 10388 40572 12012 40628
rect 12068 40572 12078 40628
rect 14914 40572 14924 40628
rect 14980 40572 22204 40628
rect 22260 40572 23660 40628
rect 23716 40572 23726 40628
rect 24556 40572 24668 40628
rect 24724 40572 25228 40628
rect 25284 40572 25294 40628
rect 27010 40572 27020 40628
rect 27076 40572 29484 40628
rect 29540 40572 29550 40628
rect 40450 40572 40460 40628
rect 40516 40572 41244 40628
rect 41300 40572 41310 40628
rect 43026 40572 43036 40628
rect 43092 40572 43932 40628
rect 43988 40572 43998 40628
rect 44258 40572 44268 40628
rect 44324 40572 45164 40628
rect 45220 40572 45724 40628
rect 45780 40572 45790 40628
rect 2706 40460 2716 40516
rect 2772 40460 3164 40516
rect 3220 40460 3836 40516
rect 3892 40460 3902 40516
rect 7522 40460 7532 40516
rect 7588 40460 8092 40516
rect 8148 40460 8158 40516
rect 16828 40460 17948 40516
rect 18004 40460 22092 40516
rect 22148 40460 22158 40516
rect 25666 40460 25676 40516
rect 25732 40460 27580 40516
rect 27636 40460 27646 40516
rect 36082 40460 36092 40516
rect 36148 40460 37212 40516
rect 37268 40460 37278 40516
rect 38322 40460 38332 40516
rect 38388 40460 40908 40516
rect 40964 40460 42028 40516
rect 42084 40460 45276 40516
rect 45332 40460 45342 40516
rect 9874 40348 9884 40404
rect 9940 40348 11340 40404
rect 11396 40348 11406 40404
rect 14550 40348 14588 40404
rect 14644 40348 14654 40404
rect 2370 40236 2380 40292
rect 2436 40236 3388 40292
rect 3444 40236 3454 40292
rect 7074 40236 7084 40292
rect 7140 40236 8876 40292
rect 8932 40236 8942 40292
rect 13122 40236 13132 40292
rect 13188 40236 15484 40292
rect 15540 40236 15550 40292
rect 16828 40180 16884 40460
rect 46060 40404 46116 40684
rect 56914 40572 56924 40628
rect 56980 40572 58268 40628
rect 58324 40572 58334 40628
rect 61170 40572 61180 40628
rect 61236 40572 62300 40628
rect 62356 40572 62366 40628
rect 47170 40460 47180 40516
rect 47236 40460 49980 40516
rect 50036 40460 53228 40516
rect 53284 40460 53294 40516
rect 54198 40460 54236 40516
rect 54292 40460 54302 40516
rect 55794 40460 55804 40516
rect 55860 40460 56700 40516
rect 56756 40460 56766 40516
rect 57026 40460 57036 40516
rect 57092 40460 60620 40516
rect 60676 40460 60686 40516
rect 61394 40460 61404 40516
rect 61460 40460 61740 40516
rect 61796 40460 61806 40516
rect 18162 40348 18172 40404
rect 18228 40348 20412 40404
rect 20468 40348 21420 40404
rect 21476 40348 21486 40404
rect 29026 40348 29036 40404
rect 29092 40348 30492 40404
rect 30548 40348 30558 40404
rect 34178 40348 34188 40404
rect 34244 40348 34860 40404
rect 34916 40348 34926 40404
rect 36866 40348 36876 40404
rect 36932 40348 37436 40404
rect 37492 40348 37502 40404
rect 46050 40348 46060 40404
rect 46116 40348 46126 40404
rect 49746 40348 49756 40404
rect 49812 40348 50428 40404
rect 50484 40348 50494 40404
rect 54674 40348 54684 40404
rect 54740 40348 56364 40404
rect 56420 40348 57820 40404
rect 57876 40348 57886 40404
rect 61058 40348 61068 40404
rect 61124 40348 61134 40404
rect 61506 40348 61516 40404
rect 61572 40348 62076 40404
rect 62132 40348 62142 40404
rect 61068 40292 61124 40348
rect 19058 40236 19068 40292
rect 19124 40236 20188 40292
rect 20244 40236 20254 40292
rect 27346 40236 27356 40292
rect 27412 40236 27916 40292
rect 27972 40236 27982 40292
rect 30034 40236 30044 40292
rect 30100 40236 31276 40292
rect 31332 40236 31724 40292
rect 31780 40236 31790 40292
rect 33506 40236 33516 40292
rect 33572 40236 34636 40292
rect 34692 40236 35420 40292
rect 35476 40236 35486 40292
rect 40338 40236 40348 40292
rect 40404 40236 42924 40292
rect 42980 40236 42990 40292
rect 45490 40236 45500 40292
rect 45556 40236 48636 40292
rect 48692 40236 48702 40292
rect 48850 40236 48860 40292
rect 48916 40236 53788 40292
rect 53844 40236 53854 40292
rect 56018 40236 56028 40292
rect 56084 40236 57260 40292
rect 57316 40236 60228 40292
rect 60386 40236 60396 40292
rect 60452 40236 61124 40292
rect 60172 40180 60228 40236
rect 13346 40124 13356 40180
rect 13412 40124 14252 40180
rect 14308 40124 14700 40180
rect 14756 40124 14766 40180
rect 16818 40124 16828 40180
rect 16884 40124 16894 40180
rect 18050 40124 18060 40180
rect 18116 40124 23884 40180
rect 23940 40124 23950 40180
rect 26852 40124 38668 40180
rect 49634 40124 49644 40180
rect 49700 40124 54348 40180
rect 54404 40124 54414 40180
rect 55122 40124 55132 40180
rect 55188 40124 57932 40180
rect 57988 40124 57998 40180
rect 60172 40124 60508 40180
rect 60564 40124 60574 40180
rect 61926 40124 61964 40180
rect 62020 40124 62030 40180
rect 22418 40012 22428 40068
rect 22484 40012 23212 40068
rect 23268 40012 26124 40068
rect 26180 40012 26190 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 26852 39956 26908 40124
rect 38612 40068 38668 40124
rect 62132 40068 62188 40292
rect 62244 40236 62254 40292
rect 29138 40012 29148 40068
rect 29204 40012 31164 40068
rect 31220 40012 31230 40068
rect 38612 40012 39564 40068
rect 39620 40012 39630 40068
rect 44258 40012 44268 40068
rect 44324 40012 44940 40068
rect 44996 40012 46844 40068
rect 46900 40012 49084 40068
rect 49140 40012 49150 40068
rect 53218 40012 53228 40068
rect 53284 40012 62188 40068
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 6066 39900 6076 39956
rect 6132 39900 13692 39956
rect 13748 39900 13758 39956
rect 16482 39900 16492 39956
rect 16548 39900 26908 39956
rect 28242 39900 28252 39956
rect 28308 39900 28588 39956
rect 28644 39900 28654 39956
rect 28914 39900 28924 39956
rect 28980 39900 31052 39956
rect 31108 39900 31118 39956
rect 54786 39900 54796 39956
rect 54852 39900 55580 39956
rect 55636 39900 55646 39956
rect 55906 39900 55916 39956
rect 55972 39900 62076 39956
rect 62132 39900 62142 39956
rect 7858 39788 7868 39844
rect 7924 39788 9772 39844
rect 9828 39788 9838 39844
rect 14018 39788 14028 39844
rect 14084 39788 16828 39844
rect 16884 39788 16894 39844
rect 28466 39788 28476 39844
rect 28532 39788 29820 39844
rect 29876 39788 29886 39844
rect 32610 39788 32620 39844
rect 32676 39788 34524 39844
rect 34580 39788 36428 39844
rect 36484 39788 36494 39844
rect 38658 39788 38668 39844
rect 38724 39788 39228 39844
rect 39284 39788 40012 39844
rect 40068 39788 40078 39844
rect 54002 39788 54012 39844
rect 54068 39788 56364 39844
rect 56420 39788 56430 39844
rect 58258 39788 58268 39844
rect 58324 39788 60956 39844
rect 61012 39788 61022 39844
rect 4162 39676 4172 39732
rect 4228 39676 5628 39732
rect 5684 39676 5694 39732
rect 6066 39676 6076 39732
rect 6132 39676 6972 39732
rect 7028 39676 7038 39732
rect 7298 39676 7308 39732
rect 7364 39676 8540 39732
rect 8596 39676 8606 39732
rect 11778 39676 11788 39732
rect 11844 39676 34020 39732
rect 43922 39676 43932 39732
rect 43988 39676 47404 39732
rect 47460 39676 47470 39732
rect 50306 39676 50316 39732
rect 50372 39676 53564 39732
rect 53620 39676 53630 39732
rect 57250 39676 57260 39732
rect 57316 39676 59500 39732
rect 59556 39676 59566 39732
rect 6402 39564 6412 39620
rect 6468 39564 6860 39620
rect 6916 39564 7868 39620
rect 7924 39564 7934 39620
rect 9986 39564 9996 39620
rect 10052 39564 11004 39620
rect 11060 39564 11070 39620
rect 11442 39564 11452 39620
rect 11508 39564 13804 39620
rect 13860 39564 14028 39620
rect 14084 39564 14094 39620
rect 14466 39564 14476 39620
rect 14532 39564 15036 39620
rect 15092 39564 15102 39620
rect 15250 39564 15260 39620
rect 15316 39564 15820 39620
rect 15876 39564 16660 39620
rect 16930 39564 16940 39620
rect 16996 39564 18396 39620
rect 18452 39564 18462 39620
rect 27458 39564 27468 39620
rect 27524 39564 29596 39620
rect 29652 39564 29662 39620
rect 16604 39508 16660 39564
rect 33964 39508 34020 39676
rect 47954 39564 47964 39620
rect 48020 39564 48748 39620
rect 48804 39564 48814 39620
rect 50418 39564 50428 39620
rect 50484 39564 51436 39620
rect 51492 39564 51502 39620
rect 55346 39564 55356 39620
rect 55412 39564 59836 39620
rect 59892 39564 59902 39620
rect 1474 39452 1484 39508
rect 1540 39452 2268 39508
rect 2324 39452 2334 39508
rect 6290 39452 6300 39508
rect 6356 39452 8540 39508
rect 8596 39452 8606 39508
rect 14802 39452 14812 39508
rect 14868 39452 15932 39508
rect 15988 39452 15998 39508
rect 16594 39452 16604 39508
rect 16660 39452 17612 39508
rect 17668 39452 17678 39508
rect 17938 39452 17948 39508
rect 18004 39452 21308 39508
rect 21364 39452 21374 39508
rect 22306 39452 22316 39508
rect 22372 39452 25228 39508
rect 25284 39452 26460 39508
rect 26516 39452 26526 39508
rect 27346 39452 27356 39508
rect 27412 39452 28252 39508
rect 28308 39452 29148 39508
rect 29204 39452 29214 39508
rect 33954 39452 33964 39508
rect 34020 39452 34030 39508
rect 36428 39452 38220 39508
rect 38276 39452 38286 39508
rect 41122 39452 41132 39508
rect 41188 39452 42700 39508
rect 42756 39452 42766 39508
rect 47282 39452 47292 39508
rect 47348 39452 49980 39508
rect 50036 39452 50046 39508
rect 50306 39452 50316 39508
rect 50372 39452 51212 39508
rect 51268 39452 51278 39508
rect 55570 39452 55580 39508
rect 55636 39452 57148 39508
rect 57204 39452 57214 39508
rect 36428 39396 36484 39452
rect 3714 39340 3724 39396
rect 3780 39340 4396 39396
rect 4452 39340 4462 39396
rect 4722 39340 4732 39396
rect 4788 39340 5292 39396
rect 5348 39340 5358 39396
rect 14690 39340 14700 39396
rect 14756 39340 18508 39396
rect 18564 39340 18574 39396
rect 31602 39340 31612 39396
rect 31668 39340 36484 39396
rect 36642 39340 36652 39396
rect 36708 39340 40460 39396
rect 40516 39340 40526 39396
rect 47394 39340 47404 39396
rect 47460 39340 51772 39396
rect 51828 39340 51838 39396
rect 57250 39340 57260 39396
rect 57316 39340 58156 39396
rect 58212 39340 61292 39396
rect 61348 39340 61358 39396
rect 17574 39228 17612 39284
rect 17668 39228 17678 39284
rect 19366 39228 19404 39284
rect 19460 39228 19470 39284
rect 26114 39228 26124 39284
rect 26180 39228 26796 39284
rect 26852 39228 26862 39284
rect 42802 39228 42812 39284
rect 42868 39228 47516 39284
rect 47572 39228 50428 39284
rect 52098 39228 52108 39284
rect 52164 39228 61404 39284
rect 61460 39228 61470 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 1586 39116 1596 39172
rect 1652 39116 8652 39172
rect 8708 39116 8718 39172
rect 16482 39116 16492 39172
rect 16548 39116 17276 39172
rect 17332 39116 17948 39172
rect 18004 39116 18014 39172
rect 42018 39116 42028 39172
rect 42084 39116 43036 39172
rect 43092 39116 43102 39172
rect 46508 39116 49196 39172
rect 49252 39116 49262 39172
rect 46508 39060 46564 39116
rect 3938 39004 3948 39060
rect 4004 39004 30716 39060
rect 30772 39004 30782 39060
rect 41122 39004 41132 39060
rect 41188 39004 41692 39060
rect 41748 39004 42140 39060
rect 42196 39004 42206 39060
rect 46498 39004 46508 39060
rect 46564 39004 46574 39060
rect 47954 39004 47964 39060
rect 48020 39004 50148 39060
rect 50372 39004 50428 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 50484 39004 50494 39060
rect 53106 39004 53116 39060
rect 53172 39004 53182 39060
rect 57810 39004 57820 39060
rect 57876 39004 58212 39060
rect 58482 39004 58492 39060
rect 58548 39004 59052 39060
rect 59108 39004 59724 39060
rect 59780 39004 59790 39060
rect 50092 38948 50148 39004
rect 53116 38948 53172 39004
rect 1138 38892 1148 38948
rect 1204 38892 1596 38948
rect 1652 38892 1662 38948
rect 4722 38892 4732 38948
rect 4788 38892 5068 38948
rect 5124 38892 5134 38948
rect 9762 38892 9772 38948
rect 9828 38892 12684 38948
rect 12740 38892 13356 38948
rect 13412 38892 15148 38948
rect 17154 38892 17164 38948
rect 17220 38892 17724 38948
rect 17780 38892 17790 38948
rect 20066 38892 20076 38948
rect 20132 38892 23548 38948
rect 23604 38892 23614 38948
rect 25554 38892 25564 38948
rect 25620 38892 25900 38948
rect 25956 38892 29484 38948
rect 29540 38892 30380 38948
rect 30436 38892 30446 38948
rect 31938 38892 31948 38948
rect 32004 38892 34188 38948
rect 34244 38892 34254 38948
rect 40338 38892 40348 38948
rect 40404 38892 41356 38948
rect 41412 38892 41422 38948
rect 46722 38892 46732 38948
rect 46788 38892 47628 38948
rect 47684 38892 48748 38948
rect 48804 38892 48814 38948
rect 50092 38892 50316 38948
rect 50372 38892 50382 38948
rect 51324 38892 53172 38948
rect 58156 38948 58212 39004
rect 58156 38892 59612 38948
rect 59668 38892 60508 38948
rect 60564 38892 60574 38948
rect 60946 38892 60956 38948
rect 61012 38892 61852 38948
rect 61908 38892 61918 38948
rect 15092 38836 15148 38892
rect 51324 38836 51380 38892
rect 4386 38780 4396 38836
rect 4452 38780 5404 38836
rect 5460 38780 5964 38836
rect 6020 38780 6030 38836
rect 10098 38780 10108 38836
rect 10164 38780 10556 38836
rect 10612 38780 10622 38836
rect 10770 38780 10780 38836
rect 10836 38780 11228 38836
rect 11284 38780 11788 38836
rect 11844 38780 14364 38836
rect 14420 38780 14430 38836
rect 15092 38780 16156 38836
rect 16212 38780 16222 38836
rect 19170 38780 19180 38836
rect 19236 38780 21196 38836
rect 21252 38780 21262 38836
rect 23986 38780 23996 38836
rect 24052 38780 25788 38836
rect 25844 38780 25854 38836
rect 26898 38780 26908 38836
rect 26964 38780 32508 38836
rect 32564 38780 33404 38836
rect 33460 38780 33470 38836
rect 41570 38780 41580 38836
rect 41636 38780 43484 38836
rect 43540 38780 43550 38836
rect 45042 38780 45052 38836
rect 45108 38780 45836 38836
rect 45892 38780 46956 38836
rect 47012 38780 47022 38836
rect 47730 38780 47740 38836
rect 47796 38780 49532 38836
rect 49588 38780 49868 38836
rect 49924 38780 51380 38836
rect 51538 38780 51548 38836
rect 51604 38780 52444 38836
rect 52500 38780 52510 38836
rect 52994 38780 53004 38836
rect 53060 38780 53788 38836
rect 53844 38780 53854 38836
rect 55906 38780 55916 38836
rect 55972 38780 60732 38836
rect 60788 38780 61404 38836
rect 61460 38780 61470 38836
rect 7298 38668 7308 38724
rect 7364 38668 9996 38724
rect 10052 38668 11004 38724
rect 11060 38668 11070 38724
rect 11666 38668 11676 38724
rect 11732 38668 13244 38724
rect 13300 38668 14700 38724
rect 14756 38668 14766 38724
rect 22194 38668 22204 38724
rect 22260 38668 22652 38724
rect 22708 38668 22718 38724
rect 25666 38668 25676 38724
rect 25732 38668 25742 38724
rect 31266 38668 31276 38724
rect 31332 38668 32060 38724
rect 32116 38668 32126 38724
rect 41234 38668 41244 38724
rect 41300 38668 42980 38724
rect 49410 38668 49420 38724
rect 49476 38668 50764 38724
rect 50820 38668 50830 38724
rect 53330 38668 53340 38724
rect 53396 38668 56700 38724
rect 56756 38668 56766 38724
rect 25676 38612 25732 38668
rect 42924 38612 42980 38668
rect 49420 38612 49476 38668
rect 2034 38556 2044 38612
rect 2100 38556 20412 38612
rect 20468 38556 20860 38612
rect 20916 38556 23324 38612
rect 23380 38556 23390 38612
rect 25676 38556 26124 38612
rect 26180 38556 26190 38612
rect 30594 38556 30604 38612
rect 30660 38556 32172 38612
rect 32228 38556 32238 38612
rect 37314 38556 37324 38612
rect 37380 38556 42140 38612
rect 42196 38556 42206 38612
rect 42914 38556 42924 38612
rect 42980 38556 42990 38612
rect 46722 38556 46732 38612
rect 46788 38556 47516 38612
rect 47572 38556 47582 38612
rect 48178 38556 48188 38612
rect 48244 38556 49476 38612
rect 51202 38556 51212 38612
rect 51268 38556 51548 38612
rect 51604 38556 52108 38612
rect 52164 38556 52174 38612
rect 54786 38556 54796 38612
rect 54852 38556 58044 38612
rect 58100 38556 59276 38612
rect 59332 38556 59342 38612
rect 51212 38500 51268 38556
rect 24210 38444 24220 38500
rect 24276 38444 25564 38500
rect 25620 38444 25630 38500
rect 28914 38444 28924 38500
rect 28980 38444 32956 38500
rect 33012 38444 34300 38500
rect 34356 38444 34366 38500
rect 41794 38444 41804 38500
rect 41860 38444 41870 38500
rect 42802 38444 42812 38500
rect 42868 38444 43596 38500
rect 43652 38444 43662 38500
rect 48402 38444 48412 38500
rect 48468 38444 51268 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 41804 38388 41860 38444
rect 19478 38332 19516 38388
rect 19572 38332 21532 38388
rect 21588 38332 22540 38388
rect 22596 38332 22606 38388
rect 25666 38332 25676 38388
rect 25732 38332 27692 38388
rect 27748 38332 27758 38388
rect 28130 38332 28140 38388
rect 28196 38332 29932 38388
rect 29988 38332 29998 38388
rect 41804 38332 42028 38388
rect 42084 38332 42094 38388
rect 46694 38332 46732 38388
rect 46788 38332 46798 38388
rect 2258 38220 2268 38276
rect 2324 38220 15260 38276
rect 15316 38220 15326 38276
rect 15586 38220 15596 38276
rect 15652 38220 16268 38276
rect 16324 38220 16334 38276
rect 28466 38220 28476 38276
rect 28532 38220 31500 38276
rect 31556 38220 32956 38276
rect 33012 38220 33022 38276
rect 41458 38220 41468 38276
rect 41524 38220 42700 38276
rect 42756 38220 43596 38276
rect 43652 38220 43662 38276
rect 48038 38220 48076 38276
rect 48132 38220 48142 38276
rect 55794 38220 55804 38276
rect 55860 38220 56812 38276
rect 56868 38220 56878 38276
rect 3042 38108 3052 38164
rect 3108 38108 4956 38164
rect 5012 38108 28924 38164
rect 28980 38108 28990 38164
rect 31154 38108 31164 38164
rect 31220 38108 32060 38164
rect 32116 38108 33404 38164
rect 33460 38108 33470 38164
rect 44930 38108 44940 38164
rect 44996 38108 46620 38164
rect 46676 38108 47964 38164
rect 48020 38108 48748 38164
rect 48804 38108 48814 38164
rect 58930 38108 58940 38164
rect 58996 38108 59500 38164
rect 59556 38108 59566 38164
rect 8642 37996 8652 38052
rect 8708 37996 9548 38052
rect 9604 37996 9614 38052
rect 13458 37996 13468 38052
rect 13524 37996 14588 38052
rect 14644 37996 15596 38052
rect 15652 37996 15932 38052
rect 15988 37996 15998 38052
rect 19842 37996 19852 38052
rect 19908 37996 20748 38052
rect 20804 37996 21084 38052
rect 21140 37996 21150 38052
rect 21494 37996 21532 38052
rect 21588 37996 21598 38052
rect 28242 37996 28252 38052
rect 28308 37996 29932 38052
rect 29988 37996 29998 38052
rect 30258 37996 30268 38052
rect 30324 37996 31948 38052
rect 32004 37996 32014 38052
rect 33282 37996 33292 38052
rect 33348 37996 34076 38052
rect 34132 37996 36092 38052
rect 36148 37996 36158 38052
rect 42130 37996 42140 38052
rect 42196 37996 42700 38052
rect 42756 37996 47180 38052
rect 47236 37996 47246 38052
rect 48066 37996 48076 38052
rect 48132 37996 49308 38052
rect 49364 37996 49374 38052
rect 50754 37996 50764 38052
rect 50820 37996 51996 38052
rect 52052 37996 52062 38052
rect 54898 37996 54908 38052
rect 54964 37996 55916 38052
rect 55972 37996 55982 38052
rect 58818 37996 58828 38052
rect 58884 37996 60508 38052
rect 60564 37996 60574 38052
rect 60946 37996 60956 38052
rect 61012 37996 61292 38052
rect 61348 37996 61358 38052
rect 29932 37940 29988 37996
rect 1586 37884 1596 37940
rect 1652 37884 2716 37940
rect 2772 37884 2782 37940
rect 9090 37884 9100 37940
rect 9156 37884 12684 37940
rect 12740 37884 13692 37940
rect 13748 37884 13758 37940
rect 15138 37884 15148 37940
rect 15204 37884 15708 37940
rect 15764 37884 15774 37940
rect 18498 37884 18508 37940
rect 18564 37884 19404 37940
rect 19460 37884 21420 37940
rect 21476 37884 21486 37940
rect 27234 37884 27244 37940
rect 27300 37884 29148 37940
rect 29204 37884 29214 37940
rect 29932 37884 31164 37940
rect 31220 37884 31230 37940
rect 33506 37884 33516 37940
rect 33572 37884 34636 37940
rect 34692 37884 34702 37940
rect 43698 37884 43708 37940
rect 43764 37884 44716 37940
rect 44772 37884 47292 37940
rect 47348 37884 47358 37940
rect 49522 37884 49532 37940
rect 49588 37884 49868 37940
rect 49924 37884 49934 37940
rect 52322 37884 52332 37940
rect 52388 37884 53900 37940
rect 53956 37884 53966 37940
rect 55010 37884 55020 37940
rect 55076 37884 56588 37940
rect 56644 37884 56654 37940
rect 57698 37884 57708 37940
rect 57764 37884 60844 37940
rect 60900 37884 60910 37940
rect 4834 37772 4844 37828
rect 4900 37772 6412 37828
rect 6468 37772 6478 37828
rect 9314 37772 9324 37828
rect 9380 37772 14700 37828
rect 14756 37772 14766 37828
rect 20374 37772 20412 37828
rect 20468 37772 20478 37828
rect 22754 37772 22764 37828
rect 22820 37772 25340 37828
rect 25396 37772 25406 37828
rect 26852 37772 28700 37828
rect 28756 37772 28766 37828
rect 35074 37772 35084 37828
rect 35140 37772 37100 37828
rect 37156 37772 40348 37828
rect 40404 37772 40414 37828
rect 43138 37772 43148 37828
rect 43204 37772 43820 37828
rect 43876 37772 43886 37828
rect 45714 37772 45724 37828
rect 45780 37772 45790 37828
rect 47842 37772 47852 37828
rect 47908 37772 48412 37828
rect 48468 37772 48478 37828
rect 50194 37772 50204 37828
rect 50260 37772 51100 37828
rect 51156 37772 51166 37828
rect 2706 37660 2716 37716
rect 2772 37660 3388 37716
rect 3444 37660 3948 37716
rect 4004 37660 4014 37716
rect 4844 37492 4900 37772
rect 7858 37660 7868 37716
rect 7924 37660 8316 37716
rect 8372 37660 10220 37716
rect 10276 37660 10286 37716
rect 11106 37660 11116 37716
rect 11172 37660 11452 37716
rect 11508 37660 11518 37716
rect 15708 37660 19572 37716
rect 15708 37604 15764 37660
rect 5058 37548 5068 37604
rect 5124 37548 11788 37604
rect 13346 37548 13356 37604
rect 13412 37548 13916 37604
rect 13972 37548 13982 37604
rect 15148 37548 15764 37604
rect 11732 37492 11788 37548
rect 15148 37492 15204 37548
rect 19516 37492 19572 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 25340 37604 25396 37772
rect 26786 37660 26796 37716
rect 26852 37660 26908 37772
rect 45724 37716 45780 37772
rect 27682 37660 27692 37716
rect 27748 37660 29148 37716
rect 29204 37660 29214 37716
rect 34066 37660 34076 37716
rect 34132 37660 34524 37716
rect 34580 37660 34590 37716
rect 39442 37660 39452 37716
rect 39508 37660 45780 37716
rect 47506 37660 47516 37716
rect 47572 37660 48972 37716
rect 49028 37660 49868 37716
rect 49924 37660 49934 37716
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 25340 37548 27132 37604
rect 27188 37548 27198 37604
rect 2482 37436 2492 37492
rect 2548 37436 3276 37492
rect 3332 37436 4900 37492
rect 6066 37436 6076 37492
rect 6132 37436 8652 37492
rect 8708 37436 8718 37492
rect 11732 37436 15204 37492
rect 16044 37436 17556 37492
rect 19516 37436 26908 37492
rect 26964 37436 26974 37492
rect 32498 37436 32508 37492
rect 32564 37436 33628 37492
rect 33684 37436 33694 37492
rect 34514 37436 34524 37492
rect 34580 37436 36988 37492
rect 37044 37436 37054 37492
rect 39778 37436 39788 37492
rect 39844 37436 41468 37492
rect 41524 37436 44268 37492
rect 44324 37436 44334 37492
rect 46834 37436 46844 37492
rect 46900 37436 48860 37492
rect 48916 37436 48926 37492
rect 49186 37436 49196 37492
rect 49252 37436 54012 37492
rect 54068 37436 54078 37492
rect 59490 37436 59500 37492
rect 59556 37436 60396 37492
rect 60452 37436 61068 37492
rect 61124 37436 61628 37492
rect 61684 37436 61694 37492
rect 16044 37380 16100 37436
rect 2818 37324 2828 37380
rect 2884 37324 4060 37380
rect 4116 37324 4732 37380
rect 4788 37324 4798 37380
rect 7970 37324 7980 37380
rect 8036 37324 8988 37380
rect 9044 37324 9054 37380
rect 13346 37324 13356 37380
rect 13412 37324 16100 37380
rect 17500 37268 17556 37436
rect 36530 37324 36540 37380
rect 36596 37324 39676 37380
rect 39732 37324 39742 37380
rect 45826 37324 45836 37380
rect 45892 37324 49420 37380
rect 49476 37324 50316 37380
rect 50372 37324 51884 37380
rect 51940 37324 51950 37380
rect 56690 37324 56700 37380
rect 56756 37324 60620 37380
rect 60676 37324 60686 37380
rect 12450 37212 12460 37268
rect 12516 37212 13916 37268
rect 13972 37212 13982 37268
rect 14354 37212 14364 37268
rect 14420 37212 16044 37268
rect 16100 37212 16110 37268
rect 17490 37212 17500 37268
rect 17556 37212 17948 37268
rect 18004 37212 23548 37268
rect 23604 37212 23614 37268
rect 26226 37212 26236 37268
rect 26292 37212 28588 37268
rect 28644 37212 28654 37268
rect 29026 37212 29036 37268
rect 29092 37212 31500 37268
rect 31556 37212 31566 37268
rect 33394 37212 33404 37268
rect 33460 37212 34188 37268
rect 34244 37212 35308 37268
rect 36306 37212 36316 37268
rect 36372 37212 36876 37268
rect 36932 37212 36942 37268
rect 37874 37212 37884 37268
rect 37940 37212 41020 37268
rect 41076 37212 41086 37268
rect 44930 37212 44940 37268
rect 44996 37212 46172 37268
rect 46228 37212 46238 37268
rect 46386 37212 46396 37268
rect 46452 37212 51100 37268
rect 51156 37212 52556 37268
rect 52612 37212 52622 37268
rect 54226 37212 54236 37268
rect 54292 37212 56924 37268
rect 56980 37212 56990 37268
rect 62038 37212 62076 37268
rect 62132 37212 62142 37268
rect 35252 37156 35308 37212
rect 5730 37100 5740 37156
rect 5796 37100 22652 37156
rect 22708 37100 24668 37156
rect 24724 37100 27804 37156
rect 27860 37100 27870 37156
rect 32162 37100 32172 37156
rect 32228 37100 33852 37156
rect 33908 37100 33918 37156
rect 35252 37100 38780 37156
rect 38836 37100 38846 37156
rect 40338 37100 40348 37156
rect 40404 37100 41132 37156
rect 41188 37100 41692 37156
rect 41748 37100 41758 37156
rect 54114 37100 54124 37156
rect 54180 37100 59500 37156
rect 59556 37100 59566 37156
rect 3602 36988 3612 37044
rect 3668 36988 6636 37044
rect 6692 36988 6702 37044
rect 9874 36988 9884 37044
rect 9940 36988 11340 37044
rect 11396 36988 12236 37044
rect 12292 36988 12302 37044
rect 14018 36988 14028 37044
rect 14084 36988 15148 37044
rect 15204 36988 15214 37044
rect 20178 36988 20188 37044
rect 20244 36988 26684 37044
rect 26740 36988 26750 37044
rect 27682 36988 27692 37044
rect 27748 36988 30604 37044
rect 30660 36988 33628 37044
rect 33684 36988 33694 37044
rect 34402 36988 34412 37044
rect 34468 36988 36540 37044
rect 36596 36988 36606 37044
rect 36866 36988 36876 37044
rect 36932 36988 37436 37044
rect 37492 36988 37502 37044
rect 39666 36988 39676 37044
rect 39732 36988 43708 37044
rect 43764 36988 43774 37044
rect 46610 36988 46620 37044
rect 46676 36988 48748 37044
rect 48804 36988 49308 37044
rect 49364 36988 50204 37044
rect 50260 36988 51548 37044
rect 51604 36988 51614 37044
rect 52882 36988 52892 37044
rect 52948 36988 54012 37044
rect 54068 36988 54078 37044
rect 59602 36988 59612 37044
rect 59668 36988 60620 37044
rect 60676 36988 60686 37044
rect 5058 36876 5068 36932
rect 5124 36876 5516 36932
rect 5572 36876 15148 36932
rect 20738 36876 20748 36932
rect 20804 36876 22428 36932
rect 22484 36876 23660 36932
rect 23716 36876 23726 36932
rect 25666 36876 25676 36932
rect 25732 36876 26572 36932
rect 26628 36876 26638 36932
rect 36194 36876 36204 36932
rect 36260 36876 36652 36932
rect 36708 36876 36718 36932
rect 37202 36876 37212 36932
rect 37268 36876 37996 36932
rect 38052 36876 38062 36932
rect 41682 36876 41692 36932
rect 41748 36876 47180 36932
rect 47236 36876 47246 36932
rect 47404 36876 53340 36932
rect 53396 36876 53406 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 15092 36820 15148 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 47404 36820 47460 36876
rect 11890 36764 11900 36820
rect 11956 36764 11966 36820
rect 15092 36764 18620 36820
rect 18676 36764 18686 36820
rect 41010 36764 41020 36820
rect 41076 36764 41356 36820
rect 41412 36764 41422 36820
rect 45714 36764 45724 36820
rect 45780 36764 47460 36820
rect 48178 36764 48188 36820
rect 48244 36764 50204 36820
rect 50260 36764 50988 36820
rect 51044 36764 51054 36820
rect 53218 36764 53228 36820
rect 53284 36764 53788 36820
rect 53844 36764 53854 36820
rect 59266 36764 59276 36820
rect 59332 36764 61740 36820
rect 61796 36764 61964 36820
rect 62020 36764 62030 36820
rect 11900 36708 11956 36764
rect 6514 36652 6524 36708
rect 6580 36652 7196 36708
rect 7252 36652 7262 36708
rect 11900 36652 14700 36708
rect 14756 36652 15148 36708
rect 15204 36652 15214 36708
rect 20290 36652 20300 36708
rect 20356 36652 25452 36708
rect 25508 36652 25518 36708
rect 47842 36652 47852 36708
rect 47908 36652 49084 36708
rect 49140 36652 49150 36708
rect 49410 36652 49420 36708
rect 49476 36652 50540 36708
rect 50596 36652 50606 36708
rect 54898 36652 54908 36708
rect 54964 36652 55132 36708
rect 55188 36652 57372 36708
rect 57428 36652 57438 36708
rect 3042 36540 3052 36596
rect 3108 36540 14140 36596
rect 14196 36540 15372 36596
rect 15428 36540 15438 36596
rect 17154 36540 17164 36596
rect 17220 36540 17500 36596
rect 17556 36540 17566 36596
rect 20514 36540 20524 36596
rect 20580 36540 23996 36596
rect 24052 36540 24062 36596
rect 27010 36540 27020 36596
rect 27076 36540 27916 36596
rect 27972 36540 27982 36596
rect 39778 36540 39788 36596
rect 39844 36540 42364 36596
rect 42420 36540 42430 36596
rect 42690 36540 42700 36596
rect 42756 36540 45276 36596
rect 45332 36540 46172 36596
rect 46228 36540 46238 36596
rect 52210 36540 52220 36596
rect 52276 36540 52892 36596
rect 52948 36540 52958 36596
rect 56018 36540 56028 36596
rect 56084 36540 61068 36596
rect 61124 36540 61964 36596
rect 62020 36540 62030 36596
rect 2146 36428 2156 36484
rect 2212 36428 2828 36484
rect 2884 36428 2894 36484
rect 10098 36428 10108 36484
rect 10164 36428 11004 36484
rect 11060 36428 11564 36484
rect 11620 36428 11630 36484
rect 13570 36428 13580 36484
rect 13636 36428 20300 36484
rect 20356 36428 20366 36484
rect 21634 36428 21644 36484
rect 21700 36428 22316 36484
rect 22372 36428 22382 36484
rect 28242 36428 28252 36484
rect 28308 36428 31612 36484
rect 31668 36428 31678 36484
rect 34962 36428 34972 36484
rect 35028 36428 35644 36484
rect 35700 36428 37772 36484
rect 37828 36428 41020 36484
rect 41076 36428 41086 36484
rect 42018 36428 42028 36484
rect 42084 36428 43596 36484
rect 43652 36428 44828 36484
rect 44884 36428 45612 36484
rect 45668 36428 45678 36484
rect 51874 36428 51884 36484
rect 51940 36428 52780 36484
rect 52836 36428 52846 36484
rect 53106 36428 53116 36484
rect 53172 36428 54012 36484
rect 54068 36428 54078 36484
rect 56690 36428 56700 36484
rect 56756 36428 57260 36484
rect 57316 36428 57326 36484
rect 60050 36428 60060 36484
rect 60116 36428 60956 36484
rect 61012 36428 61022 36484
rect 61254 36428 61292 36484
rect 61348 36428 61358 36484
rect 2380 36316 4396 36372
rect 4452 36316 5628 36372
rect 5684 36316 5694 36372
rect 16034 36316 16044 36372
rect 16100 36316 18508 36372
rect 18564 36316 18574 36372
rect 20626 36316 20636 36372
rect 20692 36316 21980 36372
rect 22036 36316 24332 36372
rect 24388 36316 24398 36372
rect 34850 36316 34860 36372
rect 34916 36316 35756 36372
rect 35812 36316 36428 36372
rect 36484 36316 36494 36372
rect 39778 36316 39788 36372
rect 39844 36316 40908 36372
rect 40964 36316 40974 36372
rect 50866 36316 50876 36372
rect 50932 36316 51772 36372
rect 51828 36316 51838 36372
rect 54786 36316 54796 36372
rect 54852 36316 61516 36372
rect 61572 36316 61582 36372
rect 2380 36260 2436 36316
rect 2370 36204 2380 36260
rect 2436 36204 2446 36260
rect 2594 36204 2604 36260
rect 2660 36204 3948 36260
rect 4004 36204 4014 36260
rect 5842 36204 5852 36260
rect 5908 36204 8876 36260
rect 8932 36204 8942 36260
rect 12114 36204 12124 36260
rect 12180 36204 13916 36260
rect 13972 36204 14924 36260
rect 14980 36204 14990 36260
rect 16258 36204 16268 36260
rect 16324 36204 18284 36260
rect 18340 36204 18350 36260
rect 21522 36204 21532 36260
rect 21588 36204 22876 36260
rect 22932 36204 25676 36260
rect 25732 36204 25742 36260
rect 31042 36204 31052 36260
rect 31108 36204 33068 36260
rect 33124 36204 33134 36260
rect 35410 36204 35420 36260
rect 35476 36204 36652 36260
rect 36708 36204 37884 36260
rect 37940 36204 37950 36260
rect 38322 36204 38332 36260
rect 38388 36204 42924 36260
rect 42980 36204 42990 36260
rect 46050 36204 46060 36260
rect 46116 36204 46396 36260
rect 46452 36204 52220 36260
rect 52276 36204 53228 36260
rect 53284 36204 53294 36260
rect 58370 36204 58380 36260
rect 58436 36204 60508 36260
rect 60564 36204 60574 36260
rect 1474 36092 1484 36148
rect 1540 36092 17612 36148
rect 17668 36092 18396 36148
rect 18452 36092 18462 36148
rect 27794 36092 27804 36148
rect 27860 36092 30380 36148
rect 30436 36092 31948 36148
rect 32004 36092 32014 36148
rect 35074 36092 35084 36148
rect 35140 36092 36204 36148
rect 36260 36092 36270 36148
rect 40114 36092 40124 36148
rect 40180 36092 42812 36148
rect 42868 36092 42878 36148
rect 48038 36092 48076 36148
rect 48132 36092 48142 36148
rect 53106 36092 53116 36148
rect 53172 36092 53564 36148
rect 53620 36092 53630 36148
rect 56466 36092 56476 36148
rect 56532 36092 60844 36148
rect 60900 36092 61628 36148
rect 61684 36092 61694 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 53564 36036 53620 36092
rect 1698 35980 1708 36036
rect 1764 35980 5404 36036
rect 5460 35980 5470 36036
rect 7196 35980 11788 36036
rect 12338 35980 12348 36036
rect 12404 35980 15148 36036
rect 15204 35980 19292 36036
rect 19348 35980 19358 36036
rect 38098 35980 38108 36036
rect 38164 35980 40404 36036
rect 41010 35980 41020 36036
rect 41076 35980 44380 36036
rect 44436 35980 44446 36036
rect 44940 35980 50428 36036
rect 53564 35980 57540 36036
rect 58482 35980 58492 36036
rect 58548 35980 60732 36036
rect 60788 35980 60798 36036
rect 7196 35924 7252 35980
rect 11732 35924 11788 35980
rect 7186 35868 7196 35924
rect 7252 35868 7262 35924
rect 8866 35868 8876 35924
rect 8932 35868 11228 35924
rect 11284 35868 11294 35924
rect 11732 35868 16828 35924
rect 16884 35868 16894 35924
rect 35410 35868 35420 35924
rect 35476 35868 39900 35924
rect 39956 35868 39966 35924
rect 40348 35812 40404 35980
rect 44940 35924 44996 35980
rect 40674 35868 40684 35924
rect 40740 35868 43484 35924
rect 43540 35868 43550 35924
rect 43922 35868 43932 35924
rect 43988 35868 44996 35924
rect 45126 35868 45164 35924
rect 45220 35868 45230 35924
rect 50372 35812 50428 35980
rect 57484 35924 57540 35980
rect 52658 35868 52668 35924
rect 52724 35868 53004 35924
rect 53060 35868 57260 35924
rect 57316 35868 57326 35924
rect 57484 35868 62188 35924
rect 62244 35868 62254 35924
rect 3332 35756 4284 35812
rect 4340 35756 4350 35812
rect 7074 35756 7084 35812
rect 7140 35756 7756 35812
rect 7812 35756 7822 35812
rect 7970 35756 7980 35812
rect 8036 35756 10780 35812
rect 10836 35756 10846 35812
rect 10994 35756 11004 35812
rect 11060 35756 12012 35812
rect 12068 35756 12078 35812
rect 37986 35756 37996 35812
rect 38052 35756 38556 35812
rect 38612 35756 39788 35812
rect 39844 35756 39854 35812
rect 40338 35756 40348 35812
rect 40404 35756 45052 35812
rect 45108 35756 45118 35812
rect 46834 35756 46844 35812
rect 46900 35756 47628 35812
rect 47684 35756 47694 35812
rect 50372 35756 57596 35812
rect 57652 35756 57662 35812
rect 3332 35476 3388 35756
rect 7410 35644 7420 35700
rect 7476 35644 8540 35700
rect 8596 35644 8606 35700
rect 9762 35644 9772 35700
rect 9828 35644 10668 35700
rect 10724 35644 10734 35700
rect 15586 35644 15596 35700
rect 15652 35644 18844 35700
rect 18900 35644 18910 35700
rect 19618 35644 19628 35700
rect 19684 35644 20972 35700
rect 21028 35644 21038 35700
rect 22418 35644 22428 35700
rect 22484 35644 23212 35700
rect 23268 35644 23278 35700
rect 23538 35644 23548 35700
rect 23604 35644 25228 35700
rect 25284 35644 25294 35700
rect 34402 35644 34412 35700
rect 34468 35644 37100 35700
rect 37156 35644 37166 35700
rect 37426 35644 37436 35700
rect 37492 35644 38780 35700
rect 38836 35644 38846 35700
rect 42354 35644 42364 35700
rect 42420 35644 43148 35700
rect 43204 35644 43214 35700
rect 44258 35644 44268 35700
rect 44324 35644 44940 35700
rect 44996 35644 45612 35700
rect 45668 35644 45678 35700
rect 47170 35644 47180 35700
rect 47236 35644 47852 35700
rect 47908 35644 47918 35700
rect 49410 35644 49420 35700
rect 49476 35644 51996 35700
rect 52052 35644 52062 35700
rect 52882 35644 52892 35700
rect 52948 35644 53340 35700
rect 53396 35644 53406 35700
rect 54338 35644 54348 35700
rect 54404 35644 58828 35700
rect 58884 35644 58894 35700
rect 15250 35532 15260 35588
rect 15316 35532 20860 35588
rect 20916 35532 20926 35588
rect 21858 35532 21868 35588
rect 21924 35532 24444 35588
rect 24500 35532 24510 35588
rect 28130 35532 28140 35588
rect 28196 35532 29372 35588
rect 29428 35532 29438 35588
rect 41458 35532 41468 35588
rect 41524 35532 42476 35588
rect 42532 35532 45164 35588
rect 45220 35532 45230 35588
rect 47730 35532 47740 35588
rect 47796 35532 50988 35588
rect 51044 35532 51054 35588
rect 52770 35532 52780 35588
rect 52836 35532 54012 35588
rect 54068 35532 54078 35588
rect 55570 35532 55580 35588
rect 55636 35532 56700 35588
rect 56756 35532 56766 35588
rect 3042 35420 3052 35476
rect 3108 35420 3388 35476
rect 17042 35420 17052 35476
rect 17108 35420 23548 35476
rect 23604 35420 23614 35476
rect 42914 35420 42924 35476
rect 42980 35420 45836 35476
rect 45892 35420 45902 35476
rect 48850 35420 48860 35476
rect 48916 35420 52332 35476
rect 52388 35420 52398 35476
rect 54450 35420 54460 35476
rect 54516 35420 55692 35476
rect 55748 35420 55758 35476
rect 7634 35308 7644 35364
rect 7700 35308 8484 35364
rect 17154 35308 17164 35364
rect 17220 35308 17612 35364
rect 17668 35308 17678 35364
rect 38612 35308 39564 35364
rect 39620 35308 39630 35364
rect 39890 35308 39900 35364
rect 39956 35308 40124 35364
rect 40180 35308 40190 35364
rect 42018 35308 42028 35364
rect 42084 35308 42812 35364
rect 42868 35308 44268 35364
rect 44324 35308 44334 35364
rect 49298 35308 49308 35364
rect 49364 35308 49868 35364
rect 49924 35308 49934 35364
rect 54786 35308 54796 35364
rect 54852 35308 55244 35364
rect 55300 35308 55310 35364
rect 55906 35308 55916 35364
rect 55972 35308 57260 35364
rect 57316 35308 57326 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 8428 35252 8484 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 38612 35252 38668 35308
rect 6738 35196 6748 35252
rect 6804 35196 7420 35252
rect 7476 35196 7486 35252
rect 8428 35196 9884 35252
rect 9940 35196 15372 35252
rect 15428 35196 15438 35252
rect 28018 35196 28028 35252
rect 28084 35196 29820 35252
rect 29876 35196 32956 35252
rect 33012 35196 33022 35252
rect 36204 35196 38668 35252
rect 45154 35196 45164 35252
rect 45220 35196 49196 35252
rect 49252 35196 50428 35252
rect 50484 35196 51212 35252
rect 51268 35196 51278 35252
rect 53778 35196 53788 35252
rect 53844 35196 55468 35252
rect 55524 35196 55534 35252
rect 55794 35196 55804 35252
rect 55860 35196 56812 35252
rect 56868 35196 56878 35252
rect 57474 35196 57484 35252
rect 57540 35196 61292 35252
rect 61348 35196 61358 35252
rect 36204 35140 36260 35196
rect 10546 35084 10556 35140
rect 10612 35084 34076 35140
rect 34132 35084 34142 35140
rect 36194 35084 36204 35140
rect 36260 35084 36270 35140
rect 38612 35084 39340 35140
rect 39396 35084 40572 35140
rect 40628 35084 40638 35140
rect 41906 35084 41916 35140
rect 41972 35084 53004 35140
rect 53060 35084 53070 35140
rect 53554 35084 53564 35140
rect 53620 35084 55580 35140
rect 55636 35084 55646 35140
rect 56018 35084 56028 35140
rect 56084 35084 56252 35140
rect 56308 35084 56318 35140
rect 58034 35084 58044 35140
rect 58100 35084 58716 35140
rect 58772 35084 58782 35140
rect 38612 35028 38668 35084
rect 2146 34972 2156 35028
rect 2212 34972 4172 35028
rect 4228 34972 4238 35028
rect 6738 34972 6748 35028
rect 6804 34972 7532 35028
rect 7588 34972 11004 35028
rect 11060 34972 11070 35028
rect 15820 34972 19964 35028
rect 20020 34972 20030 35028
rect 22530 34972 22540 35028
rect 22596 34972 26572 35028
rect 26628 34972 26638 35028
rect 28466 34972 28476 35028
rect 28532 34972 29596 35028
rect 29652 34972 29662 35028
rect 35298 34972 35308 35028
rect 35364 34972 38668 35028
rect 50372 34972 51772 35028
rect 51828 34972 51838 35028
rect 53442 34972 53452 35028
rect 53508 34972 54908 35028
rect 54964 34972 54974 35028
rect 55682 34972 55692 35028
rect 55748 34972 59668 35028
rect 15820 34916 15876 34972
rect 50372 34916 50428 34972
rect 59612 34916 59668 34972
rect 2482 34860 2492 34916
rect 2548 34860 6188 34916
rect 6244 34860 6254 34916
rect 7298 34860 7308 34916
rect 7364 34860 8092 34916
rect 8148 34860 8652 34916
rect 8708 34860 8718 34916
rect 9650 34860 9660 34916
rect 9716 34860 9996 34916
rect 10052 34860 10062 34916
rect 11732 34860 15876 34916
rect 16034 34860 16044 34916
rect 16100 34860 18620 34916
rect 18676 34860 18686 34916
rect 28578 34860 28588 34916
rect 28644 34860 29932 34916
rect 29988 34860 29998 34916
rect 37538 34860 37548 34916
rect 37604 34860 38220 34916
rect 38276 34860 39564 34916
rect 39620 34860 40012 34916
rect 40068 34860 40078 34916
rect 41570 34860 41580 34916
rect 41636 34860 42700 34916
rect 42756 34860 42766 34916
rect 48738 34860 48748 34916
rect 48804 34860 49980 34916
rect 50036 34860 50428 34916
rect 53666 34860 53676 34916
rect 53732 34860 54572 34916
rect 54628 34860 54638 34916
rect 56018 34860 56028 34916
rect 56084 34860 56924 34916
rect 56980 34860 56990 34916
rect 59602 34860 59612 34916
rect 59668 34860 60732 34916
rect 60788 34860 60798 34916
rect 2594 34748 2604 34804
rect 2660 34748 3612 34804
rect 3668 34748 5964 34804
rect 6020 34748 6030 34804
rect 6290 34748 6300 34804
rect 6356 34748 6860 34804
rect 6916 34748 7868 34804
rect 7924 34748 8540 34804
rect 8596 34748 8606 34804
rect 11732 34692 11788 34860
rect 20738 34748 20748 34804
rect 20804 34748 27356 34804
rect 27412 34748 27422 34804
rect 27542 34748 27580 34804
rect 27636 34748 27646 34804
rect 28130 34748 28140 34804
rect 28196 34748 31836 34804
rect 31892 34748 31902 34804
rect 42018 34748 42028 34804
rect 42084 34748 42476 34804
rect 42532 34748 42542 34804
rect 56578 34748 56588 34804
rect 56644 34748 62188 34804
rect 62132 34692 62188 34748
rect 8306 34636 8316 34692
rect 8372 34636 8652 34692
rect 8708 34636 8718 34692
rect 9426 34636 9436 34692
rect 9492 34636 11788 34692
rect 13794 34636 13804 34692
rect 13860 34636 14812 34692
rect 14868 34636 14878 34692
rect 16818 34636 16828 34692
rect 16884 34636 18396 34692
rect 18452 34636 18462 34692
rect 20066 34636 20076 34692
rect 20132 34636 21420 34692
rect 21476 34636 21486 34692
rect 27094 34636 27132 34692
rect 27188 34636 27198 34692
rect 29334 34636 29372 34692
rect 29428 34636 29438 34692
rect 36082 34636 36092 34692
rect 36148 34636 36876 34692
rect 36932 34636 36942 34692
rect 41122 34636 41132 34692
rect 41188 34636 42812 34692
rect 42868 34636 43596 34692
rect 43652 34636 43662 34692
rect 45602 34636 45612 34692
rect 45668 34636 46508 34692
rect 46564 34636 46574 34692
rect 50372 34636 56252 34692
rect 56308 34636 56318 34692
rect 56914 34636 56924 34692
rect 56980 34636 58268 34692
rect 58324 34636 58334 34692
rect 62132 34636 62972 34692
rect 63028 34636 63038 34692
rect 2146 34524 2156 34580
rect 2212 34524 4844 34580
rect 4900 34524 5628 34580
rect 5684 34524 5694 34580
rect 7746 34524 7756 34580
rect 7812 34524 9100 34580
rect 9156 34524 10444 34580
rect 10500 34524 10510 34580
rect 15092 34524 17892 34580
rect 37202 34524 37212 34580
rect 37268 34524 43484 34580
rect 43540 34524 43550 34580
rect 15092 34468 15148 34524
rect 17836 34468 17892 34524
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50372 34468 50428 34636
rect 54338 34524 54348 34580
rect 54404 34524 57036 34580
rect 57092 34524 57102 34580
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 1922 34412 1932 34468
rect 1988 34412 15148 34468
rect 15334 34412 15372 34468
rect 15428 34412 15438 34468
rect 17826 34412 17836 34468
rect 17892 34412 17902 34468
rect 36530 34412 36540 34468
rect 36596 34412 37324 34468
rect 37380 34412 38668 34468
rect 38724 34412 38734 34468
rect 38882 34412 38892 34468
rect 38948 34412 39900 34468
rect 39956 34412 39966 34468
rect 41234 34412 41244 34468
rect 41300 34412 50428 34468
rect 2370 34300 2380 34356
rect 2436 34300 2940 34356
rect 2996 34300 3006 34356
rect 10210 34300 10220 34356
rect 10276 34300 11788 34356
rect 11844 34300 11854 34356
rect 14018 34300 14028 34356
rect 14084 34300 17276 34356
rect 17332 34300 17342 34356
rect 29250 34300 29260 34356
rect 29316 34300 29652 34356
rect 32386 34300 32396 34356
rect 32452 34300 33180 34356
rect 33236 34300 33246 34356
rect 36092 34300 40348 34356
rect 40404 34300 40414 34356
rect 42018 34300 42028 34356
rect 42084 34300 45836 34356
rect 45892 34300 45902 34356
rect 46834 34300 46844 34356
rect 46900 34300 48188 34356
rect 48244 34300 48254 34356
rect 50418 34300 50428 34356
rect 50484 34300 57148 34356
rect 57204 34300 57214 34356
rect 3378 34188 3388 34244
rect 3444 34188 3612 34244
rect 3668 34188 3678 34244
rect 15260 34188 17500 34244
rect 17556 34188 17566 34244
rect 18162 34188 18172 34244
rect 18228 34188 23324 34244
rect 23380 34188 23390 34244
rect 24546 34188 24556 34244
rect 24612 34188 25676 34244
rect 25732 34188 29372 34244
rect 29428 34188 29438 34244
rect 15260 34132 15316 34188
rect 29596 34132 29652 34300
rect 36092 34244 36148 34300
rect 35522 34188 35532 34244
rect 35588 34188 35868 34244
rect 35924 34188 36092 34244
rect 36148 34188 36158 34244
rect 39330 34188 39340 34244
rect 39396 34188 39788 34244
rect 39844 34188 40908 34244
rect 40964 34188 42588 34244
rect 42644 34188 42654 34244
rect 46946 34188 46956 34244
rect 47012 34188 49084 34244
rect 49140 34188 49150 34244
rect 59378 34188 59388 34244
rect 59444 34188 60732 34244
rect 60788 34188 61740 34244
rect 61796 34188 61806 34244
rect 62850 34188 62860 34244
rect 62916 34188 62926 34244
rect 62860 34132 62916 34188
rect 7746 34076 7756 34132
rect 7812 34076 10556 34132
rect 10612 34076 10622 34132
rect 15026 34076 15036 34132
rect 15092 34076 15316 34132
rect 15810 34076 15820 34132
rect 15876 34076 17612 34132
rect 17668 34076 17678 34132
rect 23426 34076 23436 34132
rect 23492 34076 29652 34132
rect 36306 34076 36316 34132
rect 36372 34076 37212 34132
rect 37268 34076 37278 34132
rect 37986 34076 37996 34132
rect 38052 34076 40796 34132
rect 40852 34076 40862 34132
rect 42130 34076 42140 34132
rect 42196 34076 43484 34132
rect 43540 34076 43550 34132
rect 44146 34076 44156 34132
rect 44212 34076 44492 34132
rect 44548 34076 47180 34132
rect 47236 34076 47246 34132
rect 50166 34076 50204 34132
rect 50260 34076 50270 34132
rect 50372 34076 53788 34132
rect 53844 34076 53854 34132
rect 54002 34076 54012 34132
rect 54068 34076 62916 34132
rect 2034 33964 2044 34020
rect 2100 33964 2492 34020
rect 2548 33964 4060 34020
rect 4116 33964 4126 34020
rect 6402 33964 6412 34020
rect 6468 33964 8428 34020
rect 8484 33964 8494 34020
rect 16604 33964 23548 34020
rect 24322 33964 24332 34020
rect 24388 33964 25788 34020
rect 25844 33964 25854 34020
rect 26852 33964 28140 34020
rect 28196 33964 28206 34020
rect 37874 33964 37884 34020
rect 37940 33964 38892 34020
rect 38948 33964 38958 34020
rect 40002 33964 40012 34020
rect 40068 33964 41356 34020
rect 41412 33964 43708 34020
rect 43764 33964 43774 34020
rect 45714 33964 45724 34020
rect 45780 33964 46284 34020
rect 46340 33964 46350 34020
rect 1362 33852 1372 33908
rect 1428 33852 7084 33908
rect 7140 33852 7150 33908
rect 8978 33852 8988 33908
rect 9044 33852 10276 33908
rect 13234 33852 13244 33908
rect 13300 33852 16044 33908
rect 16100 33852 16110 33908
rect 10220 33796 10276 33852
rect 16604 33796 16660 33964
rect 17826 33852 17836 33908
rect 17892 33852 18172 33908
rect 18228 33852 18238 33908
rect 22082 33852 22092 33908
rect 22148 33852 22876 33908
rect 22932 33852 22942 33908
rect 23492 33796 23548 33964
rect 26852 33908 26908 33964
rect 50372 33908 50428 34076
rect 50978 33964 50988 34020
rect 51044 33964 51660 34020
rect 51716 33964 51726 34020
rect 51986 33964 51996 34020
rect 52052 33964 53900 34020
rect 53956 33964 53966 34020
rect 23650 33852 23660 33908
rect 23716 33852 26908 33908
rect 28018 33852 28028 33908
rect 28084 33852 28094 33908
rect 37090 33852 37100 33908
rect 37156 33852 39340 33908
rect 39396 33852 39406 33908
rect 40338 33852 40348 33908
rect 40404 33852 41132 33908
rect 41188 33852 41580 33908
rect 41636 33852 42140 33908
rect 42196 33852 42206 33908
rect 48178 33852 48188 33908
rect 48244 33852 48972 33908
rect 49028 33852 50428 33908
rect 28028 33796 28084 33852
rect 54124 33796 54180 34076
rect 57026 33852 57036 33908
rect 57092 33852 59612 33908
rect 59668 33852 59678 33908
rect 8194 33740 8204 33796
rect 8260 33740 9996 33796
rect 10052 33740 10062 33796
rect 10220 33740 16660 33796
rect 16818 33740 16828 33796
rect 16884 33740 17388 33796
rect 17444 33740 18508 33796
rect 18564 33740 19292 33796
rect 19348 33740 19358 33796
rect 23492 33740 24444 33796
rect 24500 33740 24510 33796
rect 24780 33740 28084 33796
rect 37538 33740 37548 33796
rect 37604 33740 38220 33796
rect 38276 33740 38286 33796
rect 45826 33740 45836 33796
rect 45892 33740 54180 33796
rect 0 33684 800 33712
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 24780 33684 24836 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 0 33628 1764 33684
rect 0 33600 800 33628
rect 1708 33572 1764 33628
rect 5068 33628 12684 33684
rect 12740 33628 12750 33684
rect 17266 33628 17276 33684
rect 17332 33628 19852 33684
rect 19908 33628 19918 33684
rect 21074 33628 21084 33684
rect 21140 33628 23436 33684
rect 23492 33628 23502 33684
rect 24770 33628 24780 33684
rect 24836 33628 24846 33684
rect 24994 33628 25004 33684
rect 25060 33628 26460 33684
rect 26516 33628 26526 33684
rect 32470 33628 32508 33684
rect 32564 33628 32574 33684
rect 38658 33628 38668 33684
rect 38724 33628 43764 33684
rect 52098 33628 52108 33684
rect 52164 33628 53228 33684
rect 53284 33628 55020 33684
rect 55076 33628 55086 33684
rect 56102 33628 56140 33684
rect 56196 33628 56206 33684
rect 1708 33516 1932 33572
rect 1988 33516 1998 33572
rect 2146 33516 2156 33572
rect 2212 33516 2222 33572
rect 2706 33516 2716 33572
rect 2772 33516 4284 33572
rect 4340 33516 4350 33572
rect 2156 33124 2212 33516
rect 5068 33460 5124 33628
rect 43708 33572 43764 33628
rect 5954 33516 5964 33572
rect 6020 33516 6860 33572
rect 6916 33516 7644 33572
rect 7700 33516 7710 33572
rect 11330 33516 11340 33572
rect 11396 33516 13132 33572
rect 13188 33516 13198 33572
rect 13346 33516 13356 33572
rect 13412 33516 38668 33572
rect 39442 33516 39452 33572
rect 39508 33516 41020 33572
rect 41076 33516 41086 33572
rect 43708 33516 47068 33572
rect 47124 33516 47134 33572
rect 48626 33516 48636 33572
rect 48692 33516 50428 33572
rect 54226 33516 54236 33572
rect 54292 33516 54908 33572
rect 54964 33516 54974 33572
rect 55682 33516 55692 33572
rect 55748 33516 57148 33572
rect 57204 33516 60508 33572
rect 60564 33516 60574 33572
rect 38612 33460 38668 33516
rect 50372 33460 50428 33516
rect 4050 33404 4060 33460
rect 4116 33404 5124 33460
rect 7074 33404 7084 33460
rect 7140 33404 8092 33460
rect 8148 33404 10556 33460
rect 10612 33404 10622 33460
rect 12786 33404 12796 33460
rect 12852 33404 16940 33460
rect 16996 33404 19068 33460
rect 19124 33404 19134 33460
rect 26674 33404 26684 33460
rect 26740 33404 27804 33460
rect 27860 33404 28252 33460
rect 28308 33404 28318 33460
rect 29334 33404 29372 33460
rect 29428 33404 29438 33460
rect 31714 33404 31724 33460
rect 31780 33404 32732 33460
rect 32788 33404 32798 33460
rect 38612 33404 41692 33460
rect 41748 33404 45836 33460
rect 45892 33404 45902 33460
rect 47394 33404 47404 33460
rect 47460 33404 48860 33460
rect 48916 33404 50092 33460
rect 50148 33404 50158 33460
rect 50372 33404 55468 33460
rect 55524 33404 55534 33460
rect 4946 33292 4956 33348
rect 5012 33292 7196 33348
rect 7252 33292 7532 33348
rect 7588 33292 7598 33348
rect 8754 33292 8764 33348
rect 8820 33292 10220 33348
rect 10276 33292 10286 33348
rect 12338 33292 12348 33348
rect 12404 33292 15708 33348
rect 15764 33292 15774 33348
rect 16034 33292 16044 33348
rect 16100 33292 16380 33348
rect 16436 33292 16446 33348
rect 29922 33292 29932 33348
rect 29988 33292 30156 33348
rect 30212 33292 30828 33348
rect 30884 33292 30894 33348
rect 31826 33292 31836 33348
rect 31892 33292 33068 33348
rect 33124 33292 33134 33348
rect 33730 33292 33740 33348
rect 33796 33292 34412 33348
rect 34468 33292 34478 33348
rect 35410 33292 35420 33348
rect 35476 33292 38220 33348
rect 38276 33292 38286 33348
rect 44146 33292 44156 33348
rect 44212 33292 45724 33348
rect 45780 33292 45790 33348
rect 51314 33292 51324 33348
rect 51380 33292 51548 33348
rect 51604 33292 52892 33348
rect 52948 33292 52958 33348
rect 53330 33292 53340 33348
rect 53396 33292 53900 33348
rect 53956 33292 54684 33348
rect 54740 33292 54750 33348
rect 56242 33292 56252 33348
rect 56308 33292 56812 33348
rect 56868 33292 56878 33348
rect 58146 33292 58156 33348
rect 58212 33292 60732 33348
rect 60788 33292 60798 33348
rect 61394 33292 61404 33348
rect 61460 33292 61740 33348
rect 61796 33292 62412 33348
rect 62468 33292 62478 33348
rect 8530 33180 8540 33236
rect 8596 33180 10780 33236
rect 10836 33180 10846 33236
rect 19058 33180 19068 33236
rect 19124 33180 21868 33236
rect 21924 33180 21934 33236
rect 26002 33180 26012 33236
rect 26068 33180 28812 33236
rect 28868 33180 28878 33236
rect 32050 33180 32060 33236
rect 32116 33180 33292 33236
rect 33348 33180 34524 33236
rect 34580 33180 34590 33236
rect 37772 33180 40348 33236
rect 40404 33180 40414 33236
rect 43138 33180 43148 33236
rect 43204 33180 44268 33236
rect 44324 33180 44334 33236
rect 45042 33180 45052 33236
rect 45108 33180 46844 33236
rect 46900 33180 46910 33236
rect 48066 33180 48076 33236
rect 48132 33180 48748 33236
rect 48804 33180 49308 33236
rect 49364 33180 49374 33236
rect 52770 33180 52780 33236
rect 52836 33180 55804 33236
rect 55860 33180 60508 33236
rect 60564 33180 60574 33236
rect 37772 33124 37828 33180
rect 2146 33068 2156 33124
rect 2212 33068 2222 33124
rect 2370 33068 2380 33124
rect 2436 33068 4060 33124
rect 4116 33068 4126 33124
rect 7858 33068 7868 33124
rect 7924 33068 10220 33124
rect 10276 33068 10286 33124
rect 14214 33068 14252 33124
rect 14308 33068 14700 33124
rect 14756 33068 14766 33124
rect 15922 33068 15932 33124
rect 15988 33068 15998 33124
rect 18162 33068 18172 33124
rect 18228 33068 20748 33124
rect 20804 33068 24108 33124
rect 24164 33068 25004 33124
rect 25060 33068 25070 33124
rect 32162 33068 32172 33124
rect 32228 33068 36988 33124
rect 37044 33068 37054 33124
rect 37762 33068 37772 33124
rect 37828 33068 37838 33124
rect 41122 33068 41132 33124
rect 41188 33068 44044 33124
rect 44100 33068 44110 33124
rect 47842 33068 47852 33124
rect 47908 33068 50988 33124
rect 51044 33068 51054 33124
rect 10322 32956 10332 33012
rect 10388 32956 13804 33012
rect 13860 32956 13870 33012
rect 14476 32956 14588 33012
rect 14644 32956 14654 33012
rect 14476 32900 14532 32956
rect 5394 32844 5404 32900
rect 5460 32844 14924 32900
rect 14980 32844 14990 32900
rect 15932 32788 15988 33068
rect 63200 33012 64000 33040
rect 30482 32956 30492 33012
rect 30548 32956 31164 33012
rect 31220 32956 34412 33012
rect 34468 32956 36652 33012
rect 36708 32956 36718 33012
rect 61618 32956 61628 33012
rect 61684 32956 64000 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 63200 32928 64000 32956
rect 32162 32844 32172 32900
rect 32228 32844 35084 32900
rect 35140 32844 35532 32900
rect 35588 32844 35598 32900
rect 5282 32732 5292 32788
rect 5348 32732 11844 32788
rect 12002 32732 12012 32788
rect 12068 32732 16324 32788
rect 25778 32732 25788 32788
rect 25844 32732 28252 32788
rect 28308 32732 28318 32788
rect 28802 32732 28812 32788
rect 28868 32732 29932 32788
rect 29988 32732 29998 32788
rect 33506 32732 33516 32788
rect 33572 32732 36092 32788
rect 36148 32732 36158 32788
rect 38770 32732 38780 32788
rect 38836 32732 39788 32788
rect 39844 32732 39854 32788
rect 49186 32732 49196 32788
rect 49252 32732 52220 32788
rect 52276 32732 52286 32788
rect 56802 32732 56812 32788
rect 56868 32732 57484 32788
rect 57540 32732 57550 32788
rect 11788 32676 11844 32732
rect 1810 32620 1820 32676
rect 1876 32620 2268 32676
rect 2324 32620 2334 32676
rect 2482 32620 2492 32676
rect 2548 32620 3612 32676
rect 3668 32620 4844 32676
rect 4900 32620 4910 32676
rect 5842 32620 5852 32676
rect 5908 32620 6524 32676
rect 6580 32620 10108 32676
rect 10164 32620 10174 32676
rect 11788 32620 13356 32676
rect 13412 32620 13422 32676
rect 16268 32564 16324 32732
rect 16482 32620 16492 32676
rect 16548 32620 17388 32676
rect 17444 32620 17454 32676
rect 21410 32620 21420 32676
rect 21476 32620 22316 32676
rect 22372 32620 22876 32676
rect 22932 32620 25228 32676
rect 25284 32620 25294 32676
rect 27906 32620 27916 32676
rect 27972 32620 28476 32676
rect 28532 32620 28542 32676
rect 37986 32620 37996 32676
rect 38052 32620 38556 32676
rect 38612 32620 39676 32676
rect 39732 32620 39742 32676
rect 49522 32620 49532 32676
rect 49588 32620 49598 32676
rect 4050 32508 4060 32564
rect 4116 32508 5964 32564
rect 6020 32508 6030 32564
rect 14914 32508 14924 32564
rect 14980 32508 16044 32564
rect 16100 32508 16110 32564
rect 16258 32508 16268 32564
rect 16324 32508 18508 32564
rect 18564 32508 18574 32564
rect 28914 32508 28924 32564
rect 28980 32508 29372 32564
rect 29428 32508 30380 32564
rect 30436 32508 31836 32564
rect 31892 32508 31902 32564
rect 33842 32508 33852 32564
rect 33908 32508 34356 32564
rect 37650 32508 37660 32564
rect 37716 32508 39452 32564
rect 39508 32508 39518 32564
rect 40114 32508 40124 32564
rect 40180 32508 42028 32564
rect 42084 32508 42094 32564
rect 45378 32508 45388 32564
rect 45444 32508 45454 32564
rect 34300 32452 34356 32508
rect 45388 32452 45444 32508
rect 49532 32452 49588 32620
rect 51202 32508 51212 32564
rect 51268 32508 51278 32564
rect 56466 32508 56476 32564
rect 56532 32508 58492 32564
rect 58548 32508 58558 32564
rect 60498 32508 60508 32564
rect 60564 32508 61180 32564
rect 61236 32508 61246 32564
rect 51212 32452 51268 32508
rect 1810 32396 1820 32452
rect 1876 32396 2380 32452
rect 2436 32396 4172 32452
rect 4228 32396 4508 32452
rect 4564 32396 4574 32452
rect 12562 32396 12572 32452
rect 12628 32396 13356 32452
rect 13412 32396 13422 32452
rect 15474 32396 15484 32452
rect 15540 32396 16380 32452
rect 16436 32396 17612 32452
rect 17668 32396 17678 32452
rect 18722 32396 18732 32452
rect 18788 32396 20860 32452
rect 20916 32396 20926 32452
rect 32470 32396 32508 32452
rect 32564 32396 33068 32452
rect 33124 32396 33134 32452
rect 34290 32396 34300 32452
rect 34356 32396 34366 32452
rect 34514 32396 34524 32452
rect 34580 32396 37884 32452
rect 37940 32396 39228 32452
rect 39284 32396 39294 32452
rect 41682 32396 41692 32452
rect 41748 32396 43148 32452
rect 43204 32396 43214 32452
rect 45388 32396 51268 32452
rect 51986 32396 51996 32452
rect 52052 32396 52780 32452
rect 52836 32396 52846 32452
rect 53666 32396 53676 32452
rect 53732 32396 54124 32452
rect 54180 32396 62076 32452
rect 62132 32396 62142 32452
rect 15484 32340 15540 32396
rect 11554 32284 11564 32340
rect 11620 32284 13132 32340
rect 13188 32284 15540 32340
rect 19058 32284 19068 32340
rect 19124 32284 21196 32340
rect 21252 32284 21262 32340
rect 35970 32284 35980 32340
rect 36036 32284 36204 32340
rect 36260 32284 37100 32340
rect 37156 32284 37166 32340
rect 48290 32284 48300 32340
rect 48356 32284 59724 32340
rect 59780 32284 59790 32340
rect 10882 32172 10892 32228
rect 10948 32172 12236 32228
rect 12292 32172 12302 32228
rect 17714 32172 17724 32228
rect 17780 32172 18060 32228
rect 18116 32172 18126 32228
rect 43810 32172 43820 32228
rect 43876 32172 56252 32228
rect 56308 32172 56318 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 3154 32060 3164 32116
rect 3220 32060 3500 32116
rect 3556 32060 3566 32116
rect 5170 32060 5180 32116
rect 5236 32060 9660 32116
rect 9716 32060 9726 32116
rect 10658 32060 10668 32116
rect 10724 32060 11228 32116
rect 11284 32060 11294 32116
rect 14018 32060 14028 32116
rect 14084 32060 23772 32116
rect 23828 32060 26012 32116
rect 26068 32060 26078 32116
rect 41682 32060 41692 32116
rect 41748 32060 43148 32116
rect 43204 32060 43932 32116
rect 43988 32060 49980 32116
rect 50036 32060 51100 32116
rect 51156 32060 51166 32116
rect 52994 32060 53004 32116
rect 53060 32060 56812 32116
rect 56868 32060 56878 32116
rect 2818 31948 2828 32004
rect 2884 31948 4732 32004
rect 4788 31948 4798 32004
rect 5058 31948 5068 32004
rect 5124 31948 6188 32004
rect 6244 31948 6254 32004
rect 8530 31948 8540 32004
rect 8596 31948 9772 32004
rect 9828 31948 9838 32004
rect 10892 31948 13020 32004
rect 13076 31948 13086 32004
rect 17052 31948 20412 32004
rect 20468 31948 20478 32004
rect 21858 31948 21868 32004
rect 21924 31948 22316 32004
rect 22372 31948 22382 32004
rect 22530 31948 22540 32004
rect 22596 31948 22606 32004
rect 24658 31948 24668 32004
rect 24724 31948 31948 32004
rect 32004 31948 32014 32004
rect 34178 31948 34188 32004
rect 34244 31948 34412 32004
rect 34468 31948 34478 32004
rect 42242 31948 42252 32004
rect 42308 31948 46508 32004
rect 46564 31948 46574 32004
rect 50530 31948 50540 32004
rect 50596 31948 51660 32004
rect 51716 31948 51726 32004
rect 52210 31948 52220 32004
rect 52276 31948 53564 32004
rect 53620 31948 53630 32004
rect 2930 31836 2940 31892
rect 2996 31836 9212 31892
rect 9268 31836 9278 31892
rect 10892 31780 10948 31948
rect 12226 31836 12236 31892
rect 12292 31836 12684 31892
rect 12740 31836 15260 31892
rect 15316 31836 15326 31892
rect 15586 31836 15596 31892
rect 15652 31836 16268 31892
rect 16324 31836 16334 31892
rect 2146 31724 2156 31780
rect 2212 31724 2828 31780
rect 2884 31724 2894 31780
rect 3938 31724 3948 31780
rect 4004 31724 4284 31780
rect 4340 31724 5516 31780
rect 5572 31724 5582 31780
rect 6402 31724 6412 31780
rect 6468 31724 8988 31780
rect 9044 31724 9054 31780
rect 9762 31724 9772 31780
rect 9828 31724 10948 31780
rect 14326 31724 14364 31780
rect 14420 31724 14430 31780
rect 14578 31724 14588 31780
rect 14644 31724 16828 31780
rect 16884 31724 16894 31780
rect 14364 31668 14420 31724
rect 3266 31612 3276 31668
rect 3332 31612 6188 31668
rect 6244 31612 6254 31668
rect 6822 31612 6860 31668
rect 6916 31612 6926 31668
rect 7718 31612 7756 31668
rect 7812 31612 7822 31668
rect 14364 31612 14700 31668
rect 14756 31612 14766 31668
rect 15138 31612 15148 31668
rect 15204 31612 16660 31668
rect 16604 31556 16660 31612
rect 17052 31556 17108 31948
rect 22540 31892 22596 31948
rect 22540 31836 23212 31892
rect 23268 31836 23278 31892
rect 24322 31836 24332 31892
rect 24388 31836 25564 31892
rect 25620 31836 25630 31892
rect 26226 31836 26236 31892
rect 26292 31836 28364 31892
rect 28420 31836 28430 31892
rect 28690 31836 28700 31892
rect 28756 31836 29708 31892
rect 29764 31836 30940 31892
rect 30996 31836 31006 31892
rect 34962 31836 34972 31892
rect 35028 31836 35980 31892
rect 36036 31836 37436 31892
rect 37492 31836 37502 31892
rect 37660 31836 39676 31892
rect 39732 31836 39742 31892
rect 43586 31836 43596 31892
rect 43652 31836 43932 31892
rect 43988 31836 44716 31892
rect 44772 31836 44782 31892
rect 45154 31836 45164 31892
rect 45220 31836 46284 31892
rect 46340 31836 48748 31892
rect 48804 31836 48814 31892
rect 52658 31836 52668 31892
rect 52724 31836 53340 31892
rect 53396 31836 53406 31892
rect 54562 31836 54572 31892
rect 54628 31836 55692 31892
rect 55748 31836 57484 31892
rect 57540 31836 57550 31892
rect 37660 31780 37716 31836
rect 45164 31780 45220 31836
rect 17826 31724 17836 31780
rect 17892 31724 20300 31780
rect 20356 31724 21532 31780
rect 21588 31724 22092 31780
rect 22148 31724 22158 31780
rect 22754 31724 22764 31780
rect 22820 31724 23996 31780
rect 24052 31724 24062 31780
rect 33730 31724 33740 31780
rect 33796 31724 35532 31780
rect 35588 31724 35598 31780
rect 36418 31724 36428 31780
rect 36484 31724 37716 31780
rect 38546 31724 38556 31780
rect 38612 31724 40684 31780
rect 40740 31724 40750 31780
rect 42242 31724 42252 31780
rect 42308 31724 43708 31780
rect 43764 31724 45220 31780
rect 53340 31780 53396 31836
rect 53340 31724 57820 31780
rect 57876 31724 58828 31780
rect 58884 31724 58894 31780
rect 60162 31724 60172 31780
rect 60228 31724 61628 31780
rect 61684 31724 61694 31780
rect 18498 31612 18508 31668
rect 18564 31612 21308 31668
rect 21364 31612 21374 31668
rect 21970 31612 21980 31668
rect 22036 31612 23548 31668
rect 23604 31612 23614 31668
rect 24546 31612 24556 31668
rect 24612 31612 25900 31668
rect 25956 31612 25966 31668
rect 30706 31612 30716 31668
rect 30772 31612 32396 31668
rect 32452 31612 32956 31668
rect 33012 31612 33022 31668
rect 34178 31612 34188 31668
rect 34244 31612 34524 31668
rect 34580 31612 34590 31668
rect 36306 31612 36316 31668
rect 36372 31612 37324 31668
rect 37380 31612 37390 31668
rect 42130 31612 42140 31668
rect 42196 31612 44156 31668
rect 44212 31612 62076 31668
rect 62132 31612 62142 31668
rect 3938 31500 3948 31556
rect 4004 31500 6972 31556
rect 7028 31500 7038 31556
rect 7410 31500 7420 31556
rect 7476 31500 9100 31556
rect 9156 31500 9166 31556
rect 9398 31500 9436 31556
rect 9492 31500 9502 31556
rect 10994 31500 11004 31556
rect 11060 31500 15148 31556
rect 15204 31500 15214 31556
rect 16594 31500 16604 31556
rect 16660 31500 17108 31556
rect 19628 31500 23100 31556
rect 23156 31500 23548 31556
rect 24322 31500 24332 31556
rect 24388 31500 26012 31556
rect 26068 31500 27692 31556
rect 27748 31500 27758 31556
rect 30258 31500 30268 31556
rect 30324 31500 31276 31556
rect 31332 31500 32732 31556
rect 32788 31500 33852 31556
rect 33908 31500 33918 31556
rect 34738 31500 34748 31556
rect 34804 31500 35756 31556
rect 35812 31500 38332 31556
rect 38388 31500 38398 31556
rect 41458 31500 41468 31556
rect 41524 31500 45276 31556
rect 45332 31500 46060 31556
rect 46116 31500 46126 31556
rect 48178 31500 48188 31556
rect 48244 31500 50988 31556
rect 51044 31500 51054 31556
rect 54450 31500 54460 31556
rect 54516 31500 55020 31556
rect 55076 31500 56252 31556
rect 56308 31500 56318 31556
rect 56578 31500 56588 31556
rect 56644 31500 57148 31556
rect 57204 31500 57596 31556
rect 57652 31500 57662 31556
rect 58370 31500 58380 31556
rect 58436 31500 61516 31556
rect 61572 31500 61582 31556
rect 6178 31388 6188 31444
rect 6244 31388 6860 31444
rect 6916 31388 8764 31444
rect 8820 31388 8830 31444
rect 12674 31388 12684 31444
rect 12740 31388 15036 31444
rect 15092 31388 16492 31444
rect 16548 31388 16558 31444
rect 16930 31388 16940 31444
rect 16996 31388 17500 31444
rect 17556 31388 17566 31444
rect 19628 31332 19684 31500
rect 23492 31444 23548 31500
rect 23492 31388 31948 31444
rect 32004 31388 32014 31444
rect 32834 31388 32844 31444
rect 32900 31388 41916 31444
rect 41972 31388 41982 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 4834 31276 4844 31332
rect 4900 31276 8540 31332
rect 8596 31276 8606 31332
rect 9650 31276 9660 31332
rect 9716 31276 12012 31332
rect 12068 31276 19684 31332
rect 52658 31276 52668 31332
rect 52724 31276 56588 31332
rect 56644 31276 57932 31332
rect 57988 31276 60508 31332
rect 60564 31276 60574 31332
rect 2156 31164 6636 31220
rect 6692 31164 6702 31220
rect 7970 31164 7980 31220
rect 8036 31164 8316 31220
rect 8372 31164 10108 31220
rect 10164 31164 10174 31220
rect 11666 31164 11676 31220
rect 11732 31164 12124 31220
rect 12180 31164 12190 31220
rect 12786 31164 12796 31220
rect 12852 31164 13468 31220
rect 13524 31164 13534 31220
rect 13794 31164 13804 31220
rect 13860 31164 15372 31220
rect 15428 31164 15438 31220
rect 16258 31164 16268 31220
rect 16324 31164 18732 31220
rect 18788 31164 18798 31220
rect 19058 31164 19068 31220
rect 19124 31164 23212 31220
rect 23268 31164 24556 31220
rect 24612 31164 24622 31220
rect 27234 31164 27244 31220
rect 27300 31164 28252 31220
rect 28308 31164 28318 31220
rect 30034 31164 30044 31220
rect 30100 31164 31164 31220
rect 31220 31164 31230 31220
rect 38770 31164 38780 31220
rect 38836 31164 40012 31220
rect 40068 31164 40078 31220
rect 44818 31164 44828 31220
rect 44884 31164 45948 31220
rect 46004 31164 46014 31220
rect 46274 31164 46284 31220
rect 46340 31164 47628 31220
rect 47684 31164 47694 31220
rect 51090 31164 51100 31220
rect 51156 31164 51436 31220
rect 51492 31164 51502 31220
rect 2156 31108 2212 31164
rect 19068 31108 19124 31164
rect 2146 31052 2156 31108
rect 2212 31052 2222 31108
rect 13682 31052 13692 31108
rect 13748 31052 14476 31108
rect 14532 31052 14542 31108
rect 14802 31052 14812 31108
rect 14868 31052 15148 31108
rect 15204 31052 15708 31108
rect 15764 31052 16716 31108
rect 16772 31052 16782 31108
rect 17826 31052 17836 31108
rect 17892 31052 19124 31108
rect 37650 31052 37660 31108
rect 37716 31052 40124 31108
rect 40180 31052 40190 31108
rect 50372 31052 52780 31108
rect 52836 31052 52846 31108
rect 53554 31052 53564 31108
rect 53620 31052 54572 31108
rect 54628 31052 54638 31108
rect 0 30996 800 31024
rect 50372 30996 50428 31052
rect 63200 30996 64000 31024
rect 0 30940 1596 30996
rect 1652 30940 1662 30996
rect 2706 30940 2716 30996
rect 2772 30940 3724 30996
rect 3780 30940 5852 30996
rect 5908 30940 7532 30996
rect 7588 30940 7598 30996
rect 7858 30940 7868 30996
rect 7924 30940 8876 30996
rect 8932 30940 8942 30996
rect 12450 30940 12460 30996
rect 12516 30940 12526 30996
rect 13122 30940 13132 30996
rect 13188 30940 14028 30996
rect 14084 30940 14094 30996
rect 16034 30940 16044 30996
rect 16100 30940 16492 30996
rect 16548 30940 18508 30996
rect 18564 30940 18574 30996
rect 21074 30940 21084 30996
rect 21140 30940 23100 30996
rect 23156 30940 23166 30996
rect 23762 30940 23772 30996
rect 23828 30940 24668 30996
rect 24724 30940 24734 30996
rect 27346 30940 27356 30996
rect 27412 30940 29596 30996
rect 29652 30940 29662 30996
rect 34188 30940 36540 30996
rect 36596 30940 36606 30996
rect 37090 30940 37100 30996
rect 37156 30940 38108 30996
rect 38164 30940 38174 30996
rect 48178 30940 48188 30996
rect 48244 30940 50428 30996
rect 51762 30940 51772 30996
rect 51828 30940 59612 30996
rect 59668 30940 59678 30996
rect 62132 30940 64000 30996
rect 0 30912 800 30940
rect 12460 30884 12516 30940
rect 34188 30884 34244 30940
rect 62132 30884 62188 30940
rect 63200 30912 64000 30940
rect 7074 30828 7084 30884
rect 7140 30828 10892 30884
rect 10948 30828 11228 30884
rect 11284 30828 12516 30884
rect 21298 30828 21308 30884
rect 21364 30828 22428 30884
rect 22484 30828 23660 30884
rect 23716 30828 23726 30884
rect 34178 30828 34188 30884
rect 34244 30828 34254 30884
rect 34402 30828 34412 30884
rect 34468 30828 37772 30884
rect 37828 30828 40908 30884
rect 40964 30828 40974 30884
rect 43250 30828 43260 30884
rect 43316 30828 44380 30884
rect 44436 30828 55020 30884
rect 55076 30828 55086 30884
rect 61954 30828 61964 30884
rect 62020 30828 62188 30884
rect 7634 30716 7644 30772
rect 7700 30716 8092 30772
rect 8148 30716 8158 30772
rect 20738 30716 20748 30772
rect 20804 30716 23212 30772
rect 23268 30716 23436 30772
rect 23492 30716 25676 30772
rect 25732 30716 25742 30772
rect 35634 30716 35644 30772
rect 35700 30716 41244 30772
rect 41300 30716 41310 30772
rect 51426 30716 51436 30772
rect 51492 30716 60284 30772
rect 60340 30716 60350 30772
rect 14018 30604 14028 30660
rect 14084 30604 28700 30660
rect 28756 30604 28766 30660
rect 34150 30604 34188 30660
rect 34244 30604 34254 30660
rect 37314 30604 37324 30660
rect 37380 30604 48076 30660
rect 48132 30604 48142 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 7074 30492 7084 30548
rect 7140 30492 7756 30548
rect 7812 30492 7822 30548
rect 20290 30492 20300 30548
rect 20356 30492 23548 30548
rect 23604 30492 24668 30548
rect 24724 30492 24734 30548
rect 46722 30492 46732 30548
rect 46788 30492 59276 30548
rect 59332 30492 59948 30548
rect 60004 30492 60014 30548
rect 1138 30380 1148 30436
rect 1204 30380 7756 30436
rect 7812 30380 7822 30436
rect 13682 30380 13692 30436
rect 13748 30380 14140 30436
rect 14196 30380 14206 30436
rect 23986 30380 23996 30436
rect 24052 30380 26908 30436
rect 27682 30380 27692 30436
rect 27748 30380 28476 30436
rect 28532 30380 29148 30436
rect 29204 30380 29214 30436
rect 43026 30380 43036 30436
rect 43092 30380 43932 30436
rect 43988 30380 43998 30436
rect 46610 30380 46620 30436
rect 46676 30380 51436 30436
rect 51492 30380 51502 30436
rect 56802 30380 56812 30436
rect 56868 30380 57708 30436
rect 57764 30380 57774 30436
rect 5618 30268 5628 30324
rect 5684 30268 7868 30324
rect 7924 30268 7934 30324
rect 19506 30268 19516 30324
rect 19572 30268 21420 30324
rect 21476 30268 21486 30324
rect 23202 30268 23212 30324
rect 23268 30268 25228 30324
rect 25284 30268 25294 30324
rect 25442 30268 25452 30324
rect 25508 30268 26012 30324
rect 26068 30268 26078 30324
rect 3826 30156 3836 30212
rect 3892 30156 5740 30212
rect 5796 30156 5806 30212
rect 6066 30156 6076 30212
rect 6132 30156 7308 30212
rect 7364 30156 7374 30212
rect 11554 30156 11564 30212
rect 11620 30156 12908 30212
rect 12964 30156 12974 30212
rect 19842 30156 19852 30212
rect 19908 30156 24388 30212
rect 24546 30156 24556 30212
rect 24612 30156 25564 30212
rect 25620 30156 25630 30212
rect 24332 30100 24388 30156
rect 26852 30100 26908 30380
rect 63200 30324 64000 30352
rect 30482 30268 30492 30324
rect 30548 30268 30940 30324
rect 30996 30268 31836 30324
rect 31892 30268 31902 30324
rect 40002 30268 40012 30324
rect 40068 30268 47404 30324
rect 47460 30268 47470 30324
rect 55458 30268 55468 30324
rect 55524 30268 57036 30324
rect 57092 30268 57102 30324
rect 61618 30268 61628 30324
rect 61684 30268 62636 30324
rect 62692 30268 62702 30324
rect 62962 30268 62972 30324
rect 63028 30268 64000 30324
rect 63200 30240 64000 30268
rect 33506 30156 33516 30212
rect 33572 30156 34412 30212
rect 34468 30156 34478 30212
rect 37986 30156 37996 30212
rect 38052 30156 41356 30212
rect 41412 30156 42252 30212
rect 42308 30156 42318 30212
rect 43362 30156 43372 30212
rect 43428 30156 44156 30212
rect 44212 30156 44222 30212
rect 46946 30156 46956 30212
rect 47012 30156 47628 30212
rect 47684 30156 47694 30212
rect 51874 30156 51884 30212
rect 51940 30156 52668 30212
rect 52724 30156 52734 30212
rect 53218 30156 53228 30212
rect 53284 30156 54124 30212
rect 54180 30156 54460 30212
rect 54516 30156 55132 30212
rect 55188 30156 55198 30212
rect 56018 30156 56028 30212
rect 56084 30156 56476 30212
rect 56532 30156 56542 30212
rect 60274 30156 60284 30212
rect 60340 30156 61068 30212
rect 61124 30156 61134 30212
rect 4722 30044 4732 30100
rect 4788 30044 7420 30100
rect 7476 30044 7486 30100
rect 8530 30044 8540 30100
rect 8596 30044 16380 30100
rect 16436 30044 16446 30100
rect 21858 30044 21868 30100
rect 21924 30044 23884 30100
rect 23940 30044 23950 30100
rect 24332 30044 26236 30100
rect 26292 30044 26302 30100
rect 26852 30044 27804 30100
rect 27860 30044 32060 30100
rect 32116 30044 33852 30100
rect 33908 30044 33918 30100
rect 34748 30044 38556 30100
rect 38612 30044 38622 30100
rect 41906 30044 41916 30100
rect 41972 30044 43820 30100
rect 43876 30044 43886 30100
rect 46060 30044 50204 30100
rect 50260 30044 53340 30100
rect 53396 30044 54236 30100
rect 54292 30044 54302 30100
rect 55570 30044 55580 30100
rect 55636 30044 56924 30100
rect 56980 30044 56990 30100
rect 59714 30044 59724 30100
rect 59780 30044 61404 30100
rect 61460 30044 61470 30100
rect 61618 30044 61628 30100
rect 61684 30044 62188 30100
rect 62244 30044 62254 30100
rect 34748 29988 34804 30044
rect 46060 29988 46116 30044
rect 3042 29932 3052 29988
rect 3108 29932 3500 29988
rect 3556 29932 6860 29988
rect 6916 29932 6926 29988
rect 20850 29932 20860 29988
rect 20916 29932 22204 29988
rect 22260 29932 22270 29988
rect 31938 29932 31948 29988
rect 32004 29932 34804 29988
rect 34962 29932 34972 29988
rect 35028 29932 35756 29988
rect 35812 29932 35822 29988
rect 37202 29932 37212 29988
rect 37268 29932 37436 29988
rect 37492 29932 38892 29988
rect 38948 29932 38958 29988
rect 39218 29932 39228 29988
rect 39284 29932 39788 29988
rect 39844 29932 40460 29988
rect 40516 29932 40526 29988
rect 43362 29932 43372 29988
rect 43428 29932 45052 29988
rect 45108 29932 45118 29988
rect 46050 29932 46060 29988
rect 46116 29932 46126 29988
rect 46386 29932 46396 29988
rect 46452 29932 55020 29988
rect 55076 29932 55086 29988
rect 55766 29932 55804 29988
rect 55860 29932 55870 29988
rect 56018 29932 56028 29988
rect 56084 29932 60508 29988
rect 60564 29932 60574 29988
rect 60946 29932 60956 29988
rect 61012 29932 62860 29988
rect 62916 29932 62926 29988
rect 20514 29820 20524 29876
rect 20580 29820 23884 29876
rect 23940 29820 23950 29876
rect 33730 29820 33740 29876
rect 33796 29820 35868 29876
rect 35924 29820 35934 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 3714 29708 3724 29764
rect 3780 29708 7196 29764
rect 7252 29708 7756 29764
rect 7812 29708 7822 29764
rect 25554 29708 25564 29764
rect 25620 29708 27244 29764
rect 27300 29708 27580 29764
rect 27636 29708 27646 29764
rect 63200 29652 64000 29680
rect 2034 29596 2044 29652
rect 2100 29596 4732 29652
rect 4788 29596 4798 29652
rect 9846 29596 9884 29652
rect 9940 29596 9950 29652
rect 16930 29596 16940 29652
rect 16996 29596 24332 29652
rect 24388 29596 24398 29652
rect 32386 29596 32396 29652
rect 32452 29596 33180 29652
rect 33236 29596 34580 29652
rect 35522 29596 35532 29652
rect 35588 29596 35980 29652
rect 36036 29596 36046 29652
rect 36642 29596 36652 29652
rect 36708 29596 37996 29652
rect 38052 29596 38062 29652
rect 38658 29596 38668 29652
rect 38724 29596 39340 29652
rect 39396 29596 39406 29652
rect 40114 29596 40124 29652
rect 40180 29596 41356 29652
rect 41412 29596 41422 29652
rect 59602 29596 59612 29652
rect 59668 29596 64000 29652
rect 34524 29540 34580 29596
rect 63200 29568 64000 29596
rect 16482 29484 16492 29540
rect 16548 29484 19180 29540
rect 19236 29484 19246 29540
rect 31266 29484 31276 29540
rect 31332 29484 33068 29540
rect 33124 29484 33134 29540
rect 34514 29484 34524 29540
rect 34580 29484 35084 29540
rect 35140 29484 35150 29540
rect 10098 29372 10108 29428
rect 10164 29372 13804 29428
rect 13860 29372 13870 29428
rect 14242 29372 14252 29428
rect 14308 29372 15260 29428
rect 15316 29372 16604 29428
rect 16660 29372 16670 29428
rect 19282 29372 19292 29428
rect 19348 29372 20748 29428
rect 20804 29372 21644 29428
rect 21700 29372 22652 29428
rect 22708 29372 23996 29428
rect 24052 29372 24062 29428
rect 24210 29372 24220 29428
rect 24276 29372 25004 29428
rect 25060 29372 25564 29428
rect 25620 29372 25630 29428
rect 26338 29372 26348 29428
rect 26404 29372 29036 29428
rect 29092 29372 29102 29428
rect 35252 29316 35308 29540
rect 35364 29484 36540 29540
rect 36596 29484 42476 29540
rect 42532 29484 44268 29540
rect 44324 29484 44334 29540
rect 48066 29484 48076 29540
rect 48132 29484 49756 29540
rect 49812 29484 49822 29540
rect 51202 29484 51212 29540
rect 51268 29484 52332 29540
rect 52388 29484 52398 29540
rect 55906 29484 55916 29540
rect 55972 29484 56924 29540
rect 56980 29484 56990 29540
rect 57596 29484 58828 29540
rect 58884 29484 60396 29540
rect 60452 29484 60462 29540
rect 57596 29428 57652 29484
rect 36418 29372 36428 29428
rect 36484 29372 37212 29428
rect 37268 29372 37278 29428
rect 40338 29372 40348 29428
rect 40404 29372 41244 29428
rect 41300 29372 41310 29428
rect 46050 29372 46060 29428
rect 46116 29372 47292 29428
rect 47348 29372 47358 29428
rect 47842 29372 47852 29428
rect 47908 29372 48860 29428
rect 48916 29372 48926 29428
rect 50530 29372 50540 29428
rect 50596 29372 52108 29428
rect 52164 29372 52174 29428
rect 54562 29372 54572 29428
rect 54628 29372 55468 29428
rect 55524 29372 55534 29428
rect 56690 29372 56700 29428
rect 56756 29372 56766 29428
rect 57558 29372 57596 29428
rect 57652 29372 57662 29428
rect 58034 29372 58044 29428
rect 58100 29372 60284 29428
rect 60340 29372 60350 29428
rect 60722 29372 60732 29428
rect 60788 29372 62412 29428
rect 62468 29372 62478 29428
rect 56700 29316 56756 29372
rect 3154 29260 3164 29316
rect 3220 29260 4620 29316
rect 4676 29260 6300 29316
rect 6356 29260 6972 29316
rect 7028 29260 7038 29316
rect 24658 29260 24668 29316
rect 24724 29260 27076 29316
rect 27346 29260 27356 29316
rect 27412 29260 28700 29316
rect 28756 29260 30156 29316
rect 30212 29260 30222 29316
rect 35074 29260 35084 29316
rect 35140 29260 35308 29316
rect 35634 29260 35644 29316
rect 35700 29260 35756 29316
rect 35812 29260 35822 29316
rect 36866 29260 36876 29316
rect 36932 29260 37044 29316
rect 40198 29260 40236 29316
rect 40292 29260 40302 29316
rect 43362 29260 43372 29316
rect 43428 29260 43596 29316
rect 43652 29260 43662 29316
rect 44706 29260 44716 29316
rect 44772 29260 45836 29316
rect 45892 29260 45902 29316
rect 46498 29260 46508 29316
rect 46564 29260 48748 29316
rect 48804 29260 51996 29316
rect 52052 29260 54908 29316
rect 54964 29260 54974 29316
rect 56700 29260 61180 29316
rect 61236 29260 61246 29316
rect 27020 29204 27076 29260
rect 3490 29148 3500 29204
rect 3556 29148 4508 29204
rect 4564 29148 6188 29204
rect 6244 29148 6254 29204
rect 9538 29148 9548 29204
rect 9604 29148 14476 29204
rect 14532 29148 16716 29204
rect 16772 29148 16782 29204
rect 19740 29148 22316 29204
rect 22372 29148 22382 29204
rect 26786 29148 26796 29204
rect 19740 29092 19796 29148
rect 26852 29092 26908 29204
rect 27020 29148 28476 29204
rect 28532 29148 33180 29204
rect 33236 29148 33246 29204
rect 35186 29148 35196 29204
rect 35252 29148 35868 29204
rect 35924 29148 35934 29204
rect 36988 29092 37044 29260
rect 37324 29148 38780 29204
rect 38836 29148 38846 29204
rect 42018 29148 42028 29204
rect 42084 29148 44156 29204
rect 44212 29148 44222 29204
rect 45266 29148 45276 29204
rect 45332 29148 46732 29204
rect 46788 29148 46798 29204
rect 47170 29148 47180 29204
rect 47236 29148 48972 29204
rect 49028 29148 49038 29204
rect 55794 29148 55804 29204
rect 55860 29148 56868 29204
rect 57250 29148 57260 29204
rect 57316 29148 58828 29204
rect 58884 29148 58894 29204
rect 13010 29036 13020 29092
rect 13076 29036 14364 29092
rect 14420 29036 14430 29092
rect 16146 29036 16156 29092
rect 16212 29036 19740 29092
rect 19796 29036 19806 29092
rect 22194 29036 22204 29092
rect 22260 29036 26124 29092
rect 26180 29036 29708 29092
rect 29764 29036 29774 29092
rect 36194 29036 36204 29092
rect 36260 29036 36270 29092
rect 36978 29036 36988 29092
rect 37044 29036 37054 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 36204 28980 36260 29036
rect 37324 28980 37380 29148
rect 56812 29092 56868 29148
rect 40114 29036 40124 29092
rect 40180 29036 42700 29092
rect 42756 29036 48636 29092
rect 48692 29036 48702 29092
rect 55458 29036 55468 29092
rect 55524 29036 56588 29092
rect 56644 29036 56654 29092
rect 56812 29036 60732 29092
rect 60788 29036 60798 29092
rect 63200 28980 64000 29008
rect 14130 28924 14140 28980
rect 14196 28924 15260 28980
rect 15316 28924 17276 28980
rect 17332 28924 17342 28980
rect 36204 28924 36372 28980
rect 36642 28924 36652 28980
rect 36708 28924 37380 28980
rect 46722 28924 46732 28980
rect 46788 28924 49756 28980
rect 49812 28924 52164 28980
rect 56242 28924 56252 28980
rect 56308 28924 56364 28980
rect 56420 28924 56430 28980
rect 59714 28924 59724 28980
rect 59780 28924 64000 28980
rect 36316 28868 36372 28924
rect 1698 28812 1708 28868
rect 1764 28812 2268 28868
rect 2324 28812 4396 28868
rect 4452 28812 5516 28868
rect 5572 28812 5582 28868
rect 12674 28812 12684 28868
rect 12740 28812 17052 28868
rect 17108 28812 17118 28868
rect 19506 28812 19516 28868
rect 19572 28812 20300 28868
rect 20356 28812 20524 28868
rect 20580 28812 20590 28868
rect 29922 28812 29932 28868
rect 29988 28812 31052 28868
rect 31108 28812 31118 28868
rect 32610 28812 32620 28868
rect 32676 28812 35196 28868
rect 35252 28812 35262 28868
rect 35858 28812 35868 28868
rect 35924 28812 37212 28868
rect 37268 28812 39004 28868
rect 39060 28812 39070 28868
rect 39890 28812 39900 28868
rect 39956 28812 40796 28868
rect 40852 28812 40862 28868
rect 45154 28812 45164 28868
rect 45220 28812 47236 28868
rect 48850 28812 48860 28868
rect 48916 28812 50540 28868
rect 50596 28812 50606 28868
rect 47180 28756 47236 28812
rect 52108 28756 52164 28924
rect 63200 28896 64000 28924
rect 53666 28812 53676 28868
rect 53732 28812 56588 28868
rect 56644 28812 56654 28868
rect 60050 28812 60060 28868
rect 60116 28812 60620 28868
rect 60676 28812 60686 28868
rect 1922 28700 1932 28756
rect 1988 28700 2380 28756
rect 2436 28700 2446 28756
rect 10546 28700 10556 28756
rect 10612 28700 13132 28756
rect 13188 28700 13198 28756
rect 14690 28700 14700 28756
rect 14756 28700 17388 28756
rect 17444 28700 17454 28756
rect 18610 28700 18620 28756
rect 18676 28700 19964 28756
rect 20020 28700 20030 28756
rect 24546 28700 24556 28756
rect 24612 28700 26236 28756
rect 26292 28700 26302 28756
rect 28354 28700 28364 28756
rect 28420 28700 29148 28756
rect 29204 28700 29214 28756
rect 30370 28700 30380 28756
rect 30436 28700 31444 28756
rect 32498 28700 32508 28756
rect 32564 28700 33852 28756
rect 33908 28700 33918 28756
rect 41234 28700 41244 28756
rect 41300 28700 43932 28756
rect 43988 28700 46956 28756
rect 47012 28700 47022 28756
rect 47180 28700 51772 28756
rect 51828 28700 51838 28756
rect 52098 28700 52108 28756
rect 52164 28700 55020 28756
rect 55076 28700 55086 28756
rect 56214 28700 56252 28756
rect 56308 28700 56318 28756
rect 31388 28644 31444 28700
rect 1810 28588 1820 28644
rect 1876 28588 5628 28644
rect 5684 28588 5694 28644
rect 7634 28588 7644 28644
rect 7700 28588 9436 28644
rect 9492 28588 10332 28644
rect 10388 28588 10398 28644
rect 12786 28588 12796 28644
rect 12852 28588 13468 28644
rect 13524 28588 13534 28644
rect 14354 28588 14364 28644
rect 14420 28588 16268 28644
rect 16324 28588 16334 28644
rect 19058 28588 19068 28644
rect 19124 28588 19628 28644
rect 19684 28588 19694 28644
rect 20850 28588 20860 28644
rect 20916 28588 26124 28644
rect 26180 28588 26190 28644
rect 29698 28588 29708 28644
rect 29764 28588 30492 28644
rect 30548 28588 31164 28644
rect 31220 28588 31230 28644
rect 31378 28588 31388 28644
rect 31444 28588 33292 28644
rect 33348 28588 33358 28644
rect 35186 28588 35196 28644
rect 35252 28588 35980 28644
rect 36036 28588 36988 28644
rect 37044 28588 37054 28644
rect 38518 28588 38556 28644
rect 38612 28588 38622 28644
rect 39666 28588 39676 28644
rect 39732 28588 41356 28644
rect 41412 28588 45948 28644
rect 46004 28588 46014 28644
rect 49858 28588 49868 28644
rect 49924 28588 50988 28644
rect 51044 28588 51054 28644
rect 53116 28588 54348 28644
rect 54404 28588 54414 28644
rect 56802 28588 56812 28644
rect 56868 28588 57932 28644
rect 57988 28588 57998 28644
rect 59826 28588 59836 28644
rect 59892 28588 61068 28644
rect 61124 28588 61628 28644
rect 61684 28588 61694 28644
rect 53116 28532 53172 28588
rect 17266 28476 17276 28532
rect 17332 28476 18060 28532
rect 18116 28476 20356 28532
rect 25666 28476 25676 28532
rect 25732 28476 37716 28532
rect 42018 28476 42028 28532
rect 42084 28476 42700 28532
rect 42756 28476 42766 28532
rect 48738 28476 48748 28532
rect 48804 28476 53172 28532
rect 55794 28476 55804 28532
rect 55860 28476 56476 28532
rect 56532 28476 58044 28532
rect 58100 28476 58110 28532
rect 58706 28476 58716 28532
rect 58772 28476 59276 28532
rect 59332 28476 61516 28532
rect 61572 28476 61582 28532
rect 2258 28364 2268 28420
rect 2324 28364 2604 28420
rect 2660 28364 2670 28420
rect 16594 28364 16604 28420
rect 16660 28364 18172 28420
rect 18228 28364 20244 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 20188 28196 20244 28364
rect 20300 28308 20356 28476
rect 28802 28364 28812 28420
rect 28868 28364 31164 28420
rect 31220 28364 31230 28420
rect 32386 28364 32396 28420
rect 32452 28364 34356 28420
rect 34626 28364 34636 28420
rect 34692 28364 34972 28420
rect 35028 28364 35038 28420
rect 36166 28364 36204 28420
rect 36260 28364 36270 28420
rect 34300 28308 34356 28364
rect 37660 28308 37716 28476
rect 39106 28364 39116 28420
rect 39172 28364 39788 28420
rect 39844 28364 39854 28420
rect 41234 28364 41244 28420
rect 41300 28364 52164 28420
rect 55234 28364 55244 28420
rect 55300 28364 57148 28420
rect 57204 28364 57214 28420
rect 61394 28364 61404 28420
rect 61460 28364 62188 28420
rect 62244 28364 62254 28420
rect 52108 28308 52164 28364
rect 63200 28308 64000 28336
rect 20300 28252 31500 28308
rect 31556 28252 31566 28308
rect 31938 28252 31948 28308
rect 32004 28252 32956 28308
rect 33012 28252 33022 28308
rect 34290 28252 34300 28308
rect 34356 28252 34748 28308
rect 34804 28252 34814 28308
rect 35522 28252 35532 28308
rect 35588 28252 35868 28308
rect 35924 28252 35934 28308
rect 36082 28252 36092 28308
rect 36148 28252 36428 28308
rect 36484 28252 36494 28308
rect 37650 28252 37660 28308
rect 37716 28252 37726 28308
rect 38434 28252 38444 28308
rect 38500 28252 39900 28308
rect 39956 28252 39966 28308
rect 41906 28252 41916 28308
rect 41972 28252 45164 28308
rect 45220 28252 45230 28308
rect 52098 28252 52108 28308
rect 52164 28252 53340 28308
rect 53396 28252 53406 28308
rect 56466 28252 56476 28308
rect 56532 28252 57036 28308
rect 57092 28252 57102 28308
rect 60274 28252 60284 28308
rect 60340 28252 64000 28308
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 63200 28224 64000 28252
rect 3378 28140 3388 28196
rect 3444 28140 4508 28196
rect 4564 28140 4574 28196
rect 20188 28140 38556 28196
rect 38612 28140 38622 28196
rect 40450 28140 40460 28196
rect 40516 28140 45948 28196
rect 46004 28140 47292 28196
rect 47348 28140 48300 28196
rect 48356 28140 48366 28196
rect 51986 28140 51996 28196
rect 52052 28140 52444 28196
rect 52500 28140 53004 28196
rect 53060 28140 53676 28196
rect 53732 28140 53742 28196
rect 53890 28140 53900 28196
rect 53956 28140 55580 28196
rect 55636 28140 55646 28196
rect 57698 28140 57708 28196
rect 57764 28140 61964 28196
rect 62020 28140 62030 28196
rect 1250 28028 1260 28084
rect 1316 28028 2940 28084
rect 2996 28028 5516 28084
rect 5572 28028 5582 28084
rect 6290 28028 6300 28084
rect 6356 28028 8428 28084
rect 8484 28028 8494 28084
rect 10546 28028 10556 28084
rect 10612 28028 11340 28084
rect 11396 28028 11564 28084
rect 11620 28028 12460 28084
rect 12516 28028 12526 28084
rect 18050 28028 18060 28084
rect 18116 28028 32788 28084
rect 33506 28028 33516 28084
rect 33572 28028 34076 28084
rect 34132 28028 34142 28084
rect 34300 28028 37380 28084
rect 37762 28028 37772 28084
rect 37828 28028 39228 28084
rect 39284 28028 39294 28084
rect 40002 28028 40012 28084
rect 40068 28028 40236 28084
rect 40292 28028 40302 28084
rect 41570 28028 41580 28084
rect 41636 28028 43148 28084
rect 43204 28028 43214 28084
rect 47170 28028 47180 28084
rect 47236 28028 55020 28084
rect 55076 28028 55086 28084
rect 56326 28028 56364 28084
rect 56420 28028 56430 28084
rect 32732 27972 32788 28028
rect 34300 27972 34356 28028
rect 1922 27916 1932 27972
rect 1988 27916 4060 27972
rect 4116 27916 4508 27972
rect 4564 27916 4574 27972
rect 10882 27916 10892 27972
rect 10948 27916 11676 27972
rect 11732 27916 12236 27972
rect 12292 27916 12302 27972
rect 13346 27916 13356 27972
rect 13412 27916 18620 27972
rect 18676 27916 18686 27972
rect 21074 27916 21084 27972
rect 21140 27916 21756 27972
rect 21812 27916 23436 27972
rect 23492 27916 23502 27972
rect 24658 27916 24668 27972
rect 24724 27916 26012 27972
rect 26068 27916 26078 27972
rect 26226 27916 26236 27972
rect 26292 27916 27468 27972
rect 27524 27916 28588 27972
rect 28644 27916 28654 27972
rect 32732 27916 34356 27972
rect 2258 27804 2268 27860
rect 2324 27804 3724 27860
rect 3780 27804 3790 27860
rect 3938 27804 3948 27860
rect 4004 27804 5628 27860
rect 5684 27804 5694 27860
rect 11302 27804 11340 27860
rect 11396 27804 11406 27860
rect 12338 27804 12348 27860
rect 12404 27804 13804 27860
rect 13860 27804 14588 27860
rect 14644 27804 14924 27860
rect 14980 27804 14990 27860
rect 19170 27804 19180 27860
rect 19236 27804 22764 27860
rect 22820 27804 22830 27860
rect 24210 27804 24220 27860
rect 24276 27804 25452 27860
rect 25508 27804 25518 27860
rect 26674 27804 26684 27860
rect 26740 27804 27580 27860
rect 27636 27804 27646 27860
rect 31714 27804 31724 27860
rect 31780 27804 33628 27860
rect 33684 27804 33694 27860
rect 35522 27804 35532 27860
rect 35588 27804 35756 27860
rect 35812 27804 36764 27860
rect 36820 27804 36830 27860
rect 37324 27748 37380 28028
rect 38668 27860 38724 28028
rect 38892 27916 40124 27972
rect 40180 27916 41468 27972
rect 41524 27916 41534 27972
rect 47506 27916 47516 27972
rect 47572 27916 50092 27972
rect 50148 27916 50158 27972
rect 50372 27916 52500 27972
rect 52658 27916 52668 27972
rect 52724 27916 53564 27972
rect 53620 27916 54796 27972
rect 54852 27916 54862 27972
rect 57586 27916 57596 27972
rect 57652 27916 58604 27972
rect 58660 27916 61292 27972
rect 61348 27916 61358 27972
rect 37538 27804 37548 27860
rect 37604 27804 38332 27860
rect 38388 27804 38398 27860
rect 38658 27804 38668 27860
rect 38724 27804 38734 27860
rect 38892 27748 38948 27916
rect 50372 27860 50428 27916
rect 52444 27860 52500 27916
rect 59724 27860 59780 27916
rect 9986 27692 9996 27748
rect 10052 27692 14700 27748
rect 14756 27692 14766 27748
rect 16706 27692 16716 27748
rect 16772 27692 18732 27748
rect 18788 27692 18798 27748
rect 24322 27692 24332 27748
rect 24388 27692 25676 27748
rect 25732 27692 26348 27748
rect 26404 27692 26414 27748
rect 31266 27692 31276 27748
rect 31332 27692 31500 27748
rect 31556 27692 31566 27748
rect 33730 27692 33740 27748
rect 33796 27692 34188 27748
rect 34244 27692 37100 27748
rect 37156 27692 37166 27748
rect 37324 27692 37492 27748
rect 38434 27692 38444 27748
rect 38500 27692 38948 27748
rect 39564 27804 46060 27860
rect 46116 27804 46732 27860
rect 46788 27804 46798 27860
rect 50194 27804 50204 27860
rect 50260 27804 50428 27860
rect 50754 27804 50764 27860
rect 50820 27804 51996 27860
rect 52052 27804 52062 27860
rect 52444 27804 54460 27860
rect 54516 27804 54526 27860
rect 59714 27804 59724 27860
rect 59780 27804 59790 27860
rect 1250 27580 1260 27636
rect 1316 27580 8092 27636
rect 8148 27580 8158 27636
rect 31490 27580 31500 27636
rect 31556 27580 37212 27636
rect 37268 27580 37278 27636
rect 6178 27468 6188 27524
rect 6244 27468 9548 27524
rect 9604 27468 23660 27524
rect 23716 27468 23726 27524
rect 35830 27468 35868 27524
rect 35924 27468 35934 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 37436 27412 37492 27692
rect 39564 27524 39620 27804
rect 39778 27692 39788 27748
rect 39844 27692 41692 27748
rect 41748 27692 41758 27748
rect 43148 27692 49980 27748
rect 50036 27692 51324 27748
rect 51380 27692 51390 27748
rect 52882 27692 52892 27748
rect 52948 27692 55356 27748
rect 55412 27692 55422 27748
rect 43148 27636 43204 27692
rect 63200 27636 64000 27664
rect 41570 27580 41580 27636
rect 41636 27580 43204 27636
rect 43810 27580 43820 27636
rect 43876 27580 46396 27636
rect 46452 27580 46462 27636
rect 51398 27580 51436 27636
rect 51492 27580 51502 27636
rect 52210 27580 52220 27636
rect 52276 27580 54684 27636
rect 54740 27580 54750 27636
rect 55458 27580 55468 27636
rect 55524 27580 62076 27636
rect 62132 27580 62142 27636
rect 62962 27580 62972 27636
rect 63028 27580 64000 27636
rect 63200 27552 64000 27580
rect 37650 27468 37660 27524
rect 37716 27468 39620 27524
rect 46498 27468 46508 27524
rect 46564 27468 50204 27524
rect 50260 27468 50270 27524
rect 54450 27468 54460 27524
rect 54516 27468 57596 27524
rect 57652 27468 57662 27524
rect 59714 27468 59724 27524
rect 59780 27468 60284 27524
rect 60340 27468 60350 27524
rect 10210 27356 10220 27412
rect 10276 27356 24444 27412
rect 24500 27356 24510 27412
rect 26114 27356 26124 27412
rect 26180 27356 26796 27412
rect 26852 27356 26862 27412
rect 31602 27356 31612 27412
rect 31668 27356 32508 27412
rect 32564 27356 33404 27412
rect 33460 27356 33470 27412
rect 37436 27356 39452 27412
rect 39508 27356 40348 27412
rect 40404 27356 41692 27412
rect 41748 27356 50876 27412
rect 50932 27356 57708 27412
rect 57764 27356 57774 27412
rect 9314 27244 9324 27300
rect 9380 27244 15148 27300
rect 15204 27244 15214 27300
rect 20514 27244 20524 27300
rect 20580 27244 23660 27300
rect 23716 27244 33908 27300
rect 34066 27244 34076 27300
rect 34132 27244 37772 27300
rect 37828 27244 37838 27300
rect 38322 27244 38332 27300
rect 38388 27244 40908 27300
rect 40964 27244 40974 27300
rect 45602 27244 45612 27300
rect 45668 27244 49756 27300
rect 49812 27244 49822 27300
rect 51650 27244 51660 27300
rect 51716 27244 55356 27300
rect 55412 27244 55422 27300
rect 55794 27244 55804 27300
rect 55860 27244 56812 27300
rect 56868 27244 58268 27300
rect 58324 27244 58334 27300
rect 33852 27188 33908 27244
rect 1922 27132 1932 27188
rect 1988 27132 2716 27188
rect 2772 27132 6188 27188
rect 6244 27132 6254 27188
rect 6738 27132 6748 27188
rect 6804 27132 7756 27188
rect 7812 27132 7822 27188
rect 8082 27132 8092 27188
rect 8148 27132 10220 27188
rect 10276 27132 10286 27188
rect 15092 27132 19068 27188
rect 19124 27132 19516 27188
rect 19572 27132 19582 27188
rect 25218 27132 25228 27188
rect 25284 27132 26572 27188
rect 26628 27132 26638 27188
rect 26786 27132 26796 27188
rect 26852 27132 26908 27188
rect 26964 27132 31948 27188
rect 32004 27132 33404 27188
rect 33460 27132 33470 27188
rect 33852 27132 34860 27188
rect 34916 27132 34926 27188
rect 39106 27132 39116 27188
rect 39172 27132 41132 27188
rect 41188 27132 41198 27188
rect 42690 27132 42700 27188
rect 42756 27132 43148 27188
rect 43204 27132 43214 27188
rect 50306 27132 50316 27188
rect 50372 27132 50540 27188
rect 50596 27132 50606 27188
rect 59042 27132 59052 27188
rect 59108 27132 59836 27188
rect 59892 27132 60620 27188
rect 60676 27132 61180 27188
rect 61236 27132 61246 27188
rect 61506 27132 61516 27188
rect 61572 27132 62188 27188
rect 62244 27132 62254 27188
rect 15092 27076 15148 27132
rect 4050 27020 4060 27076
rect 4116 27020 4620 27076
rect 4676 27020 4686 27076
rect 7830 27020 7868 27076
rect 7924 27020 7934 27076
rect 10994 27020 11004 27076
rect 11060 27020 14028 27076
rect 14084 27020 15148 27076
rect 18834 27020 18844 27076
rect 18900 27020 19292 27076
rect 19348 27020 19358 27076
rect 21186 27020 21196 27076
rect 21252 27020 22428 27076
rect 22484 27020 23324 27076
rect 23380 27020 23390 27076
rect 25330 27020 25340 27076
rect 25396 27020 26796 27076
rect 26852 27020 26862 27076
rect 35196 27020 35756 27076
rect 35812 27020 35822 27076
rect 37202 27020 37212 27076
rect 37268 27020 37660 27076
rect 37716 27020 37726 27076
rect 46134 27020 46172 27076
rect 46228 27020 46238 27076
rect 47282 27020 47292 27076
rect 47348 27020 48748 27076
rect 48804 27020 48814 27076
rect 50978 27020 50988 27076
rect 51044 27020 52556 27076
rect 52612 27020 52622 27076
rect 60162 27020 60172 27076
rect 60228 27020 61404 27076
rect 61460 27020 61470 27076
rect 35196 26964 35252 27020
rect 60172 26964 60228 27020
rect 4722 26908 4732 26964
rect 4788 26908 6972 26964
rect 7028 26908 7084 26964
rect 7140 26908 7150 26964
rect 8194 26908 8204 26964
rect 8260 26908 8988 26964
rect 9044 26908 10444 26964
rect 10500 26908 10510 26964
rect 10658 26908 10668 26964
rect 10724 26908 11900 26964
rect 11956 26908 12404 26964
rect 15026 26908 15036 26964
rect 15092 26908 16940 26964
rect 16996 26908 18732 26964
rect 18788 26908 18798 26964
rect 27122 26908 27132 26964
rect 27188 26908 27804 26964
rect 27860 26908 33964 26964
rect 34020 26908 34030 26964
rect 34514 26908 34524 26964
rect 34580 26908 35196 26964
rect 35252 26908 35262 26964
rect 35858 26908 35868 26964
rect 35924 26908 42812 26964
rect 42868 26908 42878 26964
rect 43474 26908 43484 26964
rect 43540 26908 43820 26964
rect 43876 26908 43886 26964
rect 44818 26908 44828 26964
rect 44884 26908 49756 26964
rect 49812 26908 49822 26964
rect 50082 26908 50092 26964
rect 50148 26908 55804 26964
rect 55860 26908 55870 26964
rect 56466 26908 56476 26964
rect 56532 26908 57036 26964
rect 57092 26908 60228 26964
rect 6710 26796 6748 26852
rect 6804 26796 6814 26852
rect 11442 26796 11452 26852
rect 11508 26796 11788 26852
rect 11844 26796 11854 26852
rect 12348 26740 12404 26908
rect 12562 26796 12572 26852
rect 12628 26796 13244 26852
rect 13300 26796 15484 26852
rect 15540 26796 15932 26852
rect 15988 26796 15998 26852
rect 26338 26796 26348 26852
rect 26404 26796 26684 26852
rect 26740 26796 27580 26852
rect 27636 26796 27646 26852
rect 30482 26796 30492 26852
rect 30548 26796 30828 26852
rect 30884 26796 30894 26852
rect 33058 26796 33068 26852
rect 33124 26796 36316 26852
rect 36372 26796 36382 26852
rect 37314 26796 37324 26852
rect 37380 26796 38220 26852
rect 38276 26796 38286 26852
rect 43334 26796 43372 26852
rect 43428 26796 43438 26852
rect 45612 26796 50428 26852
rect 51874 26796 51884 26852
rect 51940 26796 52780 26852
rect 52836 26796 52846 26852
rect 57138 26796 57148 26852
rect 57204 26796 58268 26852
rect 58324 26796 60172 26852
rect 60228 26796 61180 26852
rect 61236 26796 61246 26852
rect 45612 26740 45668 26796
rect 12348 26684 12908 26740
rect 12964 26684 12974 26740
rect 17042 26684 17052 26740
rect 17108 26684 17118 26740
rect 38546 26684 38556 26740
rect 38612 26684 44828 26740
rect 44884 26684 45668 26740
rect 17052 26628 17108 26684
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 11778 26572 11788 26628
rect 11844 26572 12460 26628
rect 12516 26572 12526 26628
rect 15474 26572 15484 26628
rect 15540 26572 17276 26628
rect 17332 26572 17342 26628
rect 29026 26572 29036 26628
rect 29092 26572 30604 26628
rect 30660 26572 40460 26628
rect 40516 26572 40526 26628
rect 42914 26572 42924 26628
rect 42980 26572 43820 26628
rect 43876 26572 45164 26628
rect 45220 26572 45230 26628
rect 6748 26460 8540 26516
rect 8596 26460 8606 26516
rect 12226 26460 12236 26516
rect 12292 26460 14588 26516
rect 14644 26460 15820 26516
rect 15876 26460 15886 26516
rect 17714 26460 17724 26516
rect 17780 26460 18396 26516
rect 18452 26460 18462 26516
rect 26226 26460 26236 26516
rect 26292 26460 29148 26516
rect 29204 26460 29214 26516
rect 38612 26460 46508 26516
rect 46564 26460 46574 26516
rect 47058 26460 47068 26516
rect 47124 26460 48188 26516
rect 48244 26460 48254 26516
rect 6748 26404 6804 26460
rect 38612 26404 38668 26460
rect 2146 26348 2156 26404
rect 2212 26348 3500 26404
rect 3556 26348 3566 26404
rect 5618 26348 5628 26404
rect 5684 26348 6804 26404
rect 9986 26348 9996 26404
rect 10052 26348 22764 26404
rect 22820 26348 22830 26404
rect 23286 26348 23324 26404
rect 23380 26348 23390 26404
rect 28354 26348 28364 26404
rect 28420 26348 38668 26404
rect 39666 26348 39676 26404
rect 39732 26348 40012 26404
rect 40068 26348 40078 26404
rect 46050 26348 46060 26404
rect 46116 26348 50092 26404
rect 50148 26348 50158 26404
rect 6748 26292 6804 26348
rect 4834 26236 4844 26292
rect 4900 26236 5964 26292
rect 6020 26236 6030 26292
rect 6738 26236 6748 26292
rect 6804 26236 6814 26292
rect 7746 26236 7756 26292
rect 7812 26236 8540 26292
rect 8596 26236 8606 26292
rect 12646 26236 12684 26292
rect 12740 26236 12750 26292
rect 13794 26236 13804 26292
rect 13860 26236 14812 26292
rect 14868 26236 15820 26292
rect 15876 26236 17612 26292
rect 17668 26236 17678 26292
rect 22194 26236 22204 26292
rect 22260 26236 24220 26292
rect 24276 26236 24286 26292
rect 26114 26236 26124 26292
rect 26180 26236 27916 26292
rect 27972 26236 27982 26292
rect 31154 26236 31164 26292
rect 31220 26236 34524 26292
rect 34580 26236 34590 26292
rect 38994 26236 39004 26292
rect 39060 26236 39452 26292
rect 39508 26236 40124 26292
rect 40180 26236 40190 26292
rect 42242 26236 42252 26292
rect 42308 26236 43708 26292
rect 43764 26236 45276 26292
rect 45332 26236 45342 26292
rect 45612 26236 49644 26292
rect 49700 26236 49710 26292
rect 45612 26180 45668 26236
rect 50372 26180 50428 26796
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 55570 26572 55580 26628
rect 55636 26572 56700 26628
rect 56756 26572 61740 26628
rect 61796 26572 61806 26628
rect 57474 26460 57484 26516
rect 57540 26460 61628 26516
rect 61684 26460 61694 26516
rect 54338 26348 54348 26404
rect 54404 26348 54684 26404
rect 54740 26348 54750 26404
rect 55794 26348 55804 26404
rect 55860 26348 56140 26404
rect 56196 26348 56206 26404
rect 57250 26348 57260 26404
rect 57316 26348 58604 26404
rect 58660 26348 58670 26404
rect 60386 26348 60396 26404
rect 60452 26348 62188 26404
rect 62244 26348 62254 26404
rect 60396 26292 60452 26348
rect 55122 26236 55132 26292
rect 55188 26236 56028 26292
rect 56084 26236 56094 26292
rect 57362 26236 57372 26292
rect 57428 26236 60452 26292
rect 4274 26124 4284 26180
rect 4340 26124 5516 26180
rect 5572 26124 5852 26180
rect 5908 26124 5918 26180
rect 6402 26124 6412 26180
rect 6468 26124 8428 26180
rect 8484 26124 8494 26180
rect 12786 26124 12796 26180
rect 12852 26124 15596 26180
rect 15652 26124 15662 26180
rect 17042 26124 17052 26180
rect 17108 26124 23772 26180
rect 23828 26124 24892 26180
rect 24948 26124 24958 26180
rect 31378 26124 31388 26180
rect 31444 26124 32172 26180
rect 32228 26124 34748 26180
rect 34804 26124 34814 26180
rect 41682 26124 41692 26180
rect 41748 26124 45612 26180
rect 45668 26124 45678 26180
rect 47618 26124 47628 26180
rect 47684 26124 48748 26180
rect 48804 26124 48814 26180
rect 50372 26124 62188 26180
rect 4284 26012 7028 26068
rect 13458 26012 13468 26068
rect 13524 26012 16492 26068
rect 16548 26012 17612 26068
rect 17668 26012 17678 26068
rect 18508 26012 22876 26068
rect 22932 26012 22942 26068
rect 25890 26012 25900 26068
rect 25956 26012 29148 26068
rect 29204 26012 29214 26068
rect 30482 26012 30492 26068
rect 30548 26012 44044 26068
rect 44100 26012 45500 26068
rect 45556 26012 45566 26068
rect 46610 26012 46620 26068
rect 46676 26012 52220 26068
rect 52276 26012 52286 26068
rect 56018 26012 56028 26068
rect 56084 26012 58044 26068
rect 58100 26012 58110 26068
rect 4284 25956 4340 26012
rect 6972 25956 7028 26012
rect 18508 25956 18564 26012
rect 62132 25956 62188 26124
rect 4274 25900 4284 25956
rect 4340 25900 4350 25956
rect 6972 25900 18564 25956
rect 18722 25900 18732 25956
rect 18788 25900 19404 25956
rect 19460 25900 19470 25956
rect 24658 25900 24668 25956
rect 24724 25900 26124 25956
rect 26180 25900 26190 25956
rect 32386 25900 32396 25956
rect 32452 25900 32956 25956
rect 33012 25900 33022 25956
rect 37762 25900 37772 25956
rect 37828 25900 38108 25956
rect 38164 25900 38174 25956
rect 42812 25900 47740 25956
rect 47796 25900 57708 25956
rect 57764 25900 57774 25956
rect 62132 25900 62524 25956
rect 62580 25900 62590 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 10322 25788 10332 25844
rect 10388 25788 15484 25844
rect 15540 25788 15550 25844
rect 15708 25788 21644 25844
rect 21700 25788 21710 25844
rect 26852 25788 34076 25844
rect 34132 25788 34142 25844
rect 15708 25732 15764 25788
rect 26852 25732 26908 25788
rect 42812 25732 42868 25900
rect 45378 25788 45388 25844
rect 45444 25788 46396 25844
rect 46452 25788 49868 25844
rect 49924 25788 49934 25844
rect 50306 25788 50316 25844
rect 50372 25788 50540 25844
rect 50596 25788 50606 25844
rect 54226 25788 54236 25844
rect 54292 25788 56028 25844
rect 56084 25788 56094 25844
rect 56914 25788 56924 25844
rect 56980 25788 58492 25844
rect 58548 25788 59724 25844
rect 59780 25788 59790 25844
rect 2930 25676 2940 25732
rect 2996 25676 5740 25732
rect 5796 25676 5806 25732
rect 12002 25676 12012 25732
rect 12068 25676 15764 25732
rect 17938 25676 17948 25732
rect 18004 25676 18956 25732
rect 19012 25676 19022 25732
rect 19618 25676 19628 25732
rect 19684 25676 20300 25732
rect 20356 25676 20366 25732
rect 20524 25676 26908 25732
rect 28466 25676 28476 25732
rect 28532 25676 30492 25732
rect 30548 25676 30558 25732
rect 38098 25676 38108 25732
rect 38164 25676 38668 25732
rect 42578 25676 42588 25732
rect 42644 25676 42812 25732
rect 42868 25676 42878 25732
rect 45042 25676 45052 25732
rect 45108 25676 46060 25732
rect 46116 25676 46126 25732
rect 49420 25676 50988 25732
rect 51044 25676 53788 25732
rect 53844 25676 53854 25732
rect 54898 25676 54908 25732
rect 54964 25676 56476 25732
rect 56532 25676 56542 25732
rect 4274 25564 4284 25620
rect 4340 25564 4396 25620
rect 4452 25564 4462 25620
rect 4946 25564 4956 25620
rect 5012 25564 9660 25620
rect 9716 25564 9726 25620
rect 16034 25564 16044 25620
rect 16100 25564 17724 25620
rect 17780 25564 18508 25620
rect 18564 25564 18574 25620
rect 20524 25508 20580 25676
rect 38612 25620 38668 25676
rect 20738 25564 20748 25620
rect 20804 25564 22092 25620
rect 22148 25564 22158 25620
rect 22306 25564 22316 25620
rect 22372 25564 24556 25620
rect 24612 25564 24622 25620
rect 34290 25564 34300 25620
rect 34356 25564 35084 25620
rect 35140 25564 35150 25620
rect 38210 25564 38220 25620
rect 38276 25564 38286 25620
rect 38612 25564 40684 25620
rect 40740 25564 41356 25620
rect 41412 25564 41422 25620
rect 45154 25564 45164 25620
rect 45220 25564 47068 25620
rect 47124 25564 47134 25620
rect 38220 25508 38276 25564
rect 49420 25508 49476 25676
rect 55122 25564 55132 25620
rect 55188 25564 55692 25620
rect 55748 25564 55758 25620
rect 3490 25452 3500 25508
rect 3556 25452 6748 25508
rect 6804 25452 6814 25508
rect 12562 25452 12572 25508
rect 12628 25452 13020 25508
rect 13076 25452 13086 25508
rect 15138 25452 15148 25508
rect 15204 25452 17052 25508
rect 17108 25452 17118 25508
rect 18358 25452 18396 25508
rect 18452 25452 20580 25508
rect 20850 25452 20860 25508
rect 20916 25452 21868 25508
rect 21924 25452 21934 25508
rect 22530 25452 22540 25508
rect 22596 25452 26236 25508
rect 26292 25452 26302 25508
rect 35410 25452 35420 25508
rect 35476 25452 35756 25508
rect 35812 25452 36988 25508
rect 37044 25452 37054 25508
rect 38220 25452 38668 25508
rect 40114 25452 40124 25508
rect 40180 25452 41692 25508
rect 41748 25452 42588 25508
rect 42644 25452 42654 25508
rect 44230 25452 44268 25508
rect 44324 25452 47964 25508
rect 48020 25452 48030 25508
rect 48962 25452 48972 25508
rect 49028 25452 49420 25508
rect 49476 25452 49486 25508
rect 50082 25452 50092 25508
rect 50148 25452 50876 25508
rect 50932 25452 50942 25508
rect 52770 25452 52780 25508
rect 52836 25452 55188 25508
rect 38612 25396 38668 25452
rect 55132 25396 55188 25452
rect 2370 25340 2380 25396
rect 2436 25340 4284 25396
rect 4340 25340 4350 25396
rect 10770 25340 10780 25396
rect 10836 25340 13132 25396
rect 13188 25340 13198 25396
rect 18022 25340 18060 25396
rect 18116 25340 18126 25396
rect 19506 25340 19516 25396
rect 19572 25340 21532 25396
rect 21588 25340 21598 25396
rect 22194 25340 22204 25396
rect 22260 25340 22270 25396
rect 23202 25340 23212 25396
rect 23268 25340 29484 25396
rect 29540 25340 29550 25396
rect 30818 25340 30828 25396
rect 30884 25340 35084 25396
rect 35140 25340 35150 25396
rect 38612 25340 39116 25396
rect 39172 25340 39182 25396
rect 46162 25340 46172 25396
rect 46228 25340 47068 25396
rect 47124 25340 47134 25396
rect 49298 25340 49308 25396
rect 49364 25340 50540 25396
rect 50596 25340 50606 25396
rect 51314 25340 51324 25396
rect 51380 25340 52892 25396
rect 52948 25340 52958 25396
rect 55122 25340 55132 25396
rect 55188 25340 60620 25396
rect 60676 25340 60686 25396
rect 22204 25284 22260 25340
rect 5282 25228 5292 25284
rect 5348 25228 5852 25284
rect 5908 25228 5918 25284
rect 6962 25228 6972 25284
rect 7028 25228 7756 25284
rect 7812 25228 7822 25284
rect 8418 25228 8428 25284
rect 8484 25228 11004 25284
rect 11060 25228 11070 25284
rect 11974 25228 12012 25284
rect 12068 25228 12078 25284
rect 12422 25228 12460 25284
rect 12516 25228 12526 25284
rect 13570 25228 13580 25284
rect 13636 25228 14476 25284
rect 14532 25228 14542 25284
rect 18620 25228 22260 25284
rect 22754 25228 22764 25284
rect 22820 25228 22876 25284
rect 22932 25228 22942 25284
rect 24546 25228 24556 25284
rect 24612 25228 28140 25284
rect 28196 25228 29820 25284
rect 29876 25228 29886 25284
rect 30034 25228 30044 25284
rect 30100 25228 34412 25284
rect 34468 25228 35756 25284
rect 35812 25228 35822 25284
rect 38882 25228 38892 25284
rect 38948 25228 41020 25284
rect 41076 25228 41086 25284
rect 43586 25228 43596 25284
rect 43652 25228 44940 25284
rect 44996 25228 45006 25284
rect 45490 25228 45500 25284
rect 45556 25228 46620 25284
rect 46676 25228 46686 25284
rect 48626 25228 48636 25284
rect 48692 25228 49756 25284
rect 49812 25228 49822 25284
rect 53666 25228 53676 25284
rect 53732 25228 56812 25284
rect 56868 25228 57260 25284
rect 57316 25228 57326 25284
rect 5954 25116 5964 25172
rect 6020 25116 9436 25172
rect 9492 25116 9502 25172
rect 16818 25116 16828 25172
rect 16884 25116 18060 25172
rect 18116 25116 18396 25172
rect 18452 25116 18462 25172
rect 18620 25060 18676 25228
rect 26674 25116 26684 25172
rect 26740 25116 30828 25172
rect 30884 25116 30894 25172
rect 31266 25116 31276 25172
rect 31332 25116 32732 25172
rect 32788 25116 44604 25172
rect 44660 25116 44670 25172
rect 53778 25116 53788 25172
rect 53844 25116 59276 25172
rect 59332 25116 59342 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 2594 25004 2604 25060
rect 2660 25004 3836 25060
rect 3892 25004 3902 25060
rect 5842 25004 5852 25060
rect 5908 25004 8876 25060
rect 8932 25004 8942 25060
rect 12898 25004 12908 25060
rect 12964 25004 13580 25060
rect 13636 25004 13646 25060
rect 15026 25004 15036 25060
rect 15092 25004 18676 25060
rect 28130 25004 28140 25060
rect 28196 25004 31164 25060
rect 31220 25004 31230 25060
rect 41906 25004 41916 25060
rect 41972 25004 43148 25060
rect 43204 25004 43214 25060
rect 50166 25004 50204 25060
rect 50260 25004 50270 25060
rect 54002 25004 54012 25060
rect 54068 25004 57260 25060
rect 57316 25004 57326 25060
rect 0 24948 800 24976
rect 0 24892 1708 24948
rect 1764 24892 1774 24948
rect 2482 24892 2492 24948
rect 2548 24892 3388 24948
rect 12674 24892 12684 24948
rect 12740 24892 13132 24948
rect 13188 24892 13198 24948
rect 13346 24892 13356 24948
rect 13412 24892 13692 24948
rect 13748 24892 13758 24948
rect 14690 24892 14700 24948
rect 14756 24892 16604 24948
rect 16660 24892 16670 24948
rect 18834 24892 18844 24948
rect 18900 24892 19404 24948
rect 19460 24892 19470 24948
rect 25442 24892 25452 24948
rect 25508 24892 25900 24948
rect 25956 24892 25966 24948
rect 30566 24892 30604 24948
rect 30660 24892 31388 24948
rect 31444 24892 31454 24948
rect 34738 24892 34748 24948
rect 34804 24892 41020 24948
rect 41076 24892 41086 24948
rect 47954 24892 47964 24948
rect 48020 24892 50428 24948
rect 50530 24892 50540 24948
rect 50596 24892 51436 24948
rect 51492 24892 51502 24948
rect 57026 24892 57036 24948
rect 57092 24892 58604 24948
rect 58660 24892 58670 24948
rect 0 24864 800 24892
rect 3332 24836 3388 24892
rect 50372 24836 50428 24892
rect 3332 24780 4060 24836
rect 4116 24780 4732 24836
rect 4788 24780 5628 24836
rect 5684 24780 5694 24836
rect 6738 24780 6748 24836
rect 6804 24780 7420 24836
rect 7476 24780 7486 24836
rect 12338 24780 12348 24836
rect 12404 24780 13468 24836
rect 13524 24780 13534 24836
rect 14242 24780 14252 24836
rect 14308 24780 22876 24836
rect 22932 24780 22942 24836
rect 25666 24780 25676 24836
rect 25732 24780 31836 24836
rect 31892 24780 31902 24836
rect 32050 24780 32060 24836
rect 32116 24780 33404 24836
rect 33460 24780 33470 24836
rect 47618 24780 47628 24836
rect 47684 24780 49868 24836
rect 49924 24780 49934 24836
rect 50082 24780 50092 24836
rect 50148 24780 50186 24836
rect 50372 24780 56980 24836
rect 57138 24780 57148 24836
rect 57204 24780 57820 24836
rect 57876 24780 57886 24836
rect 56924 24724 56980 24780
rect 3490 24668 3500 24724
rect 3556 24668 5852 24724
rect 5908 24668 5918 24724
rect 7522 24668 7532 24724
rect 7588 24668 7980 24724
rect 8036 24668 8046 24724
rect 13346 24668 13356 24724
rect 13412 24668 16828 24724
rect 16884 24668 16894 24724
rect 17266 24668 17276 24724
rect 17332 24668 17500 24724
rect 17556 24668 18396 24724
rect 18452 24668 18462 24724
rect 19954 24668 19964 24724
rect 20020 24668 20972 24724
rect 21028 24668 21038 24724
rect 21298 24668 21308 24724
rect 21364 24668 23660 24724
rect 23716 24668 23726 24724
rect 31378 24668 31388 24724
rect 31444 24668 31500 24724
rect 31556 24668 31566 24724
rect 31724 24668 35532 24724
rect 35588 24668 35598 24724
rect 36642 24668 36652 24724
rect 36708 24668 38668 24724
rect 38724 24668 38734 24724
rect 44258 24668 44268 24724
rect 44324 24668 45052 24724
rect 45108 24668 45388 24724
rect 45444 24668 46396 24724
rect 46452 24668 46462 24724
rect 49522 24668 49532 24724
rect 49588 24668 49598 24724
rect 49746 24668 49756 24724
rect 49812 24668 51996 24724
rect 52052 24668 52062 24724
rect 52994 24668 53004 24724
rect 53060 24668 54684 24724
rect 54740 24668 54750 24724
rect 56924 24668 58156 24724
rect 58212 24668 58222 24724
rect 1362 24556 1372 24612
rect 1428 24556 8204 24612
rect 8260 24556 10164 24612
rect 10322 24556 10332 24612
rect 10388 24556 11788 24612
rect 11844 24556 11854 24612
rect 16594 24556 16604 24612
rect 16660 24556 21084 24612
rect 21140 24556 21150 24612
rect 10108 24500 10164 24556
rect 21308 24500 21364 24668
rect 24322 24556 24332 24612
rect 24388 24556 25676 24612
rect 25732 24556 25742 24612
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 2930 24444 2940 24500
rect 2996 24444 3388 24500
rect 6738 24444 6748 24500
rect 6804 24444 9548 24500
rect 9604 24444 9614 24500
rect 10108 24444 11900 24500
rect 11956 24444 11966 24500
rect 15586 24444 15596 24500
rect 15652 24444 21364 24500
rect 23650 24444 23660 24500
rect 23716 24444 24108 24500
rect 24164 24444 24174 24500
rect 25890 24444 25900 24500
rect 25956 24444 27132 24500
rect 27188 24444 27198 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 0 24220 1988 24276
rect 3332 24276 3388 24444
rect 31724 24388 31780 24668
rect 49532 24612 49588 24668
rect 31938 24556 31948 24612
rect 32004 24556 48860 24612
rect 48916 24556 48926 24612
rect 49532 24556 51884 24612
rect 51940 24556 51950 24612
rect 53330 24556 53340 24612
rect 53396 24556 53788 24612
rect 53844 24556 53854 24612
rect 33506 24444 33516 24500
rect 33572 24444 50540 24500
rect 50596 24444 50606 24500
rect 50978 24444 50988 24500
rect 51044 24444 52892 24500
rect 52948 24444 52958 24500
rect 56914 24444 56924 24500
rect 56980 24444 59500 24500
rect 59556 24444 60956 24500
rect 61012 24444 61022 24500
rect 8866 24332 8876 24388
rect 8932 24332 19292 24388
rect 19348 24332 19628 24388
rect 19684 24332 19694 24388
rect 20962 24332 20972 24388
rect 21028 24332 31780 24388
rect 36530 24332 36540 24388
rect 36596 24332 45444 24388
rect 50978 24332 50988 24388
rect 51044 24332 61852 24388
rect 61908 24332 61918 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 45388 24276 45444 24332
rect 3332 24220 3836 24276
rect 3892 24220 3902 24276
rect 6626 24220 6636 24276
rect 6692 24220 7196 24276
rect 7252 24220 7262 24276
rect 10882 24220 10892 24276
rect 10948 24220 28476 24276
rect 28532 24220 28542 24276
rect 30370 24220 30380 24276
rect 30436 24220 30446 24276
rect 39666 24220 39676 24276
rect 39732 24220 44156 24276
rect 44212 24220 44222 24276
rect 45378 24220 45388 24276
rect 45444 24220 45454 24276
rect 50306 24220 50316 24276
rect 50372 24220 50652 24276
rect 50708 24220 51548 24276
rect 51604 24220 51614 24276
rect 54786 24220 54796 24276
rect 54852 24220 55692 24276
rect 55748 24220 56588 24276
rect 56644 24220 56924 24276
rect 56980 24220 56990 24276
rect 0 24192 800 24220
rect 6962 24108 6972 24164
rect 7028 24108 7644 24164
rect 7700 24108 7710 24164
rect 8082 24108 8092 24164
rect 8148 24108 8764 24164
rect 8820 24108 8830 24164
rect 12226 24108 12236 24164
rect 12292 24108 12460 24164
rect 12516 24108 12526 24164
rect 13682 24108 13692 24164
rect 13748 24108 14700 24164
rect 14756 24108 14766 24164
rect 17686 24108 17724 24164
rect 17780 24108 17790 24164
rect 18946 24108 18956 24164
rect 19012 24108 19180 24164
rect 19236 24108 19628 24164
rect 19684 24108 19694 24164
rect 22978 24108 22988 24164
rect 23044 24108 24668 24164
rect 24724 24108 26348 24164
rect 26404 24108 26414 24164
rect 30380 24052 30436 24220
rect 32162 24108 32172 24164
rect 32228 24108 32238 24164
rect 34290 24108 34300 24164
rect 34356 24108 35084 24164
rect 35140 24108 35150 24164
rect 37314 24108 37324 24164
rect 37380 24108 38108 24164
rect 38164 24108 38174 24164
rect 40338 24108 40348 24164
rect 40404 24108 42924 24164
rect 42980 24108 42990 24164
rect 44370 24108 44380 24164
rect 44436 24108 46732 24164
rect 46788 24108 46798 24164
rect 50530 24108 50540 24164
rect 50596 24108 52668 24164
rect 52724 24108 52734 24164
rect 60050 24108 60060 24164
rect 60116 24108 60956 24164
rect 61012 24108 61516 24164
rect 61572 24108 61582 24164
rect 5058 23996 5068 24052
rect 5124 23996 10108 24052
rect 10164 23996 10174 24052
rect 19394 23996 19404 24052
rect 19460 23996 20188 24052
rect 20244 23996 20254 24052
rect 22418 23996 22428 24052
rect 22484 23996 23100 24052
rect 23156 23996 23166 24052
rect 23314 23996 23324 24052
rect 23380 23996 23418 24052
rect 23650 23996 23660 24052
rect 23716 23996 24332 24052
rect 24388 23996 24398 24052
rect 26786 23996 26796 24052
rect 26852 23996 30436 24052
rect 32172 24052 32228 24108
rect 32172 23996 49644 24052
rect 49700 23996 49710 24052
rect 50082 23996 50092 24052
rect 50148 23996 51436 24052
rect 51492 23996 52780 24052
rect 52836 23996 52846 24052
rect 57138 23996 57148 24052
rect 57204 23996 58156 24052
rect 58212 23996 58222 24052
rect 2594 23884 2604 23940
rect 2660 23884 4060 23940
rect 4116 23884 4126 23940
rect 5068 23828 5124 23996
rect 6710 23884 6748 23940
rect 6804 23884 6814 23940
rect 7046 23884 7084 23940
rect 7140 23884 7150 23940
rect 18722 23884 18732 23940
rect 18788 23884 20076 23940
rect 20132 23884 24444 23940
rect 24500 23884 24510 23940
rect 28140 23884 29372 23940
rect 29428 23884 29438 23940
rect 31602 23884 31612 23940
rect 31668 23884 32284 23940
rect 32340 23884 32350 23940
rect 33478 23884 33516 23940
rect 33572 23884 35756 23940
rect 35812 23884 37324 23940
rect 37380 23884 38668 23940
rect 40002 23884 40012 23940
rect 40068 23884 41580 23940
rect 41636 23884 41646 23940
rect 46722 23884 46732 23940
rect 46788 23884 47964 23940
rect 48020 23884 50204 23940
rect 50260 23884 51100 23940
rect 51156 23884 51166 23940
rect 54786 23884 54796 23940
rect 54852 23884 55468 23940
rect 55524 23884 55534 23940
rect 1474 23772 1484 23828
rect 1540 23772 5124 23828
rect 18834 23772 18844 23828
rect 18900 23772 19180 23828
rect 19236 23772 19964 23828
rect 20020 23772 21420 23828
rect 21476 23772 21486 23828
rect 22866 23772 22876 23828
rect 22932 23772 23212 23828
rect 23268 23772 23278 23828
rect 23538 23772 23548 23828
rect 23604 23772 24892 23828
rect 24948 23772 25116 23828
rect 25172 23772 25788 23828
rect 25844 23772 25854 23828
rect 26226 23772 26236 23828
rect 26292 23772 27356 23828
rect 27412 23772 27916 23828
rect 27972 23772 27982 23828
rect 914 23660 924 23716
rect 980 23660 9212 23716
rect 9268 23660 9436 23716
rect 9492 23660 9502 23716
rect 14130 23660 14140 23716
rect 14196 23660 16492 23716
rect 16548 23660 16558 23716
rect 16706 23660 16716 23716
rect 16772 23660 20524 23716
rect 20580 23660 20590 23716
rect 21522 23660 21532 23716
rect 21588 23660 21868 23716
rect 21924 23660 21934 23716
rect 23100 23660 23324 23716
rect 23380 23660 24108 23716
rect 24164 23660 24174 23716
rect 23100 23604 23156 23660
rect 3686 23548 3724 23604
rect 3780 23548 3790 23604
rect 5506 23548 5516 23604
rect 5572 23548 5852 23604
rect 5908 23548 5918 23604
rect 11778 23548 11788 23604
rect 11844 23548 18956 23604
rect 19012 23548 19022 23604
rect 21970 23548 21980 23604
rect 22036 23548 23100 23604
rect 23156 23548 23166 23604
rect 23874 23548 23884 23604
rect 23940 23548 26124 23604
rect 26180 23548 26190 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 28140 23492 28196 23884
rect 38612 23716 38668 23884
rect 41794 23772 41804 23828
rect 41860 23772 43596 23828
rect 43652 23772 43662 23828
rect 48850 23772 48860 23828
rect 48916 23772 49420 23828
rect 49476 23772 49486 23828
rect 49634 23772 49644 23828
rect 49700 23772 50876 23828
rect 50932 23772 51996 23828
rect 52052 23772 52062 23828
rect 57026 23772 57036 23828
rect 57092 23772 60620 23828
rect 60676 23772 60686 23828
rect 28578 23660 28588 23716
rect 28644 23660 30044 23716
rect 30100 23660 30604 23716
rect 30660 23660 30670 23716
rect 30818 23660 30828 23716
rect 30884 23660 34860 23716
rect 34916 23660 34926 23716
rect 35074 23660 35084 23716
rect 35140 23660 36092 23716
rect 36148 23660 36988 23716
rect 37044 23660 37054 23716
rect 38612 23660 39900 23716
rect 39956 23660 39966 23716
rect 40226 23660 40236 23716
rect 40292 23660 41692 23716
rect 41748 23660 41758 23716
rect 46834 23660 46844 23716
rect 46900 23660 50092 23716
rect 50148 23660 50158 23716
rect 50418 23660 50428 23716
rect 50484 23660 51100 23716
rect 51156 23660 51166 23716
rect 51314 23660 51324 23716
rect 51380 23660 53788 23716
rect 53844 23660 53854 23716
rect 54226 23660 54236 23716
rect 54292 23660 56364 23716
rect 56420 23660 56430 23716
rect 30828 23604 30884 23660
rect 30482 23548 30492 23604
rect 30548 23548 30884 23604
rect 31378 23548 31388 23604
rect 31444 23548 33404 23604
rect 33460 23548 33470 23604
rect 38630 23548 38668 23604
rect 38724 23548 38734 23604
rect 41570 23548 41580 23604
rect 41636 23548 42476 23604
rect 42532 23548 45052 23604
rect 45108 23548 45118 23604
rect 45378 23548 45388 23604
rect 45444 23548 46172 23604
rect 46228 23548 46238 23604
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 6626 23436 6636 23492
rect 6692 23436 7868 23492
rect 7924 23436 10220 23492
rect 10276 23436 10286 23492
rect 11890 23436 11900 23492
rect 11956 23436 13580 23492
rect 13636 23436 13646 23492
rect 13906 23436 13916 23492
rect 13972 23436 14812 23492
rect 14868 23436 14878 23492
rect 17378 23436 17388 23492
rect 17444 23436 19180 23492
rect 19236 23436 19246 23492
rect 23314 23436 23324 23492
rect 23380 23436 28196 23492
rect 36978 23436 36988 23492
rect 37044 23436 37436 23492
rect 37492 23436 39004 23492
rect 39060 23436 39070 23492
rect 39778 23436 39788 23492
rect 39844 23436 41804 23492
rect 41860 23436 43036 23492
rect 43092 23436 43102 23492
rect 46610 23436 46620 23492
rect 46676 23436 47404 23492
rect 47460 23436 47470 23492
rect 53442 23436 53452 23492
rect 53508 23436 56588 23492
rect 56644 23436 56654 23492
rect 57250 23436 57260 23492
rect 57316 23436 58716 23492
rect 58772 23436 58782 23492
rect 2034 23324 2044 23380
rect 2100 23324 7420 23380
rect 7476 23324 7486 23380
rect 9762 23324 9772 23380
rect 9828 23324 16716 23380
rect 16772 23324 16782 23380
rect 17826 23324 17836 23380
rect 17892 23324 19628 23380
rect 19684 23324 19694 23380
rect 24070 23324 24108 23380
rect 24164 23324 24174 23380
rect 24742 23324 24780 23380
rect 24836 23324 24846 23380
rect 29922 23324 29932 23380
rect 29988 23324 30268 23380
rect 30324 23324 31052 23380
rect 31108 23324 31118 23380
rect 36642 23324 36652 23380
rect 36708 23324 36718 23380
rect 38210 23324 38220 23380
rect 38276 23324 39620 23380
rect 40114 23324 40124 23380
rect 40180 23324 41132 23380
rect 41188 23324 41692 23380
rect 41748 23324 41758 23380
rect 43922 23324 43932 23380
rect 43988 23324 47516 23380
rect 47572 23324 47582 23380
rect 51986 23324 51996 23380
rect 52052 23324 54348 23380
rect 54404 23324 54414 23380
rect 36652 23268 36708 23324
rect 4050 23212 4060 23268
rect 4116 23212 8764 23268
rect 8820 23212 8830 23268
rect 14018 23212 14028 23268
rect 14084 23212 14588 23268
rect 14644 23212 14654 23268
rect 18050 23212 18060 23268
rect 18116 23212 23268 23268
rect 26450 23212 26460 23268
rect 26516 23212 27580 23268
rect 27636 23212 27916 23268
rect 27972 23212 29372 23268
rect 29428 23212 29438 23268
rect 33170 23212 33180 23268
rect 33236 23212 33852 23268
rect 33908 23212 34188 23268
rect 34244 23212 35868 23268
rect 35924 23212 35934 23268
rect 36652 23212 36988 23268
rect 37044 23212 37054 23268
rect 23212 23156 23268 23212
rect 39564 23156 39620 23324
rect 42018 23212 42028 23268
rect 42084 23212 44604 23268
rect 44660 23212 45612 23268
rect 45668 23212 45678 23268
rect 45938 23212 45948 23268
rect 46004 23212 47180 23268
rect 47236 23212 47246 23268
rect 52994 23212 53004 23268
rect 53060 23212 54572 23268
rect 54628 23212 57484 23268
rect 57540 23212 57550 23268
rect 60918 23212 60956 23268
rect 61012 23212 61022 23268
rect 3154 23100 3164 23156
rect 3220 23100 3500 23156
rect 3556 23100 3566 23156
rect 6626 23100 6636 23156
rect 6692 23100 8428 23156
rect 8484 23100 8494 23156
rect 13906 23100 13916 23156
rect 13972 23100 15148 23156
rect 15204 23100 15214 23156
rect 18274 23100 18284 23156
rect 18340 23100 19068 23156
rect 19124 23100 19134 23156
rect 23202 23100 23212 23156
rect 23268 23100 23278 23156
rect 24546 23100 24556 23156
rect 24612 23100 25228 23156
rect 25284 23100 25294 23156
rect 27794 23100 27804 23156
rect 27860 23100 29708 23156
rect 29764 23100 30380 23156
rect 30436 23100 30446 23156
rect 35410 23100 35420 23156
rect 35476 23100 36092 23156
rect 36148 23100 36158 23156
rect 36418 23100 36428 23156
rect 36484 23100 36652 23156
rect 36708 23100 37996 23156
rect 38052 23100 38062 23156
rect 39554 23100 39564 23156
rect 39620 23100 39630 23156
rect 42354 23100 42364 23156
rect 42420 23100 43260 23156
rect 43316 23100 43326 23156
rect 44930 23100 44940 23156
rect 44996 23100 46396 23156
rect 46452 23100 46462 23156
rect 46834 23100 46844 23156
rect 46900 23100 47852 23156
rect 47908 23100 47918 23156
rect 49858 23100 49868 23156
rect 49924 23100 50540 23156
rect 50596 23100 50606 23156
rect 51538 23100 51548 23156
rect 51604 23100 52892 23156
rect 52948 23100 52958 23156
rect 58594 23100 58604 23156
rect 58660 23100 61180 23156
rect 61236 23100 61246 23156
rect 4610 22988 4620 23044
rect 4676 22988 5628 23044
rect 5684 22988 5694 23044
rect 6962 22988 6972 23044
rect 7028 22988 7038 23044
rect 8082 22988 8092 23044
rect 8148 22988 9772 23044
rect 9828 22988 11004 23044
rect 11060 22988 11070 23044
rect 11228 22988 23548 23044
rect 23604 22988 27580 23044
rect 27636 22988 27646 23044
rect 29586 22988 29596 23044
rect 29652 22988 30492 23044
rect 30548 22988 30558 23044
rect 38322 22988 38332 23044
rect 38388 22988 41356 23044
rect 41412 22988 41422 23044
rect 48150 22988 48188 23044
rect 48244 22988 48254 23044
rect 52658 22988 52668 23044
rect 52724 22988 53452 23044
rect 53508 22988 54796 23044
rect 54852 22988 55580 23044
rect 55636 22988 55646 23044
rect 56018 22988 56028 23044
rect 56084 22988 57036 23044
rect 57092 22988 57102 23044
rect 6972 22932 7028 22988
rect 11228 22932 11284 22988
rect 3490 22876 3500 22932
rect 3556 22876 6412 22932
rect 6468 22876 6478 22932
rect 6972 22876 11284 22932
rect 13458 22876 13468 22932
rect 13524 22876 14140 22932
rect 14196 22876 15372 22932
rect 15428 22876 15438 22932
rect 16902 22876 16940 22932
rect 16996 22876 17006 22932
rect 18022 22876 18060 22932
rect 18116 22876 18126 22932
rect 28018 22876 28028 22932
rect 28084 22876 29260 22932
rect 29316 22876 29326 22932
rect 35858 22876 35868 22932
rect 35924 22876 37996 22932
rect 38052 22876 38062 22932
rect 39330 22876 39340 22932
rect 39396 22876 40012 22932
rect 40068 22876 41020 22932
rect 41076 22876 41086 22932
rect 46162 22876 46172 22932
rect 46228 22876 50428 22932
rect 51650 22876 51660 22932
rect 51716 22876 57260 22932
rect 57316 22876 57326 22932
rect 50372 22820 50428 22876
rect 1698 22764 1708 22820
rect 1764 22764 3164 22820
rect 3220 22764 3230 22820
rect 14886 22764 14924 22820
rect 14980 22764 14990 22820
rect 31042 22764 31052 22820
rect 31108 22764 31500 22820
rect 31556 22764 31566 22820
rect 34486 22764 34524 22820
rect 34580 22764 34590 22820
rect 39106 22764 39116 22820
rect 39172 22764 40572 22820
rect 40628 22764 40638 22820
rect 44706 22764 44716 22820
rect 44772 22764 47068 22820
rect 47124 22764 47134 22820
rect 50372 22764 58828 22820
rect 58884 22764 58894 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 13570 22652 13580 22708
rect 13636 22652 18956 22708
rect 19012 22652 26908 22708
rect 31266 22652 31276 22708
rect 31332 22652 32172 22708
rect 32228 22652 33068 22708
rect 33124 22652 33134 22708
rect 38612 22652 51996 22708
rect 52052 22652 52062 22708
rect 26852 22596 26908 22652
rect 38612 22596 38668 22652
rect 1698 22540 1708 22596
rect 1764 22540 2604 22596
rect 2660 22540 2670 22596
rect 10770 22540 10780 22596
rect 10836 22540 11788 22596
rect 11844 22540 11854 22596
rect 12002 22540 12012 22596
rect 12068 22540 12106 22596
rect 14438 22540 14476 22596
rect 14532 22540 14542 22596
rect 15026 22540 15036 22596
rect 15092 22540 15820 22596
rect 15876 22540 15886 22596
rect 26852 22540 29932 22596
rect 29988 22540 32060 22596
rect 32116 22540 32126 22596
rect 34514 22540 34524 22596
rect 34580 22540 35196 22596
rect 35252 22540 38668 22596
rect 41794 22540 41804 22596
rect 41860 22540 44828 22596
rect 44884 22540 44894 22596
rect 47842 22540 47852 22596
rect 47908 22540 49980 22596
rect 50036 22540 50046 22596
rect 59042 22540 59052 22596
rect 59108 22540 60620 22596
rect 60676 22540 60686 22596
rect 11218 22428 11228 22484
rect 11284 22428 16940 22484
rect 16996 22428 17276 22484
rect 17332 22428 17342 22484
rect 21634 22428 21644 22484
rect 21700 22428 25228 22484
rect 25284 22428 27468 22484
rect 27524 22428 29148 22484
rect 29204 22428 29214 22484
rect 32694 22428 32732 22484
rect 32788 22428 32798 22484
rect 33254 22428 33292 22484
rect 33348 22428 33358 22484
rect 43474 22428 43484 22484
rect 43540 22428 45276 22484
rect 45332 22428 45342 22484
rect 45490 22428 45500 22484
rect 45556 22428 45836 22484
rect 45892 22428 45902 22484
rect 4610 22316 4620 22372
rect 4676 22316 6972 22372
rect 7028 22316 8652 22372
rect 8708 22316 8718 22372
rect 11554 22316 11564 22372
rect 11620 22316 15988 22372
rect 16146 22316 16156 22372
rect 16212 22316 19516 22372
rect 19572 22316 19582 22372
rect 21746 22316 21756 22372
rect 21812 22316 22148 22372
rect 22418 22316 22428 22372
rect 22484 22316 23324 22372
rect 23380 22316 23390 22372
rect 24434 22316 24444 22372
rect 24500 22316 26460 22372
rect 26516 22316 26526 22372
rect 28466 22316 28476 22372
rect 28532 22316 29372 22372
rect 29428 22316 29438 22372
rect 31490 22316 31500 22372
rect 31556 22316 33964 22372
rect 34020 22316 34030 22372
rect 36306 22316 36316 22372
rect 36372 22316 37548 22372
rect 37604 22316 37614 22372
rect 39554 22316 39564 22372
rect 39620 22316 40684 22372
rect 40740 22316 41020 22372
rect 41076 22316 41086 22372
rect 43250 22316 43260 22372
rect 43316 22316 44828 22372
rect 44884 22316 44894 22372
rect 46610 22316 46620 22372
rect 46676 22316 51100 22372
rect 51156 22316 52108 22372
rect 52164 22316 52174 22372
rect 55794 22316 55804 22372
rect 55860 22316 58156 22372
rect 58212 22316 58222 22372
rect 8866 22204 8876 22260
rect 8932 22204 9660 22260
rect 9716 22204 10892 22260
rect 10948 22204 11676 22260
rect 11732 22204 11742 22260
rect 12310 22204 12348 22260
rect 12404 22204 12414 22260
rect 12898 22204 12908 22260
rect 12964 22204 15260 22260
rect 15316 22204 15326 22260
rect 15932 22148 15988 22316
rect 22092 22260 22148 22316
rect 16818 22204 16828 22260
rect 16884 22204 17612 22260
rect 17668 22204 22036 22260
rect 22092 22204 22316 22260
rect 22372 22204 22382 22260
rect 32274 22204 32284 22260
rect 32340 22204 33068 22260
rect 33124 22204 33134 22260
rect 47058 22204 47068 22260
rect 47124 22204 47852 22260
rect 47908 22204 48524 22260
rect 48580 22204 48590 22260
rect 49046 22204 49084 22260
rect 49140 22204 49150 22260
rect 49298 22204 49308 22260
rect 49364 22204 49644 22260
rect 49700 22204 51548 22260
rect 51604 22204 52668 22260
rect 52724 22204 52734 22260
rect 56018 22204 56028 22260
rect 56084 22204 57820 22260
rect 57876 22204 57886 22260
rect 21980 22148 22036 22204
rect 5058 22092 5068 22148
rect 5124 22092 5404 22148
rect 5460 22092 5470 22148
rect 6066 22092 6076 22148
rect 6132 22092 6412 22148
rect 6468 22092 6636 22148
rect 6692 22092 6702 22148
rect 12002 22092 12012 22148
rect 12068 22092 12572 22148
rect 12628 22092 13916 22148
rect 13972 22092 14924 22148
rect 14980 22092 14990 22148
rect 15932 22092 16940 22148
rect 16996 22092 18732 22148
rect 18788 22092 18798 22148
rect 21970 22092 21980 22148
rect 22036 22092 22046 22148
rect 24966 22092 25004 22148
rect 25060 22092 25070 22148
rect 28242 22092 28252 22148
rect 28308 22092 30716 22148
rect 30772 22092 30782 22148
rect 36390 22092 36428 22148
rect 36484 22092 36494 22148
rect 39330 22092 39340 22148
rect 39396 22092 40012 22148
rect 40068 22092 52108 22148
rect 52164 22092 52174 22148
rect 57138 22092 57148 22148
rect 57204 22092 57708 22148
rect 57764 22092 57774 22148
rect 59378 22092 59388 22148
rect 59444 22092 60956 22148
rect 61012 22092 61022 22148
rect 21410 21980 21420 22036
rect 21476 21980 21868 22036
rect 21924 21980 21934 22036
rect 32050 21980 32060 22036
rect 32116 21980 33516 22036
rect 33572 21980 33582 22036
rect 43362 21980 43372 22036
rect 43428 21980 43596 22036
rect 43652 21980 43662 22036
rect 51874 21980 51884 22036
rect 51940 21980 51950 22036
rect 57026 21980 57036 22036
rect 57092 21980 62188 22036
rect 62244 21980 62254 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 51884 21924 51940 21980
rect 1698 21868 1708 21924
rect 1764 21868 2156 21924
rect 2212 21868 2222 21924
rect 3378 21868 3388 21924
rect 3444 21868 9156 21924
rect 10994 21868 11004 21924
rect 11060 21868 11788 21924
rect 32162 21868 32172 21924
rect 32228 21868 32732 21924
rect 32788 21868 32798 21924
rect 43026 21868 43036 21924
rect 43092 21868 44548 21924
rect 47730 21868 47740 21924
rect 47796 21868 49420 21924
rect 49476 21868 49486 21924
rect 51538 21868 51548 21924
rect 51604 21868 53228 21924
rect 53284 21868 54012 21924
rect 54068 21868 54078 21924
rect 1810 21756 1820 21812
rect 1876 21756 3948 21812
rect 4004 21756 4014 21812
rect 4246 21756 4284 21812
rect 4340 21756 4350 21812
rect 5170 21756 5180 21812
rect 5236 21756 7532 21812
rect 7588 21756 7598 21812
rect 9100 21700 9156 21868
rect 11732 21812 11788 21868
rect 44492 21812 44548 21868
rect 9314 21756 9324 21812
rect 9380 21756 11116 21812
rect 11172 21756 11182 21812
rect 11732 21756 12012 21812
rect 12068 21756 12078 21812
rect 18610 21756 18620 21812
rect 18676 21756 19628 21812
rect 19684 21756 20076 21812
rect 20132 21756 20142 21812
rect 21298 21756 21308 21812
rect 21364 21756 23100 21812
rect 23156 21756 24668 21812
rect 24724 21756 24734 21812
rect 30930 21756 30940 21812
rect 30996 21756 31836 21812
rect 31892 21756 31902 21812
rect 32386 21756 32396 21812
rect 32452 21756 33292 21812
rect 33348 21756 33358 21812
rect 40114 21756 40124 21812
rect 40180 21756 41020 21812
rect 41076 21756 41086 21812
rect 41244 21756 42140 21812
rect 42196 21756 43148 21812
rect 43204 21756 43214 21812
rect 44482 21756 44492 21812
rect 44548 21756 45836 21812
rect 45892 21756 45902 21812
rect 47954 21756 47964 21812
rect 48020 21756 53340 21812
rect 53396 21756 53406 21812
rect 55346 21756 55356 21812
rect 55412 21756 60508 21812
rect 60564 21756 60574 21812
rect 41244 21700 41300 21756
rect 3490 21644 3500 21700
rect 3556 21644 4172 21700
rect 4228 21644 4238 21700
rect 9100 21644 11788 21700
rect 12674 21644 12684 21700
rect 12740 21644 15596 21700
rect 15652 21644 15662 21700
rect 16930 21644 16940 21700
rect 16996 21644 17612 21700
rect 17668 21644 19404 21700
rect 19460 21644 19470 21700
rect 19954 21644 19964 21700
rect 20020 21644 20030 21700
rect 20402 21644 20412 21700
rect 20468 21644 20972 21700
rect 21028 21644 22876 21700
rect 22932 21644 22942 21700
rect 23426 21644 23436 21700
rect 23492 21644 24220 21700
rect 24276 21644 25116 21700
rect 25172 21644 26460 21700
rect 26516 21644 26526 21700
rect 30258 21644 30268 21700
rect 30324 21644 34524 21700
rect 34580 21644 34590 21700
rect 35522 21644 35532 21700
rect 35588 21644 39116 21700
rect 39172 21644 39182 21700
rect 39442 21644 39452 21700
rect 39508 21644 41300 21700
rect 41458 21644 41468 21700
rect 41524 21644 42364 21700
rect 42420 21644 42430 21700
rect 43810 21644 43820 21700
rect 43876 21644 44716 21700
rect 44772 21644 44782 21700
rect 48290 21644 48300 21700
rect 48356 21644 48860 21700
rect 48916 21644 48926 21700
rect 49410 21644 49420 21700
rect 49476 21644 49644 21700
rect 49700 21644 49710 21700
rect 52434 21644 52444 21700
rect 52500 21644 55244 21700
rect 55300 21644 57372 21700
rect 57428 21644 57438 21700
rect 11732 21588 11788 21644
rect 19964 21588 20020 21644
rect 2482 21532 2492 21588
rect 2548 21532 3052 21588
rect 3108 21532 3118 21588
rect 4386 21532 4396 21588
rect 4452 21532 6188 21588
rect 6244 21532 6254 21588
rect 9090 21532 9100 21588
rect 9156 21532 11116 21588
rect 11172 21532 11182 21588
rect 11732 21532 20020 21588
rect 20626 21532 20636 21588
rect 20692 21532 20972 21588
rect 21028 21532 21084 21588
rect 21140 21532 21150 21588
rect 22306 21532 22316 21588
rect 22372 21532 24556 21588
rect 24612 21532 25340 21588
rect 25396 21532 25406 21588
rect 31154 21532 31164 21588
rect 31220 21532 33292 21588
rect 33348 21532 33358 21588
rect 34710 21532 34748 21588
rect 34804 21532 34814 21588
rect 35746 21532 35756 21588
rect 35812 21532 42028 21588
rect 42084 21532 42094 21588
rect 43586 21532 43596 21588
rect 43652 21532 44380 21588
rect 44436 21532 45052 21588
rect 45108 21532 45724 21588
rect 45780 21532 45790 21588
rect 47618 21532 47628 21588
rect 47684 21532 48972 21588
rect 49028 21532 49038 21588
rect 49494 21532 49532 21588
rect 49588 21532 49598 21588
rect 55010 21532 55020 21588
rect 55076 21532 57708 21588
rect 57764 21532 57774 21588
rect 57922 21532 57932 21588
rect 57988 21532 59052 21588
rect 59108 21532 60396 21588
rect 60452 21532 60462 21588
rect 4722 21420 4732 21476
rect 4788 21420 6300 21476
rect 6356 21420 6366 21476
rect 9874 21420 9884 21476
rect 9940 21420 9950 21476
rect 10770 21420 10780 21476
rect 10836 21420 12572 21476
rect 12628 21420 13020 21476
rect 13076 21420 13086 21476
rect 15026 21420 15036 21476
rect 15092 21420 17276 21476
rect 17332 21420 17342 21476
rect 19282 21420 19292 21476
rect 19348 21420 20076 21476
rect 20132 21420 20142 21476
rect 21634 21420 21644 21476
rect 21700 21420 23436 21476
rect 23492 21420 23502 21476
rect 29250 21420 29260 21476
rect 29316 21420 30044 21476
rect 30100 21420 34300 21476
rect 34356 21420 34366 21476
rect 47842 21420 47852 21476
rect 47908 21420 48860 21476
rect 48916 21420 48926 21476
rect 49074 21420 49084 21476
rect 49140 21420 49980 21476
rect 50036 21420 50046 21476
rect 53890 21420 53900 21476
rect 53956 21420 59500 21476
rect 59556 21420 59566 21476
rect 9884 21252 9940 21420
rect 10546 21308 10556 21364
rect 10612 21308 12012 21364
rect 12068 21308 12460 21364
rect 12516 21308 12526 21364
rect 14018 21308 14028 21364
rect 14084 21308 14700 21364
rect 14756 21308 14766 21364
rect 15922 21308 15932 21364
rect 15988 21308 16268 21364
rect 16324 21308 17836 21364
rect 17892 21308 17902 21364
rect 21970 21308 21980 21364
rect 22036 21308 23772 21364
rect 23828 21308 27356 21364
rect 27412 21308 27422 21364
rect 29922 21308 29932 21364
rect 29988 21308 31388 21364
rect 31444 21308 31454 21364
rect 32610 21308 32620 21364
rect 32676 21308 33068 21364
rect 33124 21308 44324 21364
rect 48402 21308 48412 21364
rect 48468 21308 49308 21364
rect 49364 21308 51436 21364
rect 51492 21308 53452 21364
rect 53508 21308 53518 21364
rect 53666 21308 53676 21364
rect 53732 21308 54460 21364
rect 54516 21308 54526 21364
rect 57250 21308 57260 21364
rect 57316 21308 59276 21364
rect 59332 21308 59342 21364
rect 60162 21308 60172 21364
rect 60228 21308 60844 21364
rect 60900 21308 61292 21364
rect 61348 21308 61358 21364
rect 9884 21196 24108 21252
rect 24164 21196 24174 21252
rect 24994 21196 25004 21252
rect 25060 21196 28028 21252
rect 28084 21196 33516 21252
rect 33572 21196 33582 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 44268 21140 44324 21308
rect 49634 21196 49644 21252
rect 49700 21196 53004 21252
rect 53060 21196 53070 21252
rect 54002 21196 54012 21252
rect 54068 21196 54684 21252
rect 54740 21196 57932 21252
rect 57988 21196 57998 21252
rect 58828 21140 58884 21308
rect 15586 21084 15596 21140
rect 15652 21084 16492 21140
rect 16548 21084 16558 21140
rect 22418 21084 22428 21140
rect 22484 21084 25228 21140
rect 25284 21084 25294 21140
rect 31602 21084 31612 21140
rect 31668 21084 32060 21140
rect 32116 21084 33068 21140
rect 33124 21084 33134 21140
rect 37986 21084 37996 21140
rect 38052 21084 39900 21140
rect 39956 21084 39966 21140
rect 44146 21084 44156 21140
rect 44212 21084 50092 21140
rect 50148 21084 50158 21140
rect 58818 21084 58828 21140
rect 58884 21084 58894 21140
rect 59826 21084 59836 21140
rect 59892 21084 60172 21140
rect 60228 21084 60238 21140
rect 2706 20972 2716 21028
rect 2772 20972 3276 21028
rect 3332 20972 3342 21028
rect 4162 20972 4172 21028
rect 4228 20972 5740 21028
rect 5796 20972 5806 21028
rect 6486 20972 6524 21028
rect 6580 20972 6590 21028
rect 14802 20972 14812 21028
rect 14868 20972 16828 21028
rect 16884 20972 17388 21028
rect 17444 20972 17454 21028
rect 19058 20972 19068 21028
rect 19124 20972 24892 21028
rect 24948 20972 24958 21028
rect 33394 20972 33404 21028
rect 33460 20972 52668 21028
rect 52724 20972 55804 21028
rect 55860 20972 55870 21028
rect 58370 20972 58380 21028
rect 58436 20972 58604 21028
rect 58660 20972 59052 21028
rect 59108 20972 59118 21028
rect 59938 20972 59948 21028
rect 60004 20972 61628 21028
rect 61684 20972 61694 21028
rect 5506 20860 5516 20916
rect 5572 20860 7756 20916
rect 7812 20860 7822 20916
rect 11890 20860 11900 20916
rect 11956 20860 12572 20916
rect 12628 20860 12638 20916
rect 17266 20860 17276 20916
rect 17332 20860 18844 20916
rect 18900 20860 19628 20916
rect 19684 20860 19694 20916
rect 31938 20860 31948 20916
rect 32004 20860 33852 20916
rect 33908 20860 33918 20916
rect 45938 20860 45948 20916
rect 46004 20860 49532 20916
rect 49588 20860 49868 20916
rect 49924 20860 49934 20916
rect 51174 20860 51212 20916
rect 51268 20860 51278 20916
rect 54338 20860 54348 20916
rect 54404 20860 56252 20916
rect 56308 20860 56318 20916
rect 59826 20860 59836 20916
rect 59892 20860 60620 20916
rect 60676 20860 61964 20916
rect 62020 20860 62030 20916
rect 2594 20748 2604 20804
rect 2660 20748 3052 20804
rect 3108 20748 3948 20804
rect 4004 20748 4014 20804
rect 4732 20748 5964 20804
rect 6020 20748 6030 20804
rect 8306 20748 8316 20804
rect 8372 20748 9548 20804
rect 9604 20748 9614 20804
rect 13682 20748 13692 20804
rect 13748 20748 15036 20804
rect 15092 20748 15484 20804
rect 15540 20748 15550 20804
rect 16034 20748 16044 20804
rect 16100 20748 20636 20804
rect 20692 20748 20702 20804
rect 32386 20748 32396 20804
rect 32452 20748 34972 20804
rect 35028 20748 35038 20804
rect 42130 20748 42140 20804
rect 42196 20748 43036 20804
rect 43092 20748 43102 20804
rect 43474 20748 43484 20804
rect 43540 20748 45164 20804
rect 45220 20748 45612 20804
rect 45668 20748 45678 20804
rect 54114 20748 54124 20804
rect 54180 20748 58380 20804
rect 58436 20748 58446 20804
rect 59042 20748 59052 20804
rect 59108 20748 60732 20804
rect 60788 20748 60798 20804
rect 60946 20748 60956 20804
rect 61012 20748 61022 20804
rect 4732 20580 4788 20748
rect 60956 20692 61012 20748
rect 6066 20636 6076 20692
rect 6132 20636 8092 20692
rect 8148 20636 8158 20692
rect 9426 20636 9436 20692
rect 9492 20636 10108 20692
rect 10164 20636 10174 20692
rect 14466 20636 14476 20692
rect 14532 20636 14924 20692
rect 14980 20636 15148 20692
rect 15362 20636 15372 20692
rect 15428 20636 16604 20692
rect 16660 20636 16670 20692
rect 30370 20636 30380 20692
rect 30436 20636 32508 20692
rect 32564 20636 32574 20692
rect 35074 20636 35084 20692
rect 35140 20636 37436 20692
rect 37492 20636 37502 20692
rect 48738 20636 48748 20692
rect 48804 20636 50204 20692
rect 50260 20636 50270 20692
rect 54562 20636 54572 20692
rect 54628 20636 56588 20692
rect 56644 20636 56654 20692
rect 60498 20636 60508 20692
rect 60564 20636 61012 20692
rect 15092 20580 15148 20636
rect 2594 20524 2604 20580
rect 2660 20524 3948 20580
rect 4004 20524 4788 20580
rect 5170 20524 5180 20580
rect 5236 20524 10332 20580
rect 10388 20524 10398 20580
rect 15092 20524 15596 20580
rect 15652 20524 15662 20580
rect 16482 20524 16492 20580
rect 16548 20524 17948 20580
rect 18004 20524 18014 20580
rect 26852 20524 30604 20580
rect 30660 20524 30670 20580
rect 30930 20524 30940 20580
rect 30996 20524 31500 20580
rect 31556 20524 31566 20580
rect 36306 20524 36316 20580
rect 36372 20524 42364 20580
rect 42420 20524 42430 20580
rect 42914 20524 42924 20580
rect 42980 20524 43820 20580
rect 43876 20524 43886 20580
rect 49046 20524 49084 20580
rect 49140 20524 49150 20580
rect 50988 20524 51436 20580
rect 51492 20524 51502 20580
rect 59042 20524 59052 20580
rect 59108 20524 61068 20580
rect 61124 20524 61134 20580
rect 7522 20412 7532 20468
rect 7588 20412 8988 20468
rect 9044 20412 9054 20468
rect 17266 20412 17276 20468
rect 17332 20412 17342 20468
rect 2146 20300 2156 20356
rect 2212 20300 2492 20356
rect 2548 20300 2558 20356
rect 8306 20300 8316 20356
rect 8372 20300 14476 20356
rect 14532 20300 14924 20356
rect 14980 20300 14990 20356
rect 6962 20188 6972 20244
rect 7028 20188 7756 20244
rect 7812 20188 8540 20244
rect 8596 20188 11900 20244
rect 11956 20188 11966 20244
rect 17276 20132 17332 20412
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 26852 20356 26908 20524
rect 50988 20468 51044 20524
rect 30706 20412 30716 20468
rect 30772 20412 30940 20468
rect 30996 20412 32620 20468
rect 32676 20412 32686 20468
rect 38994 20412 39004 20468
rect 39060 20412 40684 20468
rect 40740 20412 40750 20468
rect 50978 20412 50988 20468
rect 51044 20412 51054 20468
rect 61142 20412 61180 20468
rect 61236 20412 61246 20468
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 23426 20300 23436 20356
rect 23492 20300 26908 20356
rect 30146 20300 30156 20356
rect 30212 20300 31052 20356
rect 31108 20300 31118 20356
rect 40338 20300 40348 20356
rect 40404 20300 41356 20356
rect 41412 20300 41804 20356
rect 41860 20300 42252 20356
rect 42308 20300 42318 20356
rect 43138 20300 43148 20356
rect 43204 20300 47628 20356
rect 47684 20300 47694 20356
rect 59826 20300 59836 20356
rect 59892 20300 62076 20356
rect 62132 20300 62142 20356
rect 20178 20188 20188 20244
rect 20244 20188 21756 20244
rect 21812 20188 21822 20244
rect 23314 20188 23324 20244
rect 23380 20188 24332 20244
rect 24388 20188 24398 20244
rect 29810 20188 29820 20244
rect 29876 20188 30940 20244
rect 30996 20188 31006 20244
rect 32498 20188 32508 20244
rect 32564 20188 32956 20244
rect 33012 20188 33022 20244
rect 34748 20188 35308 20244
rect 35364 20188 35374 20244
rect 38546 20188 38556 20244
rect 38612 20188 40124 20244
rect 40180 20188 41692 20244
rect 41748 20188 44156 20244
rect 44212 20188 44222 20244
rect 51762 20188 51772 20244
rect 51828 20188 52892 20244
rect 52948 20188 52958 20244
rect 55010 20188 55020 20244
rect 55076 20188 56140 20244
rect 56196 20188 56206 20244
rect 57586 20188 57596 20244
rect 57652 20188 57662 20244
rect 61394 20188 61404 20244
rect 61460 20188 61470 20244
rect 34748 20132 34804 20188
rect 57596 20132 57652 20188
rect 61404 20132 61460 20188
rect 1922 20076 1932 20132
rect 1988 20076 5180 20132
rect 5236 20076 5246 20132
rect 6626 20076 6636 20132
rect 6692 20076 8988 20132
rect 9044 20076 11788 20132
rect 11844 20076 11854 20132
rect 12562 20076 12572 20132
rect 12628 20076 14700 20132
rect 14756 20076 14766 20132
rect 15474 20076 15484 20132
rect 15540 20076 17332 20132
rect 20626 20076 20636 20132
rect 20692 20076 22092 20132
rect 22148 20076 22158 20132
rect 24098 20076 24108 20132
rect 24164 20076 24174 20132
rect 24658 20076 24668 20132
rect 24724 20076 26684 20132
rect 26740 20076 26750 20132
rect 27234 20076 27244 20132
rect 27300 20076 30492 20132
rect 30548 20076 31164 20132
rect 31220 20076 31230 20132
rect 34738 20076 34748 20132
rect 34804 20076 34814 20132
rect 34962 20076 34972 20132
rect 35028 20076 35756 20132
rect 35812 20076 35822 20132
rect 35970 20076 35980 20132
rect 36036 20076 37772 20132
rect 37828 20076 37838 20132
rect 47730 20076 47740 20132
rect 47796 20076 48860 20132
rect 48916 20076 48926 20132
rect 50866 20076 50876 20132
rect 50932 20076 52220 20132
rect 52276 20076 52286 20132
rect 54450 20076 54460 20132
rect 54516 20076 57652 20132
rect 60274 20076 60284 20132
rect 60340 20076 61460 20132
rect 24108 20020 24164 20076
rect 5254 19964 5292 20020
rect 5348 19964 5358 20020
rect 5954 19964 5964 20020
rect 6020 19964 6524 20020
rect 6580 19964 7196 20020
rect 7252 19964 7262 20020
rect 7858 19964 7868 20020
rect 7924 19964 9772 20020
rect 9828 19964 9838 20020
rect 9986 19964 9996 20020
rect 10052 19964 12012 20020
rect 12068 19964 12078 20020
rect 13122 19964 13132 20020
rect 13188 19964 15372 20020
rect 15428 19964 15438 20020
rect 15586 19964 15596 20020
rect 15652 19964 16268 20020
rect 16324 19964 16334 20020
rect 16706 19964 16716 20020
rect 16772 19964 20524 20020
rect 20580 19964 20590 20020
rect 21410 19964 21420 20020
rect 21476 19964 21868 20020
rect 21924 19964 21934 20020
rect 24108 19964 24892 20020
rect 24948 19964 25452 20020
rect 25508 19964 25518 20020
rect 27122 19964 27132 20020
rect 27188 19964 28252 20020
rect 28308 19964 29820 20020
rect 29876 19964 33516 20020
rect 33572 19964 34188 20020
rect 34244 19964 34254 20020
rect 36082 19964 36092 20020
rect 36148 19964 37212 20020
rect 37268 19964 37660 20020
rect 37716 19964 37726 20020
rect 45490 19964 45500 20020
rect 45556 19964 47068 20020
rect 47124 19964 47134 20020
rect 47282 19964 47292 20020
rect 47348 19964 49308 20020
rect 49364 19964 49374 20020
rect 52098 19964 52108 20020
rect 52164 19964 52174 20020
rect 53666 19964 53676 20020
rect 53732 19964 55692 20020
rect 55748 19964 57036 20020
rect 57092 19964 57102 20020
rect 58258 19964 58268 20020
rect 58324 19964 61404 20020
rect 61460 19964 61470 20020
rect 6402 19852 6412 19908
rect 6468 19852 8652 19908
rect 8708 19852 12348 19908
rect 12404 19852 12414 19908
rect 18050 19852 18060 19908
rect 18116 19852 18620 19908
rect 18676 19852 18686 19908
rect 24098 19852 24108 19908
rect 24164 19852 26236 19908
rect 26292 19852 26302 19908
rect 26852 19852 27692 19908
rect 27748 19852 27758 19908
rect 29362 19852 29372 19908
rect 29428 19852 32732 19908
rect 32788 19852 33292 19908
rect 33348 19852 33358 19908
rect 34514 19852 34524 19908
rect 34580 19852 35196 19908
rect 35252 19852 35262 19908
rect 35970 19852 35980 19908
rect 36036 19852 37324 19908
rect 37380 19852 39116 19908
rect 39172 19852 39182 19908
rect 45602 19852 45612 19908
rect 45668 19852 48748 19908
rect 48804 19852 48814 19908
rect 26852 19796 26908 19852
rect 52108 19796 52164 19964
rect 54562 19852 54572 19908
rect 54628 19852 56588 19908
rect 56644 19852 56654 19908
rect 57586 19852 57596 19908
rect 57652 19852 61964 19908
rect 62020 19852 62030 19908
rect 2930 19740 2940 19796
rect 2996 19740 3836 19796
rect 3892 19740 4620 19796
rect 4676 19740 4686 19796
rect 4946 19740 4956 19796
rect 5012 19740 6300 19796
rect 6356 19740 7756 19796
rect 7812 19740 7822 19796
rect 12338 19740 12348 19796
rect 12404 19740 13468 19796
rect 13524 19740 14700 19796
rect 14756 19740 14766 19796
rect 18722 19740 18732 19796
rect 18788 19740 24220 19796
rect 24276 19740 24286 19796
rect 26338 19740 26348 19796
rect 26404 19740 26908 19796
rect 40674 19740 40684 19796
rect 40740 19740 43596 19796
rect 43652 19740 43662 19796
rect 52108 19740 58156 19796
rect 58212 19740 58716 19796
rect 58772 19740 58782 19796
rect 6486 19628 6524 19684
rect 6580 19628 6590 19684
rect 25218 19628 25228 19684
rect 25284 19628 30380 19684
rect 30436 19628 30446 19684
rect 41570 19628 41580 19684
rect 41636 19628 59052 19684
rect 59108 19628 59118 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 4946 19516 4956 19572
rect 5012 19516 9884 19572
rect 9940 19516 9950 19572
rect 11452 19516 13692 19572
rect 13748 19516 25564 19572
rect 25620 19516 25630 19572
rect 40338 19516 40348 19572
rect 40404 19516 41244 19572
rect 41300 19516 41310 19572
rect 43026 19516 43036 19572
rect 43092 19516 51660 19572
rect 51716 19516 51726 19572
rect 58034 19516 58044 19572
rect 58100 19516 61852 19572
rect 61908 19516 61918 19572
rect 3266 19404 3276 19460
rect 3332 19348 3388 19460
rect 8642 19404 8652 19460
rect 8708 19404 11228 19460
rect 11284 19404 11294 19460
rect 11452 19348 11508 19516
rect 13794 19404 13804 19460
rect 13860 19404 14588 19460
rect 14644 19404 15148 19460
rect 19506 19404 19516 19460
rect 19572 19404 20076 19460
rect 20132 19404 21420 19460
rect 21476 19404 21486 19460
rect 26674 19404 26684 19460
rect 26740 19404 29820 19460
rect 29876 19404 33292 19460
rect 33348 19404 33358 19460
rect 39890 19404 39900 19460
rect 39956 19404 47236 19460
rect 49410 19404 49420 19460
rect 49476 19404 52108 19460
rect 52164 19404 52174 19460
rect 59826 19404 59836 19460
rect 59892 19404 62860 19460
rect 62916 19404 62926 19460
rect 3332 19292 11508 19348
rect 15092 19348 15148 19404
rect 15092 19292 16940 19348
rect 16996 19292 17006 19348
rect 30146 19292 30156 19348
rect 30212 19292 31948 19348
rect 32004 19292 32014 19348
rect 33842 19292 33852 19348
rect 33908 19292 34972 19348
rect 35028 19292 35038 19348
rect 35410 19292 35420 19348
rect 35476 19292 36540 19348
rect 36596 19292 36606 19348
rect 40226 19292 40236 19348
rect 40292 19292 42252 19348
rect 42308 19292 42318 19348
rect 45602 19292 45612 19348
rect 45668 19292 46060 19348
rect 46116 19292 46126 19348
rect 46386 19292 46396 19348
rect 46452 19292 46844 19348
rect 46900 19292 46910 19348
rect 6962 19180 6972 19236
rect 7028 19180 8092 19236
rect 8148 19180 9436 19236
rect 9492 19180 9884 19236
rect 9940 19180 9950 19236
rect 10210 19180 10220 19236
rect 10276 19180 11788 19236
rect 11844 19180 11854 19236
rect 12310 19180 12348 19236
rect 12404 19180 12414 19236
rect 15698 19180 15708 19236
rect 15764 19180 16828 19236
rect 16884 19180 16894 19236
rect 24668 19180 26348 19236
rect 26404 19180 26414 19236
rect 34178 19180 34188 19236
rect 34244 19180 35756 19236
rect 35812 19180 35822 19236
rect 39106 19180 39116 19236
rect 39172 19180 41020 19236
rect 41076 19180 41086 19236
rect 45164 19180 46172 19236
rect 46228 19180 46238 19236
rect 24668 19124 24724 19180
rect 45164 19124 45220 19180
rect 47180 19124 47236 19404
rect 47730 19180 47740 19236
rect 47796 19180 49084 19236
rect 49140 19180 49150 19236
rect 54674 19180 54684 19236
rect 54740 19180 56252 19236
rect 56308 19180 56318 19236
rect 56690 19180 56700 19236
rect 56756 19180 58156 19236
rect 58212 19180 58222 19236
rect 60498 19180 60508 19236
rect 60564 19180 61628 19236
rect 61684 19180 61694 19236
rect 4722 19068 4732 19124
rect 4788 19068 5628 19124
rect 5684 19068 6636 19124
rect 6692 19068 6702 19124
rect 10546 19068 10556 19124
rect 10612 19068 12124 19124
rect 12180 19068 14252 19124
rect 14308 19068 14318 19124
rect 18274 19068 18284 19124
rect 18340 19068 22316 19124
rect 22372 19068 22382 19124
rect 24322 19068 24332 19124
rect 24388 19068 24668 19124
rect 24724 19068 24734 19124
rect 26226 19068 26236 19124
rect 26292 19068 30492 19124
rect 30548 19068 30558 19124
rect 34066 19068 34076 19124
rect 34132 19068 34142 19124
rect 35756 19068 45220 19124
rect 45490 19068 45500 19124
rect 45556 19068 46844 19124
rect 46900 19068 46910 19124
rect 47180 19068 53116 19124
rect 53172 19068 54348 19124
rect 54404 19068 54414 19124
rect 55794 19068 55804 19124
rect 55860 19068 56812 19124
rect 56868 19068 56878 19124
rect 59938 19068 59948 19124
rect 60004 19068 61404 19124
rect 61460 19068 61470 19124
rect 6738 18956 6748 19012
rect 6804 18956 13020 19012
rect 13076 18956 13086 19012
rect 23650 18956 23660 19012
rect 23716 18956 24220 19012
rect 24276 18956 24286 19012
rect 24882 18956 24892 19012
rect 24948 18956 25004 19012
rect 25060 18956 27020 19012
rect 27076 18956 29036 19012
rect 29092 18956 29102 19012
rect 34076 18900 34132 19068
rect 35756 19012 35812 19068
rect 34290 18956 34300 19012
rect 34356 18956 35812 19012
rect 36082 18956 36092 19012
rect 36148 18956 37100 19012
rect 37156 18956 38108 19012
rect 38164 18956 38174 19012
rect 43922 18956 43932 19012
rect 43988 18956 47068 19012
rect 47124 18956 47134 19012
rect 51538 18956 51548 19012
rect 51604 18956 53228 19012
rect 53284 18956 53294 19012
rect 59826 18956 59836 19012
rect 59892 18956 60284 19012
rect 60340 18956 61628 19012
rect 61684 18956 61694 19012
rect 7746 18844 7756 18900
rect 7812 18844 8316 18900
rect 8372 18844 8382 18900
rect 24546 18844 24556 18900
rect 24612 18844 26684 18900
rect 26740 18844 34132 18900
rect 44930 18844 44940 18900
rect 44996 18844 45612 18900
rect 45668 18844 46956 18900
rect 47012 18844 47022 18900
rect 49382 18844 49420 18900
rect 49476 18844 49486 18900
rect 53666 18844 53676 18900
rect 53732 18844 61404 18900
rect 61460 18844 62188 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 3574 18732 3612 18788
rect 3668 18732 3678 18788
rect 29698 18732 29708 18788
rect 29764 18732 35532 18788
rect 35588 18732 35598 18788
rect 36194 18732 36204 18788
rect 36260 18732 36270 18788
rect 58034 18732 58044 18788
rect 58100 18732 58492 18788
rect 58548 18732 60508 18788
rect 60564 18732 60574 18788
rect 62132 18732 62188 18844
rect 62244 18732 62254 18788
rect 1586 18620 1596 18676
rect 1652 18620 5292 18676
rect 5348 18620 5358 18676
rect 10322 18620 10332 18676
rect 10388 18620 12236 18676
rect 12292 18620 12302 18676
rect 13010 18620 13020 18676
rect 13076 18620 13356 18676
rect 13412 18620 13422 18676
rect 15026 18620 15036 18676
rect 15092 18620 15484 18676
rect 15540 18620 15550 18676
rect 24658 18620 24668 18676
rect 24724 18620 25900 18676
rect 25956 18620 25966 18676
rect 30482 18620 30492 18676
rect 30548 18620 34748 18676
rect 34804 18620 34814 18676
rect 36204 18564 36260 18732
rect 38322 18620 38332 18676
rect 38388 18620 39452 18676
rect 39508 18620 39518 18676
rect 42690 18620 42700 18676
rect 42756 18620 44044 18676
rect 44100 18620 44110 18676
rect 49606 18620 49644 18676
rect 49700 18620 50988 18676
rect 51044 18620 51054 18676
rect 53778 18620 53788 18676
rect 53844 18620 56252 18676
rect 56308 18620 56318 18676
rect 60834 18620 60844 18676
rect 60900 18620 60956 18676
rect 61012 18620 61022 18676
rect 2034 18508 2044 18564
rect 2100 18508 3948 18564
rect 4004 18508 4014 18564
rect 11890 18508 11900 18564
rect 11956 18508 12684 18564
rect 12740 18508 12750 18564
rect 22418 18508 22428 18564
rect 22484 18508 25788 18564
rect 25844 18508 27244 18564
rect 27300 18508 27310 18564
rect 32722 18508 32732 18564
rect 32788 18508 33796 18564
rect 36204 18508 42812 18564
rect 42868 18508 44156 18564
rect 44212 18508 44222 18564
rect 46722 18508 46732 18564
rect 46788 18508 48748 18564
rect 48804 18508 48814 18564
rect 51762 18508 51772 18564
rect 51828 18508 52556 18564
rect 52612 18508 52622 18564
rect 59378 18508 59388 18564
rect 59444 18508 59948 18564
rect 60004 18508 60014 18564
rect 1474 18396 1484 18452
rect 1540 18396 2716 18452
rect 2772 18396 2782 18452
rect 3332 18396 3612 18452
rect 3668 18396 5516 18452
rect 5572 18396 5582 18452
rect 5954 18396 5964 18452
rect 6020 18396 6524 18452
rect 6580 18396 6590 18452
rect 6738 18396 6748 18452
rect 6804 18396 6972 18452
rect 7028 18396 7038 18452
rect 11330 18396 11340 18452
rect 11396 18396 13468 18452
rect 13524 18396 13534 18452
rect 13794 18396 13804 18452
rect 13860 18396 14364 18452
rect 14420 18396 14430 18452
rect 15138 18396 15148 18452
rect 15204 18396 16492 18452
rect 16548 18396 18956 18452
rect 19012 18396 20300 18452
rect 20356 18396 20366 18452
rect 20514 18396 20524 18452
rect 20580 18396 21980 18452
rect 22036 18396 22046 18452
rect 22194 18396 22204 18452
rect 22260 18396 24892 18452
rect 24948 18396 24958 18452
rect 29474 18396 29484 18452
rect 29540 18396 30716 18452
rect 30772 18396 30782 18452
rect 30930 18396 30940 18452
rect 30996 18396 32396 18452
rect 32452 18396 33068 18452
rect 33124 18396 33134 18452
rect 3332 18228 3388 18396
rect 33740 18340 33796 18508
rect 34066 18396 34076 18452
rect 34132 18396 35084 18452
rect 35140 18396 36428 18452
rect 36484 18396 36494 18452
rect 36652 18396 39788 18452
rect 39844 18396 39854 18452
rect 42130 18396 42140 18452
rect 42196 18396 42700 18452
rect 42756 18396 44828 18452
rect 44884 18396 44894 18452
rect 45378 18396 45388 18452
rect 45444 18396 45948 18452
rect 46004 18396 46014 18452
rect 46274 18396 46284 18452
rect 46340 18396 48860 18452
rect 48916 18396 48926 18452
rect 52882 18396 52892 18452
rect 52948 18396 54908 18452
rect 54964 18396 56364 18452
rect 56420 18396 56430 18452
rect 57138 18396 57148 18452
rect 57204 18396 59836 18452
rect 59892 18396 59902 18452
rect 60050 18396 60060 18452
rect 60116 18396 62076 18452
rect 62132 18396 62142 18452
rect 5506 18284 5516 18340
rect 5572 18284 8316 18340
rect 8372 18284 8382 18340
rect 9762 18284 9772 18340
rect 9828 18284 15148 18340
rect 16930 18284 16940 18340
rect 16996 18284 19068 18340
rect 19124 18284 19134 18340
rect 21718 18284 21756 18340
rect 21812 18284 21822 18340
rect 23762 18284 23772 18340
rect 23828 18284 27020 18340
rect 27076 18284 29204 18340
rect 33730 18284 33740 18340
rect 33796 18284 33806 18340
rect 35186 18284 35196 18340
rect 35252 18284 36092 18340
rect 36148 18284 36158 18340
rect 2258 18172 2268 18228
rect 2324 18172 3388 18228
rect 3938 18172 3948 18228
rect 4004 18172 4900 18228
rect 8194 18172 8204 18228
rect 8260 18172 9548 18228
rect 9604 18172 10220 18228
rect 10276 18172 10286 18228
rect 4844 18116 4900 18172
rect 15092 18116 15148 18284
rect 29148 18228 29204 18284
rect 36652 18228 36708 18396
rect 38210 18284 38220 18340
rect 38276 18284 39564 18340
rect 39620 18284 39630 18340
rect 40002 18284 40012 18340
rect 40068 18284 43036 18340
rect 43092 18284 43102 18340
rect 43586 18284 43596 18340
rect 43652 18284 45500 18340
rect 45556 18284 46508 18340
rect 46564 18284 46574 18340
rect 50054 18284 50092 18340
rect 50148 18284 50158 18340
rect 51874 18284 51884 18340
rect 51940 18284 53116 18340
rect 53172 18284 53182 18340
rect 53554 18284 53564 18340
rect 53620 18284 57204 18340
rect 58818 18284 58828 18340
rect 58884 18284 61292 18340
rect 61348 18284 61358 18340
rect 61814 18284 61852 18340
rect 61908 18284 61918 18340
rect 57148 18228 57204 18284
rect 16034 18172 16044 18228
rect 16100 18172 16268 18228
rect 16324 18172 18508 18228
rect 18564 18172 18574 18228
rect 23492 18172 25004 18228
rect 25060 18172 25070 18228
rect 25554 18172 25564 18228
rect 25620 18172 28364 18228
rect 28420 18172 28430 18228
rect 29138 18172 29148 18228
rect 29204 18172 29214 18228
rect 33842 18172 33852 18228
rect 33908 18172 35420 18228
rect 35476 18172 35588 18228
rect 35858 18172 35868 18228
rect 35924 18172 36708 18228
rect 43138 18172 43148 18228
rect 43204 18172 43708 18228
rect 43764 18172 52220 18228
rect 52276 18172 52286 18228
rect 53330 18172 53340 18228
rect 53396 18172 54348 18228
rect 54404 18172 54414 18228
rect 55682 18172 55692 18228
rect 55748 18172 56588 18228
rect 56644 18172 56654 18228
rect 57138 18172 57148 18228
rect 57204 18172 58492 18228
rect 58548 18172 58558 18228
rect 23492 18116 23548 18172
rect 28364 18116 28420 18172
rect 4844 18060 11900 18116
rect 11956 18060 12908 18116
rect 12964 18060 12974 18116
rect 15092 18060 23548 18116
rect 23874 18060 23884 18116
rect 23940 18060 26796 18116
rect 26852 18060 26862 18116
rect 28364 18060 29260 18116
rect 29316 18060 29596 18116
rect 29652 18060 29662 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 35532 18004 35588 18172
rect 36978 18060 36988 18116
rect 37044 18060 42812 18116
rect 42868 18060 45836 18116
rect 45892 18060 45902 18116
rect 55570 18060 55580 18116
rect 55636 18060 56252 18116
rect 56308 18060 56318 18116
rect 6626 17948 6636 18004
rect 6692 17948 11340 18004
rect 11396 17948 11406 18004
rect 26450 17948 26460 18004
rect 26516 17948 35028 18004
rect 35532 17948 36652 18004
rect 36708 17948 36718 18004
rect 38612 17948 40796 18004
rect 40852 17948 40862 18004
rect 51874 17948 51884 18004
rect 51940 17948 53676 18004
rect 53732 17948 57036 18004
rect 57092 17948 60900 18004
rect 6636 17892 6692 17948
rect 34972 17892 35028 17948
rect 38612 17892 38668 17948
rect 3042 17836 3052 17892
rect 3108 17836 3118 17892
rect 3332 17836 6692 17892
rect 10994 17836 11004 17892
rect 11060 17836 12012 17892
rect 12068 17836 13580 17892
rect 13636 17836 13646 17892
rect 15250 17836 15260 17892
rect 15316 17836 17388 17892
rect 17444 17836 17454 17892
rect 18050 17836 18060 17892
rect 18116 17836 18732 17892
rect 18788 17836 20524 17892
rect 20580 17836 20590 17892
rect 25666 17836 25676 17892
rect 25732 17836 29708 17892
rect 29764 17836 33516 17892
rect 33572 17836 33582 17892
rect 34972 17836 37996 17892
rect 38052 17836 38668 17892
rect 44940 17836 45276 17892
rect 45332 17836 46508 17892
rect 46564 17836 46574 17892
rect 48626 17836 48636 17892
rect 48692 17836 50204 17892
rect 50260 17836 50270 17892
rect 52098 17836 52108 17892
rect 52164 17836 53564 17892
rect 53620 17836 53630 17892
rect 59490 17836 59500 17892
rect 59556 17836 60620 17892
rect 60676 17836 60686 17892
rect 3052 17780 3108 17836
rect 3332 17780 3388 17836
rect 44940 17780 44996 17836
rect 60844 17780 60900 17948
rect 914 17724 924 17780
rect 980 17724 2044 17780
rect 2100 17724 2110 17780
rect 3052 17724 3388 17780
rect 3686 17724 3724 17780
rect 3780 17724 3790 17780
rect 5618 17724 5628 17780
rect 5684 17724 6860 17780
rect 6916 17724 7980 17780
rect 8036 17724 8046 17780
rect 13122 17724 13132 17780
rect 13188 17724 14364 17780
rect 14420 17724 14430 17780
rect 18610 17724 18620 17780
rect 18676 17724 20076 17780
rect 20132 17724 20636 17780
rect 20692 17724 20702 17780
rect 25890 17724 25900 17780
rect 25956 17724 30380 17780
rect 30436 17724 30446 17780
rect 34514 17724 34524 17780
rect 34580 17724 35868 17780
rect 35924 17724 35934 17780
rect 36082 17724 36092 17780
rect 36148 17724 37884 17780
rect 37940 17724 37950 17780
rect 38434 17724 38444 17780
rect 38500 17724 44996 17780
rect 45714 17724 45724 17780
rect 45780 17724 50428 17780
rect 51650 17724 51660 17780
rect 51716 17724 53788 17780
rect 53844 17724 57372 17780
rect 57428 17724 60508 17780
rect 60564 17724 60574 17780
rect 60722 17724 60732 17780
rect 60788 17724 60900 17780
rect 61618 17724 61628 17780
rect 61684 17724 62972 17780
rect 63028 17724 63038 17780
rect 50372 17668 50428 17724
rect 4386 17612 4396 17668
rect 4452 17612 4956 17668
rect 5012 17612 5022 17668
rect 7410 17612 7420 17668
rect 7476 17612 9884 17668
rect 9940 17612 9950 17668
rect 16594 17612 16604 17668
rect 16660 17612 18172 17668
rect 18228 17612 18956 17668
rect 19012 17612 20188 17668
rect 20244 17612 20254 17668
rect 27234 17612 27244 17668
rect 27300 17612 28476 17668
rect 28532 17612 28542 17668
rect 30818 17612 30828 17668
rect 30884 17612 31052 17668
rect 31108 17612 31948 17668
rect 32004 17612 32014 17668
rect 41122 17612 41132 17668
rect 41188 17612 47852 17668
rect 47908 17612 47918 17668
rect 49046 17612 49084 17668
rect 49140 17612 49150 17668
rect 50372 17612 54740 17668
rect 57026 17612 57036 17668
rect 57092 17612 61852 17668
rect 61908 17612 61918 17668
rect 9436 17444 9492 17612
rect 54684 17556 54740 17612
rect 15586 17500 15596 17556
rect 15652 17500 16492 17556
rect 16548 17500 16558 17556
rect 24882 17500 24892 17556
rect 24948 17500 32396 17556
rect 32452 17500 32462 17556
rect 39442 17500 39452 17556
rect 39508 17500 39900 17556
rect 39956 17500 39966 17556
rect 40786 17500 40796 17556
rect 40852 17500 41356 17556
rect 41412 17500 41422 17556
rect 42242 17500 42252 17556
rect 42308 17500 43708 17556
rect 43764 17500 43774 17556
rect 48972 17500 49308 17556
rect 49364 17500 49374 17556
rect 49494 17500 49532 17556
rect 49588 17500 50204 17556
rect 50260 17500 50270 17556
rect 53218 17500 53228 17556
rect 53284 17500 54460 17556
rect 54516 17500 54526 17556
rect 54684 17500 58940 17556
rect 58996 17500 59006 17556
rect 60806 17500 60844 17556
rect 60900 17500 60910 17556
rect 4946 17388 4956 17444
rect 5012 17388 6300 17444
rect 6356 17388 6366 17444
rect 9426 17388 9436 17444
rect 9492 17388 9502 17444
rect 11666 17388 11676 17444
rect 11732 17388 14252 17444
rect 14308 17388 16100 17444
rect 24658 17388 24668 17444
rect 24724 17388 24780 17444
rect 24836 17388 25116 17444
rect 25172 17388 25182 17444
rect 27346 17388 27356 17444
rect 27412 17388 29148 17444
rect 29204 17388 32172 17444
rect 32228 17388 32238 17444
rect 35858 17388 35868 17444
rect 35924 17388 36316 17444
rect 36372 17388 36988 17444
rect 37044 17388 37054 17444
rect 43250 17388 43260 17444
rect 43316 17388 44044 17444
rect 44100 17388 44110 17444
rect 2818 17276 2828 17332
rect 2884 17276 10780 17332
rect 10836 17276 10846 17332
rect 5954 17164 5964 17220
rect 6020 17164 8316 17220
rect 8372 17164 8988 17220
rect 9044 17164 9884 17220
rect 9940 17164 10668 17220
rect 10724 17164 10734 17220
rect 16044 17108 16100 17388
rect 43586 17276 43596 17332
rect 43652 17276 45724 17332
rect 45780 17276 45790 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 48972 17220 49028 17500
rect 49158 17388 49196 17444
rect 49252 17388 49262 17444
rect 54338 17388 54348 17444
rect 54404 17388 57708 17444
rect 57764 17388 57774 17444
rect 61394 17388 61404 17444
rect 61460 17388 62076 17444
rect 62132 17388 62142 17444
rect 49970 17276 49980 17332
rect 50036 17276 50046 17332
rect 23762 17164 23772 17220
rect 23828 17164 26348 17220
rect 26404 17164 28196 17220
rect 38882 17164 38892 17220
rect 38948 17164 42084 17220
rect 48962 17164 48972 17220
rect 49028 17164 49038 17220
rect 2594 17052 2604 17108
rect 2660 17052 3388 17108
rect 3938 17052 3948 17108
rect 4004 17052 4396 17108
rect 4452 17052 4462 17108
rect 5842 17052 5852 17108
rect 5908 17052 10108 17108
rect 10164 17052 10174 17108
rect 13122 17052 13132 17108
rect 13188 17052 15484 17108
rect 15540 17052 15550 17108
rect 16034 17052 16044 17108
rect 16100 17052 16110 17108
rect 17602 17052 17612 17108
rect 17668 17052 24556 17108
rect 24612 17052 24780 17108
rect 24836 17052 25004 17108
rect 25060 17052 25070 17108
rect 26002 17052 26012 17108
rect 26068 17052 27244 17108
rect 27300 17052 27310 17108
rect 3332 16996 3388 17052
rect 28140 16996 28196 17164
rect 28914 17052 28924 17108
rect 28980 17052 30380 17108
rect 30436 17052 30446 17108
rect 33282 17052 33292 17108
rect 33348 17052 34412 17108
rect 34468 17052 34478 17108
rect 3332 16940 6748 16996
rect 6804 16940 6814 16996
rect 6962 16940 6972 16996
rect 7028 16940 8428 16996
rect 8484 16940 9548 16996
rect 9604 16940 9614 16996
rect 13794 16940 13804 16996
rect 13860 16940 14252 16996
rect 14308 16940 14476 16996
rect 14532 16940 16268 16996
rect 16324 16940 16334 16996
rect 16706 16940 16716 16996
rect 16772 16940 17388 16996
rect 17444 16940 17454 16996
rect 17938 16940 17948 16996
rect 18004 16940 20412 16996
rect 20468 16940 21644 16996
rect 21700 16940 21710 16996
rect 23202 16940 23212 16996
rect 23268 16940 23884 16996
rect 23940 16940 23950 16996
rect 25778 16940 25788 16996
rect 25844 16940 26908 16996
rect 28130 16940 28140 16996
rect 28196 16940 32060 16996
rect 32116 16940 32126 16996
rect 26852 16884 26908 16940
rect 4246 16828 4284 16884
rect 4340 16828 4350 16884
rect 6850 16828 6860 16884
rect 6916 16828 11004 16884
rect 11060 16828 11070 16884
rect 12898 16828 12908 16884
rect 12964 16828 13580 16884
rect 13636 16828 14140 16884
rect 14196 16828 15484 16884
rect 15540 16828 15550 16884
rect 21522 16828 21532 16884
rect 21588 16828 23548 16884
rect 23604 16828 23614 16884
rect 26852 16828 27020 16884
rect 27076 16828 28924 16884
rect 28980 16828 28990 16884
rect 29922 16828 29932 16884
rect 29988 16828 31948 16884
rect 32004 16828 32014 16884
rect 37874 16828 37884 16884
rect 37940 16828 38444 16884
rect 38500 16828 38510 16884
rect 39890 16828 39900 16884
rect 39956 16828 41132 16884
rect 41188 16828 41198 16884
rect 42028 16772 42084 17164
rect 49980 17108 50036 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 51100 17164 56476 17220
rect 56532 17164 56542 17220
rect 51100 17108 51156 17164
rect 48850 17052 48860 17108
rect 48916 17052 50036 17108
rect 50194 17052 50204 17108
rect 50260 17052 51156 17108
rect 53778 17052 53788 17108
rect 53844 17052 54572 17108
rect 54628 17052 54638 17108
rect 60162 17052 60172 17108
rect 60228 17052 62188 17108
rect 62244 17052 62254 17108
rect 61964 16996 62020 17052
rect 45826 16940 45836 16996
rect 45892 16940 45902 16996
rect 48738 16940 48748 16996
rect 48804 16940 50204 16996
rect 50260 16940 50270 16996
rect 50418 16940 50428 16996
rect 50484 16940 53340 16996
rect 53396 16940 53406 16996
rect 55906 16940 55916 16996
rect 55972 16940 57596 16996
rect 57652 16940 57662 16996
rect 61954 16940 61964 16996
rect 62020 16940 62030 16996
rect 45836 16884 45892 16940
rect 45836 16828 51996 16884
rect 52052 16828 52062 16884
rect 1362 16716 1372 16772
rect 1428 16716 2268 16772
rect 2324 16716 2334 16772
rect 10098 16716 10108 16772
rect 10164 16716 10332 16772
rect 10388 16716 15372 16772
rect 15428 16716 15438 16772
rect 18386 16716 18396 16772
rect 18452 16716 21868 16772
rect 21924 16716 21934 16772
rect 22754 16716 22764 16772
rect 22820 16716 23996 16772
rect 24052 16716 24062 16772
rect 25554 16716 25564 16772
rect 25620 16716 26796 16772
rect 26852 16716 26862 16772
rect 30146 16716 30156 16772
rect 30212 16716 30828 16772
rect 30884 16716 30894 16772
rect 38882 16716 38892 16772
rect 38948 16716 39228 16772
rect 39284 16716 39294 16772
rect 39666 16716 39676 16772
rect 39732 16716 40684 16772
rect 40740 16716 40750 16772
rect 42028 16716 42476 16772
rect 42532 16716 43876 16772
rect 47702 16716 47740 16772
rect 47796 16716 47806 16772
rect 48626 16716 48636 16772
rect 48692 16716 49756 16772
rect 49812 16716 51436 16772
rect 51492 16716 51502 16772
rect 54450 16716 54460 16772
rect 54516 16716 54908 16772
rect 54964 16716 54974 16772
rect 55458 16716 55468 16772
rect 55524 16716 56140 16772
rect 56196 16716 58380 16772
rect 58436 16716 58446 16772
rect 60610 16716 60620 16772
rect 60676 16716 62524 16772
rect 62580 16716 62590 16772
rect 43820 16660 43876 16716
rect 12002 16604 12012 16660
rect 12068 16604 12908 16660
rect 12964 16604 12974 16660
rect 27570 16604 27580 16660
rect 27636 16604 28252 16660
rect 28308 16604 28318 16660
rect 29698 16604 29708 16660
rect 29764 16604 30716 16660
rect 30772 16604 30782 16660
rect 33618 16604 33628 16660
rect 33684 16604 39452 16660
rect 39508 16604 43596 16660
rect 43652 16604 43662 16660
rect 43820 16604 61852 16660
rect 61908 16604 61918 16660
rect 12002 16492 12012 16548
rect 12068 16492 23548 16548
rect 23604 16492 27468 16548
rect 27524 16492 27534 16548
rect 51538 16492 51548 16548
rect 51604 16492 57652 16548
rect 57810 16492 57820 16548
rect 57876 16492 59836 16548
rect 59892 16492 61516 16548
rect 61572 16492 61582 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 57596 16436 57652 16492
rect 5170 16380 5180 16436
rect 5236 16380 5516 16436
rect 5572 16380 13132 16436
rect 13188 16380 13198 16436
rect 13794 16380 13804 16436
rect 13860 16380 14476 16436
rect 14532 16380 14542 16436
rect 28018 16380 28028 16436
rect 28084 16380 29708 16436
rect 29764 16380 32956 16436
rect 33012 16380 33022 16436
rect 37538 16380 37548 16436
rect 37604 16380 38332 16436
rect 38388 16380 38398 16436
rect 43586 16380 43596 16436
rect 43652 16380 51884 16436
rect 51940 16380 51950 16436
rect 57596 16380 61180 16436
rect 61236 16380 62020 16436
rect 4162 16268 4172 16324
rect 4228 16268 4732 16324
rect 4788 16268 5404 16324
rect 5460 16268 6300 16324
rect 6356 16268 6366 16324
rect 10434 16268 10444 16324
rect 10500 16268 13916 16324
rect 13972 16268 13982 16324
rect 22754 16268 22764 16324
rect 22820 16268 25564 16324
rect 25620 16268 25630 16324
rect 49046 16268 49084 16324
rect 49140 16268 49150 16324
rect 49522 16268 49532 16324
rect 49588 16268 50204 16324
rect 50260 16268 50270 16324
rect 51202 16268 51212 16324
rect 51268 16268 51772 16324
rect 51828 16268 58604 16324
rect 58660 16268 58670 16324
rect 61964 16212 62020 16380
rect 1138 16156 1148 16212
rect 1204 16156 3612 16212
rect 3668 16156 3678 16212
rect 4050 16156 4060 16212
rect 4116 16156 6188 16212
rect 6244 16156 6254 16212
rect 13234 16156 13244 16212
rect 13300 16156 15932 16212
rect 15988 16156 16492 16212
rect 16548 16156 16558 16212
rect 19506 16156 19516 16212
rect 19572 16156 20636 16212
rect 20692 16156 21980 16212
rect 22036 16156 22046 16212
rect 33506 16156 33516 16212
rect 33572 16156 37828 16212
rect 41458 16156 41468 16212
rect 41524 16156 46508 16212
rect 46564 16156 46574 16212
rect 48934 16156 48972 16212
rect 49028 16156 49038 16212
rect 49858 16156 49868 16212
rect 49924 16156 49934 16212
rect 53442 16156 53452 16212
rect 53508 16156 53518 16212
rect 55794 16156 55804 16212
rect 55860 16156 56140 16212
rect 56196 16156 56588 16212
rect 56644 16156 59276 16212
rect 59332 16156 59342 16212
rect 61954 16156 61964 16212
rect 62020 16156 62030 16212
rect 37772 16100 37828 16156
rect 49868 16100 49924 16156
rect 53452 16100 53508 16156
rect 5170 16044 5180 16100
rect 5236 16044 6076 16100
rect 6132 16044 6142 16100
rect 7970 16044 7980 16100
rect 8036 16044 8764 16100
rect 8820 16044 8830 16100
rect 9986 16044 9996 16100
rect 10052 16044 12684 16100
rect 12740 16044 13468 16100
rect 13524 16044 14028 16100
rect 14084 16044 14094 16100
rect 18162 16044 18172 16100
rect 18228 16044 20300 16100
rect 20356 16044 21308 16100
rect 21364 16044 21374 16100
rect 24546 16044 24556 16100
rect 24612 16044 25676 16100
rect 25732 16044 25742 16100
rect 27794 16044 27804 16100
rect 27860 16044 28364 16100
rect 28420 16044 28812 16100
rect 28868 16044 28878 16100
rect 36418 16044 36428 16100
rect 36484 16044 37548 16100
rect 37604 16044 37614 16100
rect 37772 16044 38556 16100
rect 38612 16044 39228 16100
rect 39284 16044 39294 16100
rect 42018 16044 42028 16100
rect 42084 16044 42476 16100
rect 42532 16044 44268 16100
rect 44324 16044 44334 16100
rect 47394 16044 47404 16100
rect 47460 16044 47628 16100
rect 47684 16044 48188 16100
rect 48244 16044 48254 16100
rect 49868 16044 54012 16100
rect 54068 16044 54078 16100
rect 54786 16044 54796 16100
rect 54852 16044 54862 16100
rect 58146 16044 58156 16100
rect 58212 16044 58828 16100
rect 58884 16044 58894 16100
rect 54796 15988 54852 16044
rect 2258 15932 2268 15988
rect 2324 15932 3164 15988
rect 3220 15932 3230 15988
rect 3602 15932 3612 15988
rect 3668 15932 4620 15988
rect 4676 15932 7420 15988
rect 7476 15932 7486 15988
rect 23426 15932 23436 15988
rect 23492 15932 30996 15988
rect 31602 15932 31612 15988
rect 31668 15932 33068 15988
rect 33124 15932 33134 15988
rect 37762 15932 37772 15988
rect 37828 15932 38780 15988
rect 38836 15932 38846 15988
rect 42802 15932 42812 15988
rect 42868 15932 47852 15988
rect 47908 15932 47918 15988
rect 50866 15932 50876 15988
rect 50932 15932 51548 15988
rect 51604 15932 51614 15988
rect 53442 15932 53452 15988
rect 53508 15932 55356 15988
rect 55412 15932 55422 15988
rect 57586 15932 57596 15988
rect 57652 15932 57932 15988
rect 57988 15932 59500 15988
rect 59556 15932 59566 15988
rect 30940 15876 30996 15932
rect 4946 15820 4956 15876
rect 5012 15820 5852 15876
rect 5908 15820 5918 15876
rect 21858 15820 21868 15876
rect 21924 15820 22540 15876
rect 22596 15820 22606 15876
rect 24098 15820 24108 15876
rect 24164 15820 24332 15876
rect 24388 15820 24398 15876
rect 24658 15820 24668 15876
rect 24724 15820 26124 15876
rect 26180 15820 26190 15876
rect 27458 15820 27468 15876
rect 27524 15820 28028 15876
rect 28084 15820 28094 15876
rect 29138 15820 29148 15876
rect 29204 15820 30044 15876
rect 30100 15820 30110 15876
rect 30940 15820 33908 15876
rect 34626 15820 34636 15876
rect 34692 15820 36988 15876
rect 37044 15820 37054 15876
rect 40114 15820 40124 15876
rect 40180 15820 44828 15876
rect 44884 15820 44894 15876
rect 47954 15820 47964 15876
rect 48020 15820 48636 15876
rect 48692 15820 48702 15876
rect 53106 15820 53116 15876
rect 53172 15820 57036 15876
rect 57092 15820 57102 15876
rect 58034 15820 58044 15876
rect 58100 15820 61068 15876
rect 61124 15820 61134 15876
rect 33852 15764 33908 15820
rect 3938 15708 3948 15764
rect 4004 15708 8652 15764
rect 8708 15708 8718 15764
rect 23324 15708 33628 15764
rect 33684 15708 33694 15764
rect 33852 15708 35084 15764
rect 35140 15708 35150 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 23324 15652 23380 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 2706 15596 2716 15652
rect 2772 15596 3836 15652
rect 3892 15596 11900 15652
rect 11956 15596 11966 15652
rect 23314 15596 23324 15652
rect 23380 15596 23390 15652
rect 23986 15596 23996 15652
rect 24052 15596 25116 15652
rect 25172 15596 25182 15652
rect 26852 15596 36428 15652
rect 36484 15596 44268 15652
rect 44324 15596 44334 15652
rect 49298 15596 49308 15652
rect 49364 15596 50092 15652
rect 50148 15596 50158 15652
rect 26852 15540 26908 15596
rect 1250 15484 1260 15540
rect 1316 15484 4284 15540
rect 4340 15484 4350 15540
rect 9314 15484 9324 15540
rect 9380 15484 11788 15540
rect 11844 15484 26908 15540
rect 29698 15484 29708 15540
rect 29764 15484 30716 15540
rect 30772 15484 30782 15540
rect 37650 15484 37660 15540
rect 37716 15484 38108 15540
rect 38164 15484 38174 15540
rect 41794 15484 41804 15540
rect 41860 15484 42588 15540
rect 42644 15484 44268 15540
rect 44324 15484 44334 15540
rect 45490 15484 45500 15540
rect 45556 15484 49588 15540
rect 49532 15428 49588 15484
rect 50372 15484 51212 15540
rect 51268 15484 51278 15540
rect 52770 15484 52780 15540
rect 52836 15484 53620 15540
rect 59042 15484 59052 15540
rect 59108 15484 60396 15540
rect 60452 15484 60844 15540
rect 60900 15484 60910 15540
rect 61366 15484 61404 15540
rect 61460 15484 61470 15540
rect 62178 15484 62188 15540
rect 62244 15484 62636 15540
rect 62692 15484 62702 15540
rect 50372 15428 50428 15484
rect 53564 15428 53620 15484
rect 2706 15372 2716 15428
rect 2772 15372 3388 15428
rect 3444 15372 3454 15428
rect 4722 15372 4732 15428
rect 4788 15372 5516 15428
rect 5572 15372 7308 15428
rect 7364 15372 7374 15428
rect 13794 15372 13804 15428
rect 13860 15372 15708 15428
rect 15764 15372 15774 15428
rect 16258 15372 16268 15428
rect 16324 15372 17388 15428
rect 17444 15372 17454 15428
rect 26002 15372 26012 15428
rect 26068 15372 28700 15428
rect 28756 15372 28766 15428
rect 31490 15372 31500 15428
rect 31556 15372 33180 15428
rect 33236 15372 33246 15428
rect 35252 15372 40964 15428
rect 41682 15372 41692 15428
rect 41748 15372 42924 15428
rect 42980 15372 42990 15428
rect 47058 15372 47068 15428
rect 47124 15372 47852 15428
rect 47908 15372 48748 15428
rect 48804 15372 48814 15428
rect 49522 15372 49532 15428
rect 49588 15372 49598 15428
rect 50082 15372 50092 15428
rect 50148 15372 50428 15428
rect 50978 15372 50988 15428
rect 51044 15372 51548 15428
rect 51604 15372 53116 15428
rect 53172 15372 53182 15428
rect 53554 15372 53564 15428
rect 53620 15372 56364 15428
rect 56420 15372 56430 15428
rect 35252 15316 35308 15372
rect 4834 15260 4844 15316
rect 4900 15260 4910 15316
rect 5282 15260 5292 15316
rect 5348 15260 6076 15316
rect 6132 15260 6142 15316
rect 6402 15260 6412 15316
rect 6468 15260 11452 15316
rect 11508 15260 11518 15316
rect 20514 15260 20524 15316
rect 20580 15260 23436 15316
rect 23492 15260 24332 15316
rect 24388 15260 24398 15316
rect 27906 15260 27916 15316
rect 27972 15260 30492 15316
rect 30548 15260 35308 15316
rect 37538 15260 37548 15316
rect 37604 15260 39004 15316
rect 39060 15260 39070 15316
rect 3378 15148 3388 15204
rect 3444 15148 3948 15204
rect 4004 15148 4014 15204
rect 3714 15036 3724 15092
rect 3780 15036 4284 15092
rect 4340 15036 4350 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 4844 14868 4900 15260
rect 40908 15204 40964 15372
rect 42018 15260 42028 15316
rect 42084 15260 42812 15316
rect 42868 15260 43148 15316
rect 43204 15260 44044 15316
rect 44100 15260 44110 15316
rect 48850 15260 48860 15316
rect 48916 15260 49756 15316
rect 49812 15260 50428 15316
rect 50484 15260 50494 15316
rect 50988 15204 51044 15372
rect 55346 15260 55356 15316
rect 55412 15260 56140 15316
rect 56196 15260 56206 15316
rect 5730 15148 5740 15204
rect 5796 15148 7084 15204
rect 7140 15148 7150 15204
rect 21858 15148 21868 15204
rect 21924 15148 22652 15204
rect 22708 15148 23212 15204
rect 23268 15148 24108 15204
rect 24164 15148 24174 15204
rect 24882 15148 24892 15204
rect 24948 15148 25004 15204
rect 25060 15148 25070 15204
rect 26002 15148 26012 15204
rect 26068 15148 26460 15204
rect 26516 15148 26526 15204
rect 40898 15148 40908 15204
rect 40964 15148 40974 15204
rect 41458 15148 41468 15204
rect 41524 15148 42252 15204
rect 42308 15148 42318 15204
rect 48514 15148 48524 15204
rect 48580 15148 49868 15204
rect 49924 15148 51044 15204
rect 51874 15148 51884 15204
rect 51940 15148 52332 15204
rect 52388 15148 53676 15204
rect 53732 15148 56812 15204
rect 56868 15148 56878 15204
rect 18722 15036 18732 15092
rect 18788 15036 19292 15092
rect 19348 15036 22092 15092
rect 22148 15036 22158 15092
rect 26114 15036 26124 15092
rect 26180 15036 26796 15092
rect 26852 15036 27692 15092
rect 27748 15036 27758 15092
rect 35858 15036 35868 15092
rect 35924 15036 37100 15092
rect 37156 15036 37166 15092
rect 45266 15036 45276 15092
rect 45332 15036 47404 15092
rect 47460 15036 47470 15092
rect 48178 15036 48188 15092
rect 48244 15036 49308 15092
rect 49364 15036 49532 15092
rect 49588 15036 49598 15092
rect 13766 14924 13804 14980
rect 13860 14924 13870 14980
rect 19506 14924 19516 14980
rect 19572 14924 20076 14980
rect 20132 14924 22204 14980
rect 22260 14924 22270 14980
rect 24434 14924 24444 14980
rect 24500 14924 26236 14980
rect 26292 14924 26302 14980
rect 26852 14924 32956 14980
rect 33012 14924 33022 14980
rect 34626 14924 34636 14980
rect 34692 14924 34972 14980
rect 35028 14924 35038 14980
rect 39106 14924 39116 14980
rect 39172 14924 39452 14980
rect 39508 14924 39518 14980
rect 40786 14924 40796 14980
rect 40852 14924 41916 14980
rect 41972 14924 47180 14980
rect 47236 14924 50204 14980
rect 50260 14924 50270 14980
rect 58594 14924 58604 14980
rect 58660 14924 59388 14980
rect 59444 14924 59454 14980
rect 4844 14812 5852 14868
rect 5908 14812 5918 14868
rect 21298 14812 21308 14868
rect 21364 14812 23436 14868
rect 23492 14812 26012 14868
rect 26068 14812 26078 14868
rect 26852 14756 26908 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 40338 14812 40348 14868
rect 40404 14812 47964 14868
rect 48020 14812 48030 14868
rect 49298 14812 49308 14868
rect 49364 14812 49374 14868
rect 49522 14812 49532 14868
rect 49588 14812 49756 14868
rect 49812 14812 49822 14868
rect 49308 14756 49364 14812
rect 3602 14700 3612 14756
rect 3668 14700 13580 14756
rect 13636 14700 14700 14756
rect 14756 14700 14766 14756
rect 18610 14700 18620 14756
rect 18676 14700 26908 14756
rect 27346 14700 27356 14756
rect 27412 14700 29596 14756
rect 29652 14700 30604 14756
rect 30660 14700 30670 14756
rect 31154 14700 31164 14756
rect 31220 14700 33068 14756
rect 33124 14700 33134 14756
rect 33366 14700 33404 14756
rect 33460 14700 33470 14756
rect 33954 14700 33964 14756
rect 34020 14700 34524 14756
rect 34580 14700 35532 14756
rect 35588 14700 35598 14756
rect 37090 14700 37100 14756
rect 37156 14700 40012 14756
rect 40068 14700 40078 14756
rect 42130 14700 42140 14756
rect 42196 14700 43708 14756
rect 43764 14700 44940 14756
rect 44996 14700 45006 14756
rect 49308 14700 50652 14756
rect 50708 14700 50718 14756
rect 56242 14700 56252 14756
rect 56308 14700 58156 14756
rect 58212 14700 58222 14756
rect 61058 14700 61068 14756
rect 61124 14700 62412 14756
rect 62468 14700 62478 14756
rect 2482 14588 2492 14644
rect 2548 14588 4172 14644
rect 4228 14588 4238 14644
rect 6262 14588 6300 14644
rect 6356 14588 6366 14644
rect 6636 14588 14812 14644
rect 14868 14588 14878 14644
rect 27794 14588 27804 14644
rect 27860 14588 29260 14644
rect 29316 14588 31612 14644
rect 31668 14588 31678 14644
rect 39890 14588 39900 14644
rect 39956 14588 40908 14644
rect 40964 14588 43316 14644
rect 6636 14532 6692 14588
rect 43260 14532 43316 14588
rect 55412 14588 58604 14644
rect 58660 14588 61292 14644
rect 61348 14588 61358 14644
rect 61590 14588 61628 14644
rect 61684 14588 61694 14644
rect 3490 14476 3500 14532
rect 3556 14476 6692 14532
rect 6850 14476 6860 14532
rect 6916 14476 7532 14532
rect 7588 14476 7598 14532
rect 11554 14476 11564 14532
rect 11620 14476 14476 14532
rect 14532 14476 14924 14532
rect 14980 14476 14990 14532
rect 15148 14476 17836 14532
rect 17892 14476 17902 14532
rect 20626 14476 20636 14532
rect 20692 14476 21420 14532
rect 21476 14476 21486 14532
rect 23762 14476 23772 14532
rect 23828 14476 25228 14532
rect 25284 14476 25294 14532
rect 25778 14476 25788 14532
rect 25844 14476 28364 14532
rect 28420 14476 28430 14532
rect 29362 14476 29372 14532
rect 29428 14476 32284 14532
rect 32340 14476 32350 14532
rect 34748 14476 35868 14532
rect 35924 14476 35934 14532
rect 37538 14476 37548 14532
rect 37604 14476 38220 14532
rect 38276 14476 39228 14532
rect 39284 14476 39294 14532
rect 42578 14476 42588 14532
rect 42644 14476 43036 14532
rect 43092 14476 43102 14532
rect 43250 14476 43260 14532
rect 43316 14476 53956 14532
rect 15148 14420 15204 14476
rect 34748 14420 34804 14476
rect 53900 14420 53956 14476
rect 55412 14420 55468 14588
rect 58818 14476 58828 14532
rect 58884 14476 60620 14532
rect 60676 14476 60686 14532
rect 5842 14364 5852 14420
rect 5908 14364 9100 14420
rect 9156 14364 9884 14420
rect 9940 14364 9950 14420
rect 11218 14364 11228 14420
rect 11284 14364 12572 14420
rect 12628 14364 12638 14420
rect 13794 14364 13804 14420
rect 13860 14364 14812 14420
rect 14868 14364 15204 14420
rect 15586 14364 15596 14420
rect 15652 14364 16044 14420
rect 16100 14364 16110 14420
rect 18946 14364 18956 14420
rect 19012 14364 22876 14420
rect 22932 14364 22942 14420
rect 23986 14364 23996 14420
rect 24052 14364 26124 14420
rect 26180 14364 26190 14420
rect 26562 14364 26572 14420
rect 26628 14364 27356 14420
rect 27412 14364 27422 14420
rect 30146 14364 30156 14420
rect 30212 14364 33068 14420
rect 33124 14364 33404 14420
rect 33460 14364 33470 14420
rect 34514 14364 34524 14420
rect 34580 14364 34748 14420
rect 34804 14364 34814 14420
rect 34962 14364 34972 14420
rect 35028 14364 36092 14420
rect 36148 14364 36540 14420
rect 36596 14364 36606 14420
rect 38882 14364 38892 14420
rect 38948 14364 39452 14420
rect 39508 14364 39518 14420
rect 41010 14364 41020 14420
rect 41076 14364 41356 14420
rect 41412 14364 43596 14420
rect 43652 14364 43662 14420
rect 46162 14364 46172 14420
rect 46228 14364 46508 14420
rect 46564 14364 47068 14420
rect 47124 14364 47134 14420
rect 49186 14364 49196 14420
rect 49252 14364 49532 14420
rect 49588 14364 49598 14420
rect 53890 14364 53900 14420
rect 53956 14364 53966 14420
rect 55010 14364 55020 14420
rect 55076 14364 55468 14420
rect 57698 14364 57708 14420
rect 57764 14364 61068 14420
rect 61124 14364 61134 14420
rect 2930 14252 2940 14308
rect 2996 14252 3500 14308
rect 3556 14252 4732 14308
rect 4788 14252 4798 14308
rect 5058 14252 5068 14308
rect 5124 14252 9212 14308
rect 9268 14252 9660 14308
rect 9716 14252 9726 14308
rect 15250 14252 15260 14308
rect 15316 14252 16268 14308
rect 16324 14252 17276 14308
rect 17332 14252 17342 14308
rect 18386 14252 18396 14308
rect 18452 14252 20244 14308
rect 21410 14252 21420 14308
rect 21476 14252 25452 14308
rect 25508 14252 25518 14308
rect 28578 14252 28588 14308
rect 28644 14252 29596 14308
rect 29652 14252 29662 14308
rect 30370 14252 30380 14308
rect 30436 14252 31836 14308
rect 31892 14252 34412 14308
rect 34468 14252 37996 14308
rect 38052 14252 38062 14308
rect 41122 14252 41132 14308
rect 41188 14252 42700 14308
rect 42756 14252 42766 14308
rect 46834 14252 46844 14308
rect 46900 14252 47516 14308
rect 47572 14252 47740 14308
rect 47796 14252 47806 14308
rect 53330 14252 53340 14308
rect 53396 14252 55916 14308
rect 55972 14252 58828 14308
rect 20188 14196 20244 14252
rect 41132 14196 41188 14252
rect 5394 14140 5404 14196
rect 5460 14140 5964 14196
rect 6020 14140 15148 14196
rect 18274 14140 18284 14196
rect 18340 14140 18732 14196
rect 18788 14140 18798 14196
rect 20188 14140 25340 14196
rect 25396 14140 25406 14196
rect 34710 14140 34748 14196
rect 34804 14140 34814 14196
rect 35858 14140 35868 14196
rect 35924 14140 36764 14196
rect 36820 14140 38892 14196
rect 38948 14140 38958 14196
rect 39554 14140 39564 14196
rect 39620 14140 41188 14196
rect 51650 14140 51660 14196
rect 51716 14140 52892 14196
rect 52948 14140 56588 14196
rect 56644 14140 56654 14196
rect 5506 14028 5516 14084
rect 5572 14028 11564 14084
rect 11620 14028 12572 14084
rect 12628 14028 12638 14084
rect 15092 13972 15148 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 58772 14084 58828 14252
rect 39564 14028 50428 14084
rect 54002 14028 54012 14084
rect 54068 14028 58492 14084
rect 58548 14028 58558 14084
rect 58772 14028 60340 14084
rect 39564 13972 39620 14028
rect 50372 13972 50428 14028
rect 58492 13972 58548 14028
rect 60284 13972 60340 14028
rect 4610 13916 4620 13972
rect 4676 13916 5852 13972
rect 5908 13916 5918 13972
rect 6178 13916 6188 13972
rect 6244 13916 7196 13972
rect 7252 13916 7262 13972
rect 10210 13916 10220 13972
rect 10276 13916 12236 13972
rect 12292 13916 12302 13972
rect 15092 13916 27244 13972
rect 27300 13916 28140 13972
rect 28196 13916 28206 13972
rect 32274 13916 32284 13972
rect 32340 13916 32732 13972
rect 32788 13916 32798 13972
rect 39554 13916 39564 13972
rect 39620 13916 39630 13972
rect 40338 13916 40348 13972
rect 40404 13916 40414 13972
rect 47506 13916 47516 13972
rect 47572 13916 49084 13972
rect 49140 13916 49150 13972
rect 50372 13916 50652 13972
rect 50708 13916 50718 13972
rect 52098 13916 52108 13972
rect 52164 13916 54012 13972
rect 54068 13916 54078 13972
rect 58492 13916 59612 13972
rect 59668 13916 59678 13972
rect 60274 13916 60284 13972
rect 60340 13916 60350 13972
rect 2370 13804 2380 13860
rect 2436 13804 3388 13860
rect 4050 13804 4060 13860
rect 4116 13804 4844 13860
rect 4900 13804 11004 13860
rect 11060 13804 11070 13860
rect 12450 13804 12460 13860
rect 12516 13804 13132 13860
rect 13188 13804 13198 13860
rect 15810 13804 15820 13860
rect 15876 13804 16940 13860
rect 16996 13804 17006 13860
rect 18610 13804 18620 13860
rect 18676 13804 20636 13860
rect 20692 13804 20702 13860
rect 33394 13804 33404 13860
rect 33460 13804 35420 13860
rect 35476 13804 35486 13860
rect 3332 13748 3388 13804
rect 40348 13748 40404 13916
rect 48066 13804 48076 13860
rect 48132 13804 52332 13860
rect 52388 13804 52398 13860
rect 53788 13804 60732 13860
rect 60788 13804 60798 13860
rect 3332 13692 5516 13748
rect 5572 13692 5582 13748
rect 8978 13692 8988 13748
rect 9044 13692 10668 13748
rect 10724 13692 10734 13748
rect 11666 13692 11676 13748
rect 11732 13692 12684 13748
rect 12740 13692 12750 13748
rect 14578 13692 14588 13748
rect 14644 13692 15036 13748
rect 15092 13692 16380 13748
rect 16436 13692 17612 13748
rect 17668 13692 17678 13748
rect 19058 13692 19068 13748
rect 19124 13692 21420 13748
rect 21476 13692 21486 13748
rect 25554 13692 25564 13748
rect 25620 13692 29932 13748
rect 29988 13692 29998 13748
rect 30902 13692 30940 13748
rect 30996 13692 31006 13748
rect 31714 13692 31724 13748
rect 31780 13692 33292 13748
rect 33348 13692 35196 13748
rect 35252 13692 35262 13748
rect 35970 13692 35980 13748
rect 36036 13692 36876 13748
rect 36932 13692 36942 13748
rect 40348 13692 41132 13748
rect 41188 13692 41198 13748
rect 42690 13692 42700 13748
rect 42756 13692 43708 13748
rect 43764 13692 46060 13748
rect 46116 13692 46126 13748
rect 46722 13692 46732 13748
rect 46788 13692 47628 13748
rect 47684 13692 47694 13748
rect 50082 13692 50092 13748
rect 50148 13692 50428 13748
rect 50484 13692 50494 13748
rect 52546 13692 52556 13748
rect 52612 13692 53340 13748
rect 53396 13692 53406 13748
rect 53788 13636 53844 13804
rect 55346 13692 55356 13748
rect 55412 13692 57148 13748
rect 57204 13692 57214 13748
rect 58146 13692 58156 13748
rect 58212 13692 59836 13748
rect 59892 13692 59902 13748
rect 5170 13580 5180 13636
rect 5236 13580 5628 13636
rect 5684 13580 7084 13636
rect 7140 13580 9436 13636
rect 9492 13580 9502 13636
rect 10444 13580 10892 13636
rect 10948 13580 10958 13636
rect 11106 13580 11116 13636
rect 11172 13580 15596 13636
rect 15652 13580 15662 13636
rect 21522 13580 21532 13636
rect 21588 13580 23660 13636
rect 23716 13580 23726 13636
rect 40002 13580 40012 13636
rect 40068 13580 40796 13636
rect 40852 13580 40862 13636
rect 41346 13580 41356 13636
rect 41412 13580 41916 13636
rect 41972 13580 41982 13636
rect 43026 13580 43036 13636
rect 43092 13580 45276 13636
rect 45332 13580 45342 13636
rect 48962 13580 48972 13636
rect 49028 13580 53844 13636
rect 10444 13524 10500 13580
rect 53788 13524 53844 13580
rect 56364 13580 57596 13636
rect 57652 13580 57662 13636
rect 56364 13524 56420 13580
rect 4722 13468 4732 13524
rect 4788 13468 4900 13524
rect 8754 13468 8764 13524
rect 8820 13468 10444 13524
rect 10500 13468 10510 13524
rect 10770 13468 10780 13524
rect 10836 13468 13692 13524
rect 13748 13468 13758 13524
rect 14354 13468 14364 13524
rect 14420 13468 16380 13524
rect 16436 13468 16446 13524
rect 22194 13468 22204 13524
rect 22260 13468 23100 13524
rect 23156 13468 24668 13524
rect 24724 13468 24734 13524
rect 25442 13468 25452 13524
rect 25508 13468 25788 13524
rect 25844 13468 25854 13524
rect 30034 13468 30044 13524
rect 30100 13468 30716 13524
rect 30772 13468 31164 13524
rect 31220 13468 31230 13524
rect 34850 13468 34860 13524
rect 34916 13468 35644 13524
rect 35700 13468 35710 13524
rect 39526 13468 39564 13524
rect 39620 13468 39630 13524
rect 40226 13468 40236 13524
rect 40292 13468 42588 13524
rect 42644 13468 42654 13524
rect 42802 13468 42812 13524
rect 42868 13468 44492 13524
rect 44548 13468 48300 13524
rect 48356 13468 48366 13524
rect 50166 13468 50204 13524
rect 50260 13468 50270 13524
rect 53778 13468 53788 13524
rect 53844 13468 53854 13524
rect 54002 13468 54012 13524
rect 54068 13468 56420 13524
rect 56578 13468 56588 13524
rect 56644 13468 57932 13524
rect 57988 13468 57998 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 4844 13300 4900 13468
rect 6262 13356 6300 13412
rect 6356 13356 6366 13412
rect 8530 13356 8540 13412
rect 8596 13356 9548 13412
rect 9604 13356 11228 13412
rect 11284 13356 11294 13412
rect 19618 13356 19628 13412
rect 19684 13356 21980 13412
rect 22036 13356 23996 13412
rect 24052 13356 24062 13412
rect 36642 13356 36652 13412
rect 36708 13356 46060 13412
rect 46116 13356 46126 13412
rect 56690 13356 56700 13412
rect 56756 13356 57820 13412
rect 57876 13356 57886 13412
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 4844 13244 6860 13300
rect 6916 13244 8428 13300
rect 8484 13244 8494 13300
rect 19730 13244 19740 13300
rect 19796 13244 21308 13300
rect 21364 13244 21374 13300
rect 22642 13244 22652 13300
rect 22708 13244 22988 13300
rect 23044 13244 25900 13300
rect 25956 13244 25966 13300
rect 30818 13244 30828 13300
rect 30884 13244 31388 13300
rect 31444 13244 31454 13300
rect 48514 13244 48524 13300
rect 48580 13244 58044 13300
rect 58100 13244 58110 13300
rect 22652 13188 22708 13244
rect 1922 13132 1932 13188
rect 1988 13132 2828 13188
rect 2884 13132 15484 13188
rect 15540 13132 15550 13188
rect 20402 13132 20412 13188
rect 20468 13132 22708 13188
rect 22866 13132 22876 13188
rect 22932 13132 23436 13188
rect 23492 13132 23502 13188
rect 24322 13132 24332 13188
rect 24388 13132 43092 13188
rect 43036 13076 43092 13132
rect 47292 13132 56924 13188
rect 56980 13132 56990 13188
rect 2034 13020 2044 13076
rect 2100 13020 3388 13076
rect 3444 13020 4060 13076
rect 4116 13020 4126 13076
rect 5058 13020 5068 13076
rect 5124 13020 8652 13076
rect 8708 13020 9996 13076
rect 10052 13020 10062 13076
rect 17826 13020 17836 13076
rect 17892 13020 21756 13076
rect 21812 13020 21822 13076
rect 30258 13020 30268 13076
rect 30324 13020 30604 13076
rect 30660 13020 30670 13076
rect 37874 13020 37884 13076
rect 37940 13020 38444 13076
rect 38500 13020 38668 13076
rect 38724 13020 38734 13076
rect 40114 13020 40124 13076
rect 40180 13020 40684 13076
rect 40740 13020 40750 13076
rect 43036 13020 47068 13076
rect 47124 13020 47134 13076
rect 47292 12964 47348 13132
rect 48178 13020 48188 13076
rect 48244 13020 49980 13076
rect 50036 13020 50046 13076
rect 53330 13020 53340 13076
rect 53396 13020 54236 13076
rect 54292 13020 55804 13076
rect 55860 13020 55870 13076
rect 57586 13020 57596 13076
rect 57652 13020 58268 13076
rect 58324 13020 59164 13076
rect 59220 13020 59230 13076
rect 3826 12908 3836 12964
rect 3892 12908 9940 12964
rect 14242 12908 14252 12964
rect 14308 12908 16604 12964
rect 16660 12908 16670 12964
rect 21074 12908 21084 12964
rect 21140 12908 22876 12964
rect 22932 12908 23212 12964
rect 23268 12908 23278 12964
rect 24994 12908 25004 12964
rect 25060 12908 25676 12964
rect 25732 12908 25742 12964
rect 31266 12908 31276 12964
rect 31332 12908 31836 12964
rect 31892 12908 31902 12964
rect 34514 12908 34524 12964
rect 34580 12908 35196 12964
rect 35252 12908 35262 12964
rect 39218 12908 39228 12964
rect 39284 12908 40460 12964
rect 40516 12908 41468 12964
rect 41524 12908 41534 12964
rect 43250 12908 43260 12964
rect 43316 12908 47348 12964
rect 50082 12908 50092 12964
rect 50148 12908 50158 12964
rect 54114 12908 54124 12964
rect 54180 12908 55244 12964
rect 55300 12908 55692 12964
rect 55748 12908 55758 12964
rect 9884 12852 9940 12908
rect 50092 12852 50148 12908
rect 6626 12796 6636 12852
rect 6692 12796 7644 12852
rect 7700 12796 8540 12852
rect 8596 12796 8606 12852
rect 9874 12796 9884 12852
rect 9940 12796 14028 12852
rect 14084 12796 14094 12852
rect 16482 12796 16492 12852
rect 16548 12796 17052 12852
rect 17108 12796 17118 12852
rect 19506 12796 19516 12852
rect 19572 12796 21644 12852
rect 21700 12796 21710 12852
rect 29698 12796 29708 12852
rect 29764 12796 30604 12852
rect 30660 12796 32620 12852
rect 32676 12796 34076 12852
rect 34132 12796 35532 12852
rect 35588 12796 35598 12852
rect 40674 12796 40684 12852
rect 40740 12796 40796 12852
rect 40852 12796 40862 12852
rect 44230 12796 44268 12852
rect 44324 12796 44940 12852
rect 44996 12796 45006 12852
rect 48290 12796 48300 12852
rect 48356 12796 49196 12852
rect 49252 12796 49262 12852
rect 50092 12796 50652 12852
rect 50708 12796 50718 12852
rect 56242 12796 56252 12852
rect 56308 12796 59500 12852
rect 59556 12796 59566 12852
rect 4050 12684 4060 12740
rect 4116 12684 5740 12740
rect 5796 12684 7084 12740
rect 7140 12684 7980 12740
rect 8036 12684 8046 12740
rect 18722 12684 18732 12740
rect 18788 12684 20188 12740
rect 20244 12684 20254 12740
rect 20514 12684 20524 12740
rect 20580 12684 21308 12740
rect 21364 12684 21374 12740
rect 22082 12684 22092 12740
rect 22148 12684 22652 12740
rect 22708 12684 22718 12740
rect 26684 12684 26908 12740
rect 26964 12684 26974 12740
rect 27580 12684 28924 12740
rect 28980 12684 28990 12740
rect 29362 12684 29372 12740
rect 29428 12684 31164 12740
rect 31220 12684 34524 12740
rect 34580 12684 34590 12740
rect 39218 12684 39228 12740
rect 39284 12684 48524 12740
rect 48580 12684 48590 12740
rect 50418 12684 50428 12740
rect 50484 12684 53340 12740
rect 53396 12684 53406 12740
rect 54114 12684 54124 12740
rect 54180 12684 55020 12740
rect 55076 12684 55086 12740
rect 22092 12572 23436 12628
rect 23492 12572 26460 12628
rect 26516 12572 26526 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 22092 12516 22148 12572
rect 26684 12516 26740 12684
rect 27580 12628 27636 12684
rect 22082 12460 22092 12516
rect 22148 12460 22158 12516
rect 22428 12460 26740 12516
rect 26852 12572 27356 12628
rect 27412 12572 27636 12628
rect 28690 12572 28700 12628
rect 28756 12572 29148 12628
rect 29204 12572 29932 12628
rect 29988 12572 29998 12628
rect 55682 12572 55692 12628
rect 55748 12572 57148 12628
rect 57204 12572 57214 12628
rect 22428 12404 22484 12460
rect 26852 12404 26908 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 27430 12460 27468 12516
rect 27524 12460 27534 12516
rect 29026 12460 29036 12516
rect 29092 12460 33292 12516
rect 33348 12460 33358 12516
rect 37426 12460 37436 12516
rect 37492 12460 38108 12516
rect 38164 12460 39116 12516
rect 39172 12460 39182 12516
rect 49410 12460 49420 12516
rect 49476 12460 50316 12516
rect 50372 12460 50382 12516
rect 15586 12348 15596 12404
rect 15652 12348 17668 12404
rect 22418 12348 22428 12404
rect 22484 12348 22494 12404
rect 22754 12348 22764 12404
rect 22820 12348 24108 12404
rect 24164 12348 24174 12404
rect 24322 12348 24332 12404
rect 24388 12348 25900 12404
rect 25956 12348 25966 12404
rect 26114 12348 26124 12404
rect 26180 12348 26908 12404
rect 28242 12348 28252 12404
rect 28308 12348 29148 12404
rect 29204 12348 29214 12404
rect 29922 12348 29932 12404
rect 29988 12348 31052 12404
rect 31108 12348 35308 12404
rect 35364 12348 35374 12404
rect 35858 12348 35868 12404
rect 35924 12348 37996 12404
rect 38052 12348 39676 12404
rect 39732 12348 39742 12404
rect 41458 12348 41468 12404
rect 41524 12348 43036 12404
rect 43092 12348 43102 12404
rect 50082 12348 50092 12404
rect 50148 12348 55468 12404
rect 55524 12348 55534 12404
rect 55794 12348 55804 12404
rect 55860 12348 56588 12404
rect 56644 12348 56654 12404
rect 58818 12348 58828 12404
rect 58884 12348 61180 12404
rect 61236 12348 61246 12404
rect 17612 12292 17668 12348
rect 8978 12236 8988 12292
rect 9044 12236 10556 12292
rect 10612 12236 11788 12292
rect 11844 12236 11854 12292
rect 13122 12236 13132 12292
rect 13188 12236 13580 12292
rect 13636 12236 13646 12292
rect 15250 12236 15260 12292
rect 15316 12236 16492 12292
rect 16548 12236 16558 12292
rect 17612 12236 18340 12292
rect 18498 12236 18508 12292
rect 18564 12236 20300 12292
rect 20356 12236 20860 12292
rect 20916 12236 20926 12292
rect 21970 12236 21980 12292
rect 22036 12236 22316 12292
rect 22372 12236 22382 12292
rect 25340 12236 29596 12292
rect 29652 12236 31276 12292
rect 31332 12236 31342 12292
rect 36978 12236 36988 12292
rect 37044 12236 38444 12292
rect 38500 12236 38510 12292
rect 41234 12236 41244 12292
rect 41300 12236 42812 12292
rect 42868 12236 42878 12292
rect 43334 12236 43372 12292
rect 43428 12236 43438 12292
rect 51174 12236 51212 12292
rect 51268 12236 51278 12292
rect 3332 12124 5964 12180
rect 6020 12124 11172 12180
rect 11862 12124 11900 12180
rect 11956 12124 11966 12180
rect 12450 12124 12460 12180
rect 12516 12124 13804 12180
rect 13860 12124 14588 12180
rect 14644 12124 14654 12180
rect 15026 12124 15036 12180
rect 3332 12068 3388 12124
rect 2818 12012 2828 12068
rect 2884 12012 3388 12068
rect 3490 12012 3500 12068
rect 3556 12012 3724 12068
rect 3780 12012 3790 12068
rect 6514 12012 6524 12068
rect 6580 12012 10108 12068
rect 10164 12012 10892 12068
rect 10948 12012 10958 12068
rect 11116 11956 11172 12124
rect 15092 12068 15148 12180
rect 16258 12124 16268 12180
rect 16324 12124 17724 12180
rect 17780 12124 17790 12180
rect 18284 12068 18340 12236
rect 25340 12180 25396 12236
rect 18946 12124 18956 12180
rect 19012 12124 20076 12180
rect 20132 12124 20142 12180
rect 20738 12124 20748 12180
rect 20804 12124 23436 12180
rect 23492 12124 23502 12180
rect 25330 12124 25340 12180
rect 25396 12124 25406 12180
rect 25666 12124 25676 12180
rect 25732 12124 28252 12180
rect 28308 12124 30604 12180
rect 30660 12124 30670 12180
rect 38108 12124 38892 12180
rect 38948 12124 38958 12180
rect 41682 12124 41692 12180
rect 41748 12124 42028 12180
rect 42084 12124 42700 12180
rect 42756 12124 42766 12180
rect 43250 12124 43260 12180
rect 43316 12124 44268 12180
rect 44324 12124 45276 12180
rect 45332 12124 45342 12180
rect 57138 12124 57148 12180
rect 57204 12124 58268 12180
rect 58324 12124 58334 12180
rect 15092 12012 17500 12068
rect 17556 12012 17948 12068
rect 18004 12012 18014 12068
rect 18284 12012 23492 12068
rect 23958 12012 23996 12068
rect 24052 12012 24062 12068
rect 24546 12012 24556 12068
rect 24612 12012 28028 12068
rect 28084 12012 28094 12068
rect 30258 12012 30268 12068
rect 30324 12012 31836 12068
rect 31892 12012 33180 12068
rect 33236 12012 33246 12068
rect 33506 12012 33516 12068
rect 33572 12012 36316 12068
rect 36372 12012 36382 12068
rect 4162 11900 4172 11956
rect 4228 11900 5628 11956
rect 5684 11900 5694 11956
rect 7308 11900 8988 11956
rect 9044 11900 9054 11956
rect 11116 11900 15148 11956
rect 15922 11900 15932 11956
rect 15988 11900 22316 11956
rect 22372 11900 22382 11956
rect 7308 11844 7364 11900
rect 15092 11844 15148 11900
rect 23436 11844 23492 12012
rect 23650 11900 23660 11956
rect 23716 11900 26236 11956
rect 26292 11900 26302 11956
rect 26786 11900 26796 11956
rect 26852 11900 28700 11956
rect 28756 11900 28766 11956
rect 33282 11900 33292 11956
rect 33348 11900 35756 11956
rect 35812 11900 35822 11956
rect 38108 11844 38164 12124
rect 47730 12012 47740 12068
rect 47796 12012 53004 12068
rect 53060 12012 57372 12068
rect 57428 12012 59164 12068
rect 59220 12012 59230 12068
rect 7298 11788 7308 11844
rect 7364 11788 7374 11844
rect 7746 11788 7756 11844
rect 7812 11788 8204 11844
rect 8260 11788 8270 11844
rect 15092 11788 16548 11844
rect 23436 11788 23604 11844
rect 25778 11788 25788 11844
rect 25844 11788 26908 11844
rect 27010 11788 27020 11844
rect 27076 11788 29036 11844
rect 29092 11788 29102 11844
rect 37650 11788 37660 11844
rect 37716 11788 38108 11844
rect 38164 11788 38174 11844
rect 41794 11788 41804 11844
rect 41860 11788 42476 11844
rect 42532 11788 42542 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 8418 11676 8428 11732
rect 8484 11676 9324 11732
rect 9380 11676 9390 11732
rect 10098 11564 10108 11620
rect 10164 11564 12124 11620
rect 12180 11564 12190 11620
rect 12338 11564 12348 11620
rect 12404 11564 12684 11620
rect 12740 11564 12750 11620
rect 14018 11564 14028 11620
rect 14084 11564 15148 11620
rect 15204 11564 15214 11620
rect 0 11508 800 11536
rect 16492 11508 16548 11788
rect 23548 11732 23604 11788
rect 26852 11732 26908 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 16706 11676 16716 11732
rect 16772 11676 17836 11732
rect 17892 11676 20580 11732
rect 22614 11676 22652 11732
rect 22708 11676 22718 11732
rect 23538 11676 23548 11732
rect 23604 11676 23614 11732
rect 26852 11676 27356 11732
rect 27412 11676 29260 11732
rect 29316 11676 29932 11732
rect 29988 11676 29998 11732
rect 38658 11676 38668 11732
rect 38724 11676 59276 11732
rect 59332 11676 59342 11732
rect 20524 11620 20580 11676
rect 16818 11564 16828 11620
rect 16884 11564 17612 11620
rect 17668 11564 17678 11620
rect 20514 11564 20524 11620
rect 20580 11564 20590 11620
rect 23650 11564 23660 11620
rect 23716 11564 23996 11620
rect 24052 11564 24062 11620
rect 28354 11564 28364 11620
rect 28420 11564 30604 11620
rect 30660 11564 30670 11620
rect 30818 11564 30828 11620
rect 30884 11564 41132 11620
rect 41188 11564 41198 11620
rect 0 11452 1708 11508
rect 1764 11452 2492 11508
rect 2548 11452 2558 11508
rect 8194 11452 8204 11508
rect 8260 11452 9884 11508
rect 9940 11452 9950 11508
rect 12534 11452 12572 11508
rect 12628 11452 12638 11508
rect 16492 11452 19348 11508
rect 23090 11452 23100 11508
rect 23156 11452 24332 11508
rect 24388 11452 24398 11508
rect 35074 11452 35084 11508
rect 35140 11452 35868 11508
rect 35924 11452 37212 11508
rect 37268 11452 37278 11508
rect 46806 11452 46844 11508
rect 46900 11452 46910 11508
rect 48066 11452 48076 11508
rect 48132 11452 48748 11508
rect 48804 11452 49420 11508
rect 49476 11452 49486 11508
rect 0 11424 800 11452
rect 6514 11340 6524 11396
rect 6580 11340 8876 11396
rect 8932 11340 8942 11396
rect 12338 11340 12348 11396
rect 12404 11340 13132 11396
rect 13188 11340 13198 11396
rect 13346 11340 13356 11396
rect 13412 11340 13916 11396
rect 13972 11340 13982 11396
rect 16482 11340 16492 11396
rect 16548 11340 17948 11396
rect 18004 11340 18014 11396
rect 19292 11284 19348 11452
rect 19506 11340 19516 11396
rect 19572 11340 20188 11396
rect 20244 11340 21868 11396
rect 21924 11340 22764 11396
rect 22820 11340 22830 11396
rect 25218 11340 25228 11396
rect 25284 11340 25676 11396
rect 25732 11340 25742 11396
rect 26562 11340 26572 11396
rect 26628 11340 29372 11396
rect 29428 11340 29438 11396
rect 41234 11340 41244 11396
rect 41300 11340 43260 11396
rect 43316 11340 43326 11396
rect 47618 11340 47628 11396
rect 47684 11340 48188 11396
rect 48244 11340 48972 11396
rect 49028 11340 49308 11396
rect 49364 11340 50988 11396
rect 51044 11340 51054 11396
rect 51986 11340 51996 11396
rect 52052 11340 53116 11396
rect 53172 11340 53182 11396
rect 4946 11228 4956 11284
rect 5012 11228 5740 11284
rect 5796 11228 6636 11284
rect 6692 11228 6702 11284
rect 13244 11228 18956 11284
rect 19012 11228 19022 11284
rect 19292 11228 23996 11284
rect 24052 11228 24062 11284
rect 28130 11228 28140 11284
rect 28196 11228 29596 11284
rect 29652 11228 29662 11284
rect 44146 11228 44156 11284
rect 44212 11228 44716 11284
rect 44772 11228 45164 11284
rect 45220 11228 45230 11284
rect 47394 11228 47404 11284
rect 47460 11228 48356 11284
rect 13244 11172 13300 11228
rect 48300 11172 48356 11228
rect 5058 11116 5068 11172
rect 5124 11116 6076 11172
rect 6132 11116 7756 11172
rect 7812 11116 7822 11172
rect 11676 11116 13244 11172
rect 13300 11116 13310 11172
rect 16594 11116 16604 11172
rect 16660 11116 20636 11172
rect 20692 11116 20702 11172
rect 23538 11116 23548 11172
rect 23604 11116 24220 11172
rect 24276 11116 25452 11172
rect 25508 11116 25518 11172
rect 26338 11116 26348 11172
rect 26404 11116 31388 11172
rect 31444 11116 31454 11172
rect 33058 11116 33068 11172
rect 33124 11116 33964 11172
rect 34020 11116 34030 11172
rect 38612 11116 47516 11172
rect 47572 11116 47582 11172
rect 48290 11116 48300 11172
rect 48356 11116 48860 11172
rect 48916 11116 48926 11172
rect 49858 11116 49868 11172
rect 49924 11116 51044 11172
rect 51202 11116 51212 11172
rect 51268 11116 52780 11172
rect 52836 11116 52846 11172
rect 11676 11060 11732 11116
rect 38612 11060 38668 11116
rect 50988 11060 51044 11116
rect 11666 11004 11676 11060
rect 11732 11004 11742 11060
rect 13010 11004 13020 11060
rect 13076 11004 13580 11060
rect 13636 11004 13646 11060
rect 18582 11004 18620 11060
rect 18676 11004 18686 11060
rect 20850 11004 20860 11060
rect 20916 11004 21196 11060
rect 21252 11004 21262 11060
rect 22642 11004 22652 11060
rect 22708 11004 38668 11060
rect 40898 11004 40908 11060
rect 40964 11004 47628 11060
rect 47684 11004 50428 11060
rect 50988 11004 51436 11060
rect 51492 11004 52220 11060
rect 52276 11004 52892 11060
rect 52948 11004 54348 11060
rect 54404 11004 54414 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 5954 10892 5964 10948
rect 6020 10892 13244 10948
rect 13300 10892 13310 10948
rect 24098 10892 24108 10948
rect 24164 10892 27804 10948
rect 27860 10892 28588 10948
rect 28644 10892 28654 10948
rect 34962 10892 34972 10948
rect 35028 10892 38668 10948
rect 43474 10892 43484 10948
rect 43540 10892 45948 10948
rect 46004 10892 47852 10948
rect 47908 10892 48524 10948
rect 48580 10892 48860 10948
rect 48916 10892 48926 10948
rect 6402 10780 6412 10836
rect 6468 10780 7756 10836
rect 7812 10780 7822 10836
rect 8306 10780 8316 10836
rect 8372 10780 9436 10836
rect 9492 10780 10220 10836
rect 10276 10780 11004 10836
rect 11060 10780 11070 10836
rect 12450 10780 12460 10836
rect 12516 10780 13020 10836
rect 13076 10780 13086 10836
rect 13682 10780 13692 10836
rect 13748 10780 19460 10836
rect 19618 10780 19628 10836
rect 19684 10780 21868 10836
rect 21924 10780 21934 10836
rect 22082 10780 22092 10836
rect 22148 10780 22876 10836
rect 22932 10780 22942 10836
rect 23986 10780 23996 10836
rect 24052 10780 25228 10836
rect 25284 10780 25294 10836
rect 25890 10780 25900 10836
rect 25956 10780 27356 10836
rect 27412 10780 27422 10836
rect 33506 10780 33516 10836
rect 33572 10780 34860 10836
rect 34916 10780 34926 10836
rect 36754 10780 36764 10836
rect 36820 10780 38220 10836
rect 38276 10780 38286 10836
rect 19404 10724 19460 10780
rect 5842 10668 5852 10724
rect 5908 10668 8540 10724
rect 8596 10668 10780 10724
rect 10836 10668 15148 10724
rect 15204 10668 15214 10724
rect 16146 10668 16156 10724
rect 16212 10668 17612 10724
rect 17668 10668 17678 10724
rect 19404 10668 22372 10724
rect 24770 10668 24780 10724
rect 24836 10668 26572 10724
rect 26628 10668 27020 10724
rect 27076 10668 27916 10724
rect 27972 10668 27982 10724
rect 33394 10668 33404 10724
rect 33460 10668 34188 10724
rect 34244 10668 34254 10724
rect 2034 10556 2044 10612
rect 2100 10556 6860 10612
rect 6916 10556 8988 10612
rect 9044 10556 9054 10612
rect 9650 10556 9660 10612
rect 9716 10556 11676 10612
rect 11732 10556 11742 10612
rect 12450 10556 12460 10612
rect 12516 10556 14476 10612
rect 14532 10556 14542 10612
rect 22316 10500 22372 10668
rect 22530 10556 22540 10612
rect 22596 10556 23548 10612
rect 23604 10556 23614 10612
rect 26674 10556 26684 10612
rect 26740 10556 30716 10612
rect 30772 10556 30782 10612
rect 33170 10556 33180 10612
rect 33236 10556 34076 10612
rect 34132 10556 34972 10612
rect 35028 10556 35038 10612
rect 6626 10444 6636 10500
rect 6692 10444 7084 10500
rect 7140 10444 7150 10500
rect 11218 10444 11228 10500
rect 11284 10444 12236 10500
rect 12292 10444 12302 10500
rect 13122 10444 13132 10500
rect 13188 10444 16044 10500
rect 16100 10444 16110 10500
rect 18274 10444 18284 10500
rect 18340 10444 19292 10500
rect 19348 10444 19358 10500
rect 22316 10444 25676 10500
rect 25732 10444 25742 10500
rect 9762 10332 9772 10388
rect 9828 10332 10220 10388
rect 10276 10332 11900 10388
rect 11956 10332 13580 10388
rect 13636 10332 13646 10388
rect 18722 10332 18732 10388
rect 18788 10332 19516 10388
rect 19572 10332 19582 10388
rect 25442 10332 25452 10388
rect 25508 10332 25900 10388
rect 25956 10332 25966 10388
rect 31238 10332 31276 10388
rect 31332 10332 31342 10388
rect 38612 10276 38668 10892
rect 50372 10836 50428 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 40562 10780 40572 10836
rect 40628 10780 43596 10836
rect 43652 10780 43662 10836
rect 46386 10780 46396 10836
rect 46452 10780 47404 10836
rect 47460 10780 48188 10836
rect 48244 10780 48254 10836
rect 50372 10780 57148 10836
rect 57204 10780 57214 10836
rect 43596 10724 43652 10780
rect 43596 10668 47964 10724
rect 48020 10668 48030 10724
rect 41346 10556 41356 10612
rect 41412 10556 42140 10612
rect 42196 10556 42206 10612
rect 47282 10556 47292 10612
rect 47348 10556 48972 10612
rect 49028 10556 49038 10612
rect 49522 10556 49532 10612
rect 49588 10556 50652 10612
rect 50708 10556 52444 10612
rect 52500 10556 52510 10612
rect 52770 10556 52780 10612
rect 52836 10556 54124 10612
rect 54180 10556 54190 10612
rect 48972 10500 49028 10556
rect 48972 10444 49420 10500
rect 49476 10444 49486 10500
rect 49298 10332 49308 10388
rect 49364 10332 52556 10388
rect 52612 10332 52622 10388
rect 12114 10220 12124 10276
rect 12180 10220 13020 10276
rect 13076 10220 13086 10276
rect 17042 10220 17052 10276
rect 17108 10220 17500 10276
rect 17556 10220 19740 10276
rect 19796 10220 21308 10276
rect 21364 10220 21374 10276
rect 23538 10220 23548 10276
rect 23604 10220 24220 10276
rect 24276 10220 24286 10276
rect 27346 10220 27356 10276
rect 27412 10220 27916 10276
rect 27972 10220 27982 10276
rect 38612 10220 50428 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 7298 10108 7308 10164
rect 7364 10108 11788 10164
rect 11844 10108 13804 10164
rect 13860 10108 13870 10164
rect 18610 10108 18620 10164
rect 18676 10108 32788 10164
rect 36866 10108 36876 10164
rect 36932 10108 44604 10164
rect 44660 10108 44670 10164
rect 50372 10108 50428 10220
rect 50484 10108 50494 10164
rect 32732 10052 32788 10108
rect 11554 9996 11564 10052
rect 11620 9996 15484 10052
rect 15540 9996 15550 10052
rect 16482 9996 16492 10052
rect 16548 9996 16558 10052
rect 16930 9996 16940 10052
rect 16996 9996 18956 10052
rect 19012 9996 19022 10052
rect 20290 9996 20300 10052
rect 20356 9996 22876 10052
rect 22932 9996 22942 10052
rect 25218 9996 25228 10052
rect 25284 9996 26796 10052
rect 26852 9996 26862 10052
rect 28578 9996 28588 10052
rect 28644 9996 30492 10052
rect 30548 9996 31276 10052
rect 31332 9996 31342 10052
rect 32732 9996 38668 10052
rect 40338 9996 40348 10052
rect 40404 9996 42252 10052
rect 42308 9996 42318 10052
rect 43586 9996 43596 10052
rect 43652 9996 47404 10052
rect 47460 9996 47470 10052
rect 16492 9940 16548 9996
rect 9986 9884 9996 9940
rect 10052 9884 12796 9940
rect 12852 9884 12862 9940
rect 14690 9884 14700 9940
rect 14756 9884 16548 9940
rect 16604 9884 26236 9940
rect 26292 9884 26302 9940
rect 31350 9884 31388 9940
rect 31444 9884 31454 9940
rect 15026 9772 15036 9828
rect 15092 9772 16380 9828
rect 16436 9772 16446 9828
rect 16604 9716 16660 9884
rect 38612 9828 38668 9996
rect 39862 9884 39900 9940
rect 39956 9884 39966 9940
rect 40674 9884 40684 9940
rect 40740 9884 43260 9940
rect 43316 9884 43326 9940
rect 16930 9772 16940 9828
rect 16996 9772 18060 9828
rect 18116 9772 19292 9828
rect 19348 9772 19358 9828
rect 20626 9772 20636 9828
rect 20692 9772 23212 9828
rect 23268 9772 23278 9828
rect 28242 9772 28252 9828
rect 28308 9772 29372 9828
rect 29428 9772 29438 9828
rect 31938 9772 31948 9828
rect 32004 9772 33292 9828
rect 33348 9772 33358 9828
rect 33954 9772 33964 9828
rect 34020 9772 34524 9828
rect 34580 9772 34590 9828
rect 36082 9772 36092 9828
rect 36148 9772 36540 9828
rect 36596 9772 37212 9828
rect 37268 9772 37278 9828
rect 38612 9772 41580 9828
rect 41636 9772 42700 9828
rect 42756 9772 43148 9828
rect 43204 9772 43214 9828
rect 44258 9772 44268 9828
rect 44324 9772 45388 9828
rect 45444 9772 45454 9828
rect 51762 9772 51772 9828
rect 51828 9772 51996 9828
rect 52052 9772 52780 9828
rect 52836 9772 52846 9828
rect 9314 9660 9324 9716
rect 9380 9660 9884 9716
rect 9940 9660 16660 9716
rect 20402 9660 20412 9716
rect 20468 9660 21420 9716
rect 21476 9660 21486 9716
rect 21634 9660 21644 9716
rect 21700 9660 21980 9716
rect 22036 9660 22046 9716
rect 22204 9660 23436 9716
rect 23492 9660 23502 9716
rect 25778 9660 25788 9716
rect 25844 9660 26796 9716
rect 26852 9660 26862 9716
rect 28354 9660 28364 9716
rect 28420 9660 29932 9716
rect 29988 9660 29998 9716
rect 33404 9660 35980 9716
rect 36036 9660 36046 9716
rect 41346 9660 41356 9716
rect 41412 9660 42476 9716
rect 42532 9660 42542 9716
rect 46946 9660 46956 9716
rect 47012 9660 48860 9716
rect 48916 9660 48926 9716
rect 50866 9660 50876 9716
rect 50932 9660 51660 9716
rect 51716 9660 51726 9716
rect 22204 9604 22260 9660
rect 33404 9604 33460 9660
rect 8306 9548 8316 9604
rect 8372 9548 9548 9604
rect 9604 9548 9614 9604
rect 14354 9548 14364 9604
rect 14420 9548 15148 9604
rect 17154 9548 17164 9604
rect 17220 9548 19740 9604
rect 19796 9548 20300 9604
rect 20356 9548 22260 9604
rect 32498 9548 32508 9604
rect 32564 9548 33404 9604
rect 33460 9548 33470 9604
rect 35522 9548 35532 9604
rect 35588 9548 38668 9604
rect 38724 9548 38734 9604
rect 39666 9548 39676 9604
rect 39732 9548 39788 9604
rect 39844 9548 39854 9604
rect 41458 9548 41468 9604
rect 41524 9548 42588 9604
rect 42644 9548 42654 9604
rect 45826 9548 45836 9604
rect 45892 9548 46620 9604
rect 46676 9548 46686 9604
rect 15092 9492 15148 9548
rect 39788 9492 39844 9548
rect 15092 9436 15708 9492
rect 15764 9436 15774 9492
rect 23314 9436 23324 9492
rect 23380 9436 24332 9492
rect 24388 9436 29708 9492
rect 29764 9436 29774 9492
rect 39788 9436 42812 9492
rect 42868 9436 42878 9492
rect 46722 9436 46732 9492
rect 46788 9436 46798 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 28812 9324 30268 9380
rect 30324 9324 31276 9380
rect 31332 9324 31342 9380
rect 38612 9324 38892 9380
rect 38948 9324 38958 9380
rect 28812 9268 28868 9324
rect 6738 9212 6748 9268
rect 6804 9212 12012 9268
rect 12068 9212 12078 9268
rect 13010 9212 13020 9268
rect 13076 9212 14252 9268
rect 14308 9212 14318 9268
rect 18050 9212 18060 9268
rect 18116 9212 20860 9268
rect 20916 9212 20926 9268
rect 24098 9212 24108 9268
rect 24164 9212 25900 9268
rect 25956 9212 25966 9268
rect 26786 9212 26796 9268
rect 26852 9212 28812 9268
rect 28868 9212 28878 9268
rect 29250 9212 29260 9268
rect 29316 9212 29820 9268
rect 29876 9212 31612 9268
rect 31668 9212 31678 9268
rect 38612 9156 38668 9324
rect 40114 9212 40124 9268
rect 40180 9212 42364 9268
rect 42420 9212 42430 9268
rect 43558 9212 43596 9268
rect 43652 9212 43662 9268
rect 44594 9212 44604 9268
rect 44660 9212 45276 9268
rect 45332 9212 46060 9268
rect 46116 9212 46126 9268
rect 46732 9156 46788 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 53330 9212 53340 9268
rect 53396 9212 54460 9268
rect 54516 9212 54526 9268
rect 8866 9100 8876 9156
rect 8932 9100 14812 9156
rect 14868 9100 14878 9156
rect 18834 9100 18844 9156
rect 18900 9100 20412 9156
rect 20468 9100 20478 9156
rect 24994 9100 25004 9156
rect 25060 9100 28028 9156
rect 28084 9100 28094 9156
rect 32386 9100 32396 9156
rect 32452 9100 32956 9156
rect 33012 9100 33852 9156
rect 33908 9100 34972 9156
rect 35028 9100 35038 9156
rect 35634 9100 35644 9156
rect 35700 9100 36988 9156
rect 37044 9100 37054 9156
rect 37538 9100 37548 9156
rect 37604 9100 38668 9156
rect 38770 9100 38780 9156
rect 38836 9100 39564 9156
rect 39620 9100 39630 9156
rect 45490 9100 45500 9156
rect 45556 9100 47180 9156
rect 47236 9100 47246 9156
rect 8754 8988 8764 9044
rect 8820 8988 10220 9044
rect 10276 8988 10286 9044
rect 19058 8988 19068 9044
rect 19124 8988 19740 9044
rect 19796 8988 19806 9044
rect 19954 8988 19964 9044
rect 20020 8988 20636 9044
rect 20692 8988 21084 9044
rect 21140 8988 21150 9044
rect 26562 8988 26572 9044
rect 26628 8988 28700 9044
rect 28756 8988 28766 9044
rect 32274 8988 32284 9044
rect 32340 8988 32508 9044
rect 32564 8988 33964 9044
rect 34020 8988 34030 9044
rect 34738 8988 34748 9044
rect 34804 8988 35532 9044
rect 35588 8988 35598 9044
rect 35746 8988 35756 9044
rect 35812 8988 36092 9044
rect 36148 8988 37772 9044
rect 37828 8988 37838 9044
rect 38612 8988 39340 9044
rect 39396 8988 39900 9044
rect 39956 8988 39966 9044
rect 40114 8988 40124 9044
rect 40180 8988 41020 9044
rect 41076 8988 41086 9044
rect 42354 8988 42364 9044
rect 42420 8988 43820 9044
rect 43876 8988 43886 9044
rect 45154 8988 45164 9044
rect 45220 8988 45612 9044
rect 45668 8988 46732 9044
rect 46788 8988 46798 9044
rect 46946 8988 46956 9044
rect 47012 8988 47964 9044
rect 48020 8988 48748 9044
rect 48804 8988 48814 9044
rect 51538 8988 51548 9044
rect 51604 8988 52668 9044
rect 52724 8988 52734 9044
rect 38612 8932 38668 8988
rect 7074 8876 7084 8932
rect 7140 8876 10444 8932
rect 10500 8876 11564 8932
rect 11620 8876 11630 8932
rect 16146 8876 16156 8932
rect 16212 8876 16492 8932
rect 16548 8876 16558 8932
rect 20738 8876 20748 8932
rect 20804 8876 21756 8932
rect 21812 8876 21822 8932
rect 22530 8876 22540 8932
rect 22596 8876 23324 8932
rect 23380 8876 23390 8932
rect 27654 8876 27692 8932
rect 27748 8876 27758 8932
rect 28130 8876 28140 8932
rect 28196 8876 30268 8932
rect 30324 8876 30334 8932
rect 33618 8876 33628 8932
rect 33684 8876 33694 8932
rect 34850 8876 34860 8932
rect 34916 8876 38668 8932
rect 39554 8876 39564 8932
rect 39620 8876 41580 8932
rect 41636 8876 44940 8932
rect 44996 8876 45006 8932
rect 47842 8876 47852 8932
rect 47908 8876 49644 8932
rect 49700 8876 49710 8932
rect 25890 8764 25900 8820
rect 25956 8764 31164 8820
rect 31220 8764 31230 8820
rect 31910 8764 31948 8820
rect 32004 8764 32014 8820
rect 33628 8708 33684 8876
rect 35410 8764 35420 8820
rect 35476 8764 37548 8820
rect 37604 8764 37614 8820
rect 38658 8764 38668 8820
rect 38724 8764 39900 8820
rect 39956 8764 39966 8820
rect 44034 8764 44044 8820
rect 44100 8764 45052 8820
rect 45108 8764 45118 8820
rect 46508 8764 53676 8820
rect 53732 8764 53742 8820
rect 46508 8708 46564 8764
rect 15250 8652 15260 8708
rect 15316 8652 16492 8708
rect 16548 8652 33684 8708
rect 38994 8652 39004 8708
rect 39060 8652 43708 8708
rect 43764 8652 43774 8708
rect 43922 8652 43932 8708
rect 43988 8652 44940 8708
rect 44996 8652 46564 8708
rect 50372 8652 55020 8708
rect 55076 8652 55086 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 50372 8596 50428 8652
rect 7970 8540 7980 8596
rect 8036 8540 8540 8596
rect 8596 8540 8606 8596
rect 15698 8540 15708 8596
rect 15764 8540 18620 8596
rect 18676 8540 18686 8596
rect 20178 8540 20188 8596
rect 20244 8540 20468 8596
rect 21410 8540 21420 8596
rect 21476 8540 22428 8596
rect 22484 8540 22494 8596
rect 26338 8540 26348 8596
rect 26404 8540 26908 8596
rect 28018 8540 28028 8596
rect 28084 8540 29260 8596
rect 29316 8540 29326 8596
rect 39890 8540 39900 8596
rect 39956 8540 40012 8596
rect 40068 8540 40078 8596
rect 43138 8540 43148 8596
rect 43204 8540 46060 8596
rect 46116 8540 50428 8596
rect 54562 8540 54572 8596
rect 54628 8540 55916 8596
rect 55972 8540 55982 8596
rect 20412 8372 20468 8540
rect 26852 8484 26908 8540
rect 20626 8428 20636 8484
rect 20692 8428 21644 8484
rect 21700 8428 21710 8484
rect 26852 8428 28252 8484
rect 28308 8428 28318 8484
rect 32162 8428 32172 8484
rect 32228 8428 32508 8484
rect 32564 8428 32574 8484
rect 35410 8428 35420 8484
rect 35476 8428 37100 8484
rect 37156 8428 37166 8484
rect 45042 8428 45052 8484
rect 45108 8428 45556 8484
rect 47730 8428 47740 8484
rect 47796 8428 48748 8484
rect 48804 8428 48814 8484
rect 45500 8372 45556 8428
rect 12534 8316 12572 8372
rect 12628 8316 12638 8372
rect 14130 8316 14140 8372
rect 14196 8316 15260 8372
rect 15316 8316 15326 8372
rect 15820 8316 16380 8372
rect 16436 8316 16446 8372
rect 16706 8316 16716 8372
rect 16772 8316 17948 8372
rect 18004 8316 18014 8372
rect 20402 8316 20412 8372
rect 20468 8316 20478 8372
rect 22978 8316 22988 8372
rect 23044 8316 24220 8372
rect 24276 8316 24286 8372
rect 32722 8316 32732 8372
rect 32788 8316 34412 8372
rect 34468 8316 37212 8372
rect 37268 8316 37278 8372
rect 45500 8316 45612 8372
rect 45668 8316 45678 8372
rect 51986 8316 51996 8372
rect 52052 8316 53004 8372
rect 53060 8316 53070 8372
rect 15820 8260 15876 8316
rect 10994 8204 11004 8260
rect 11060 8204 11564 8260
rect 11620 8204 12460 8260
rect 12516 8204 12526 8260
rect 12786 8204 12796 8260
rect 12852 8204 15876 8260
rect 16034 8204 16044 8260
rect 16100 8204 17388 8260
rect 17444 8204 17454 8260
rect 24434 8204 24444 8260
rect 24500 8204 24780 8260
rect 24836 8204 25116 8260
rect 25172 8204 27356 8260
rect 27412 8204 27422 8260
rect 31378 8204 31388 8260
rect 31444 8204 35980 8260
rect 36036 8204 37996 8260
rect 38052 8204 38062 8260
rect 48850 8204 48860 8260
rect 48916 8204 49420 8260
rect 49476 8204 49486 8260
rect 9538 8092 9548 8148
rect 9604 8092 10892 8148
rect 10948 8092 10958 8148
rect 24658 8092 24668 8148
rect 24724 8092 27132 8148
rect 27188 8092 27198 8148
rect 28690 8092 28700 8148
rect 28756 8092 29708 8148
rect 29764 8092 29774 8148
rect 32946 8092 32956 8148
rect 33012 8092 34636 8148
rect 34692 8092 34702 8148
rect 36082 8092 36092 8148
rect 36148 8092 39004 8148
rect 39060 8092 39070 8148
rect 49298 8092 49308 8148
rect 49364 8092 50428 8148
rect 50484 8092 50494 8148
rect 14802 7980 14812 8036
rect 14868 7980 15932 8036
rect 15988 7980 15998 8036
rect 26114 7980 26124 8036
rect 26180 7980 26572 8036
rect 26628 7980 26638 8036
rect 27682 7980 27692 8036
rect 27748 7980 27804 8036
rect 27860 7980 27870 8036
rect 28466 7980 28476 8036
rect 28532 7980 30828 8036
rect 30884 7980 30894 8036
rect 31490 7980 31500 8036
rect 31556 7980 33628 8036
rect 33684 7980 33694 8036
rect 35858 7980 35868 8036
rect 35924 7980 39228 8036
rect 39284 7980 39294 8036
rect 41346 7980 41356 8036
rect 41412 7980 42140 8036
rect 42196 7980 42812 8036
rect 42868 7980 42878 8036
rect 47012 7980 49196 8036
rect 49252 7980 49262 8036
rect 50372 7980 51660 8036
rect 51716 7980 51726 8036
rect 54114 7980 54124 8036
rect 54180 7980 56700 8036
rect 56756 7980 56766 8036
rect 47012 7924 47068 7980
rect 45714 7868 45724 7924
rect 45780 7868 47068 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50372 7812 50428 7980
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 26562 7756 26572 7812
rect 26628 7756 29148 7812
rect 29204 7756 29214 7812
rect 44146 7756 44156 7812
rect 44212 7756 44492 7812
rect 44548 7756 44558 7812
rect 49186 7756 49196 7812
rect 49252 7756 50428 7812
rect 17378 7644 17388 7700
rect 17444 7644 17612 7700
rect 17668 7644 17678 7700
rect 18722 7644 18732 7700
rect 18788 7644 21196 7700
rect 21252 7644 21262 7700
rect 27794 7644 27804 7700
rect 27860 7644 27870 7700
rect 28354 7644 28364 7700
rect 28420 7644 29932 7700
rect 29988 7644 29998 7700
rect 51650 7644 51660 7700
rect 51716 7644 54012 7700
rect 54068 7644 54078 7700
rect 27804 7588 27860 7644
rect 20290 7532 20300 7588
rect 20356 7532 21084 7588
rect 21140 7532 21150 7588
rect 22866 7532 22876 7588
rect 22932 7532 23436 7588
rect 23492 7532 24108 7588
rect 24164 7532 26908 7588
rect 27804 7532 28476 7588
rect 28532 7532 28542 7588
rect 33842 7532 33852 7588
rect 33908 7532 35420 7588
rect 35476 7532 35486 7588
rect 35746 7532 35756 7588
rect 35812 7532 39340 7588
rect 39396 7532 39406 7588
rect 41906 7532 41916 7588
rect 41972 7532 42924 7588
rect 42980 7532 42990 7588
rect 43362 7532 43372 7588
rect 43428 7532 44492 7588
rect 44548 7532 44558 7588
rect 47954 7532 47964 7588
rect 48020 7532 49980 7588
rect 50036 7532 50046 7588
rect 15250 7420 15260 7476
rect 15316 7420 15932 7476
rect 15988 7420 15998 7476
rect 22418 7420 22428 7476
rect 22484 7420 23660 7476
rect 23716 7420 24556 7476
rect 24612 7420 24622 7476
rect 11666 7308 11676 7364
rect 11732 7308 25564 7364
rect 25620 7308 25630 7364
rect 26852 7252 26908 7532
rect 29362 7420 29372 7476
rect 29428 7420 30492 7476
rect 30548 7420 30558 7476
rect 33506 7420 33516 7476
rect 33572 7420 36092 7476
rect 36148 7420 36158 7476
rect 36306 7420 36316 7476
rect 36372 7420 38220 7476
rect 38276 7420 38286 7476
rect 39778 7420 39788 7476
rect 39844 7420 41244 7476
rect 41300 7420 41310 7476
rect 43474 7420 43484 7476
rect 43540 7420 44156 7476
rect 44212 7420 44222 7476
rect 45602 7420 45612 7476
rect 45668 7420 47404 7476
rect 47460 7420 47470 7476
rect 51090 7420 51100 7476
rect 51156 7420 54124 7476
rect 54180 7420 54190 7476
rect 30258 7308 30268 7364
rect 30324 7308 33180 7364
rect 33236 7308 33246 7364
rect 34738 7308 34748 7364
rect 34804 7308 35644 7364
rect 35700 7308 35710 7364
rect 41906 7308 41916 7364
rect 41972 7308 42700 7364
rect 42756 7308 47740 7364
rect 47796 7308 47806 7364
rect 48178 7308 48188 7364
rect 48244 7308 48860 7364
rect 48916 7308 48926 7364
rect 50194 7308 50204 7364
rect 50260 7308 52444 7364
rect 52500 7308 52510 7364
rect 26852 7196 35588 7252
rect 37426 7196 37436 7252
rect 37492 7196 39788 7252
rect 39844 7196 39854 7252
rect 40114 7196 40124 7252
rect 40180 7196 41020 7252
rect 41076 7196 41086 7252
rect 35532 7140 35588 7196
rect 41916 7140 41972 7308
rect 46162 7196 46172 7252
rect 46228 7196 47516 7252
rect 47572 7196 47582 7252
rect 17490 7084 17500 7140
rect 17556 7084 20188 7140
rect 20244 7084 20254 7140
rect 28466 7084 28476 7140
rect 28532 7084 33852 7140
rect 33908 7084 33918 7140
rect 35532 7084 41972 7140
rect 46610 7084 46620 7140
rect 46676 7084 51212 7140
rect 51268 7084 51278 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 14690 6972 14700 7028
rect 14756 6972 15596 7028
rect 15652 6972 15662 7028
rect 24658 6972 24668 7028
rect 24724 6972 27692 7028
rect 27748 6972 27758 7028
rect 32162 6972 32172 7028
rect 32228 6972 32620 7028
rect 32676 6972 32686 7028
rect 39330 6972 39340 7028
rect 39396 6972 45220 7028
rect 45378 6972 45388 7028
rect 45444 6972 46172 7028
rect 46228 6972 46238 7028
rect 49298 6972 49308 7028
rect 49364 6972 51660 7028
rect 51716 6972 52892 7028
rect 52948 6972 52958 7028
rect 45164 6916 45220 6972
rect 27010 6860 27020 6916
rect 27076 6860 30268 6916
rect 30324 6860 30334 6916
rect 30482 6860 30492 6916
rect 30548 6860 31612 6916
rect 31668 6860 31678 6916
rect 32498 6860 32508 6916
rect 32564 6860 33292 6916
rect 33348 6860 33964 6916
rect 34020 6860 34030 6916
rect 42466 6860 42476 6916
rect 42532 6860 43596 6916
rect 43652 6860 43662 6916
rect 45164 6860 45500 6916
rect 45556 6860 45566 6916
rect 46274 6860 46284 6916
rect 46340 6860 48412 6916
rect 48468 6860 48478 6916
rect 10882 6748 10892 6804
rect 10948 6748 11788 6804
rect 11844 6748 13580 6804
rect 13636 6748 13646 6804
rect 20066 6748 20076 6804
rect 20132 6748 20860 6804
rect 20916 6748 22204 6804
rect 22260 6748 22270 6804
rect 29810 6748 29820 6804
rect 29876 6748 30940 6804
rect 30996 6748 31006 6804
rect 31836 6748 31948 6804
rect 32004 6748 32014 6804
rect 37874 6748 37884 6804
rect 37940 6748 39340 6804
rect 39396 6748 39406 6804
rect 39666 6748 39676 6804
rect 39732 6748 40460 6804
rect 40516 6748 40526 6804
rect 44146 6748 44156 6804
rect 44212 6748 45948 6804
rect 46004 6748 47852 6804
rect 47908 6748 47918 6804
rect 31836 6692 31892 6748
rect 11666 6636 11676 6692
rect 11732 6636 12236 6692
rect 12292 6636 13468 6692
rect 13524 6636 13534 6692
rect 14578 6636 14588 6692
rect 14644 6636 15820 6692
rect 15876 6636 15886 6692
rect 16258 6636 16268 6692
rect 16324 6636 17836 6692
rect 17892 6636 18956 6692
rect 19012 6636 19022 6692
rect 21634 6636 21644 6692
rect 21700 6636 22988 6692
rect 23044 6636 23054 6692
rect 23510 6636 23548 6692
rect 23604 6636 23614 6692
rect 24322 6636 24332 6692
rect 24388 6636 24892 6692
rect 24948 6636 24958 6692
rect 27234 6636 27244 6692
rect 27300 6636 27692 6692
rect 27748 6636 27758 6692
rect 28130 6636 28140 6692
rect 28196 6636 31892 6692
rect 32050 6636 32060 6692
rect 32116 6636 32956 6692
rect 33012 6636 35196 6692
rect 35252 6636 35262 6692
rect 40226 6636 40236 6692
rect 40292 6636 40572 6692
rect 40628 6636 40638 6692
rect 43250 6636 43260 6692
rect 43316 6636 45276 6692
rect 45332 6636 45342 6692
rect 45714 6636 45724 6692
rect 45780 6636 46508 6692
rect 46564 6636 46574 6692
rect 47730 6636 47740 6692
rect 47796 6636 50764 6692
rect 50820 6636 50830 6692
rect 45724 6580 45780 6636
rect 12786 6524 12796 6580
rect 12852 6524 13804 6580
rect 13860 6524 13870 6580
rect 14914 6524 14924 6580
rect 14980 6524 15372 6580
rect 15428 6524 15438 6580
rect 19618 6524 19628 6580
rect 19684 6524 20412 6580
rect 20468 6524 21980 6580
rect 22036 6524 22046 6580
rect 22306 6524 22316 6580
rect 22372 6524 25004 6580
rect 25060 6524 25070 6580
rect 25666 6524 25676 6580
rect 25732 6524 26348 6580
rect 26404 6524 26796 6580
rect 26852 6524 26862 6580
rect 28466 6524 28476 6580
rect 28532 6524 29596 6580
rect 29652 6524 29662 6580
rect 34514 6524 34524 6580
rect 34580 6524 35308 6580
rect 35364 6524 35374 6580
rect 36978 6524 36988 6580
rect 37044 6524 39228 6580
rect 39284 6524 39294 6580
rect 41010 6524 41020 6580
rect 41076 6524 42700 6580
rect 42756 6524 42766 6580
rect 44258 6524 44268 6580
rect 44324 6524 45780 6580
rect 17490 6412 17500 6468
rect 17556 6412 22204 6468
rect 22260 6412 22270 6468
rect 23202 6412 23212 6468
rect 23268 6412 23548 6468
rect 23604 6412 24668 6468
rect 24724 6412 24734 6468
rect 24882 6412 24892 6468
rect 24948 6412 25452 6468
rect 25508 6412 25518 6468
rect 27570 6412 27580 6468
rect 27636 6412 28812 6468
rect 28868 6412 28878 6468
rect 31266 6412 31276 6468
rect 31332 6412 31948 6468
rect 32004 6412 32014 6468
rect 33618 6412 33628 6468
rect 33684 6412 34972 6468
rect 35028 6412 35756 6468
rect 35812 6412 43260 6468
rect 43316 6412 43326 6468
rect 49074 6412 49084 6468
rect 49140 6412 49532 6468
rect 49588 6412 49598 6468
rect 24892 6356 24948 6412
rect 20822 6300 20860 6356
rect 20916 6300 20926 6356
rect 21074 6300 21084 6356
rect 21140 6300 22092 6356
rect 22148 6300 23436 6356
rect 23492 6300 23502 6356
rect 23762 6300 23772 6356
rect 23828 6300 24948 6356
rect 27234 6300 27244 6356
rect 27300 6300 30044 6356
rect 30100 6300 31724 6356
rect 31780 6300 31790 6356
rect 34290 6300 34300 6356
rect 34356 6300 35980 6356
rect 36036 6300 36316 6356
rect 36372 6300 36382 6356
rect 40562 6300 40572 6356
rect 40628 6300 45052 6356
rect 45108 6300 45118 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 21858 6188 21868 6244
rect 21924 6188 23436 6244
rect 23492 6188 25340 6244
rect 25396 6188 25406 6244
rect 25554 6188 25564 6244
rect 25620 6188 26684 6244
rect 26740 6188 31388 6244
rect 31444 6188 31454 6244
rect 32610 6188 32620 6244
rect 32676 6188 33516 6244
rect 33572 6188 33582 6244
rect 43708 6188 47292 6244
rect 47348 6188 49420 6244
rect 49476 6188 49486 6244
rect 43708 6132 43764 6188
rect 49420 6132 49476 6188
rect 16034 6076 16044 6132
rect 16100 6076 16492 6132
rect 16548 6076 16828 6132
rect 16884 6076 16894 6132
rect 20934 6076 20972 6132
rect 21028 6076 21420 6132
rect 21476 6076 21486 6132
rect 21634 6076 21644 6132
rect 21700 6076 21756 6132
rect 21812 6076 21980 6132
rect 22036 6076 22046 6132
rect 22194 6076 22204 6132
rect 22260 6076 23660 6132
rect 23716 6076 24332 6132
rect 24388 6076 24398 6132
rect 24742 6076 24780 6132
rect 24836 6076 24846 6132
rect 25452 6076 28476 6132
rect 28532 6076 28542 6132
rect 39778 6076 39788 6132
rect 39844 6076 43708 6132
rect 43764 6076 43774 6132
rect 44146 6076 44156 6132
rect 44212 6076 46396 6132
rect 46452 6076 47068 6132
rect 47124 6076 48188 6132
rect 48244 6076 48254 6132
rect 49420 6076 50316 6132
rect 50372 6076 52108 6132
rect 52164 6076 52174 6132
rect 13906 5964 13916 6020
rect 13972 5964 25228 6020
rect 25284 5964 25294 6020
rect 16706 5852 16716 5908
rect 16772 5852 19068 5908
rect 19124 5852 19852 5908
rect 19908 5852 19918 5908
rect 20850 5852 20860 5908
rect 20916 5852 22428 5908
rect 22484 5852 22494 5908
rect 23538 5852 23548 5908
rect 23604 5852 23660 5908
rect 23716 5852 23726 5908
rect 25452 5796 25508 6076
rect 26786 5964 26796 6020
rect 26852 5964 28140 6020
rect 28196 5964 28206 6020
rect 30146 5964 30156 6020
rect 30212 5964 31052 6020
rect 31108 5964 31118 6020
rect 31602 5964 31612 6020
rect 31668 5964 32620 6020
rect 32676 5964 34076 6020
rect 34132 5964 34142 6020
rect 35186 5964 35196 6020
rect 35252 5964 37324 6020
rect 37380 5964 38108 6020
rect 38164 5964 38174 6020
rect 45042 5964 45052 6020
rect 45108 5964 45612 6020
rect 45668 5964 46228 6020
rect 48066 5964 48076 6020
rect 48132 5964 48748 6020
rect 48804 5964 48814 6020
rect 46172 5908 46228 5964
rect 31714 5852 31724 5908
rect 31780 5852 32396 5908
rect 32452 5852 33292 5908
rect 33348 5852 33358 5908
rect 33506 5852 33516 5908
rect 33572 5852 34300 5908
rect 34356 5852 34366 5908
rect 36306 5852 36316 5908
rect 36372 5852 38444 5908
rect 38500 5852 38510 5908
rect 40002 5852 40012 5908
rect 40068 5852 41916 5908
rect 41972 5852 44828 5908
rect 44884 5852 45836 5908
rect 45892 5852 45902 5908
rect 46162 5852 46172 5908
rect 46228 5852 46238 5908
rect 16370 5740 16380 5796
rect 16436 5740 25508 5796
rect 29138 5740 29148 5796
rect 29204 5740 33068 5796
rect 33124 5740 33628 5796
rect 33684 5740 33694 5796
rect 23314 5628 23324 5684
rect 23380 5628 25900 5684
rect 25956 5628 25966 5684
rect 28354 5628 28364 5684
rect 28420 5628 29596 5684
rect 29652 5628 29662 5684
rect 32498 5628 32508 5684
rect 32564 5628 32844 5684
rect 32900 5628 32910 5684
rect 44146 5628 44156 5684
rect 44212 5628 44940 5684
rect 44996 5628 45724 5684
rect 45780 5628 45790 5684
rect 23762 5516 23772 5572
rect 23828 5516 24108 5572
rect 24164 5516 24174 5572
rect 30370 5516 30380 5572
rect 30436 5516 31500 5572
rect 31556 5516 31566 5572
rect 38322 5516 38332 5572
rect 38388 5516 40236 5572
rect 40292 5516 40302 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 32050 5404 32060 5460
rect 32116 5404 33460 5460
rect 33404 5348 33460 5404
rect 20290 5292 20300 5348
rect 20356 5292 21084 5348
rect 21140 5292 21150 5348
rect 25890 5292 25900 5348
rect 25956 5292 32788 5348
rect 33394 5292 33404 5348
rect 33460 5292 33964 5348
rect 34020 5292 34030 5348
rect 35970 5292 35980 5348
rect 36036 5292 38780 5348
rect 38836 5292 38846 5348
rect 39778 5292 39788 5348
rect 39844 5292 47292 5348
rect 47348 5292 47358 5348
rect 32732 5236 32788 5292
rect 19954 5180 19964 5236
rect 20020 5180 21644 5236
rect 21700 5180 21710 5236
rect 22978 5180 22988 5236
rect 23044 5180 23884 5236
rect 23940 5180 24668 5236
rect 24724 5180 24734 5236
rect 26674 5180 26684 5236
rect 26740 5180 27020 5236
rect 27076 5180 27086 5236
rect 32732 5180 42252 5236
rect 42308 5180 43036 5236
rect 43092 5180 50764 5236
rect 50820 5180 50830 5236
rect 15474 5068 15484 5124
rect 15540 5068 16940 5124
rect 16996 5068 17006 5124
rect 26002 5068 26012 5124
rect 26068 5068 28028 5124
rect 28084 5068 30156 5124
rect 30212 5068 30222 5124
rect 30706 5068 30716 5124
rect 30772 5068 32060 5124
rect 32116 5068 32126 5124
rect 34290 5068 34300 5124
rect 34356 5068 34972 5124
rect 35028 5068 35038 5124
rect 38322 5068 38332 5124
rect 38388 5068 40124 5124
rect 40180 5068 40190 5124
rect 46834 5068 46844 5124
rect 46900 5068 50204 5124
rect 50260 5068 51100 5124
rect 51156 5068 51166 5124
rect 23202 4956 23212 5012
rect 23268 4956 24108 5012
rect 24164 4956 24174 5012
rect 30818 4956 30828 5012
rect 30884 4956 32172 5012
rect 32228 4956 32238 5012
rect 33506 4956 33516 5012
rect 33572 4956 34860 5012
rect 34916 4956 34926 5012
rect 42018 4956 42028 5012
rect 42084 4956 43372 5012
rect 43428 4956 44940 5012
rect 44996 4956 45006 5012
rect 48486 4956 48524 5012
rect 48580 4956 48590 5012
rect 21970 4844 21980 4900
rect 22036 4844 26124 4900
rect 26180 4844 26460 4900
rect 26516 4844 26684 4900
rect 26740 4844 26750 4900
rect 35970 4844 35980 4900
rect 36036 4844 36988 4900
rect 37044 4844 37054 4900
rect 38434 4844 38444 4900
rect 38500 4844 38668 4900
rect 38724 4844 38734 4900
rect 22754 4732 22764 4788
rect 22820 4732 23660 4788
rect 23716 4732 23726 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 24220 4620 27468 4676
rect 27524 4620 27534 4676
rect 34962 4620 34972 4676
rect 35028 4620 47964 4676
rect 48020 4620 48030 4676
rect 24220 4564 24276 4620
rect 24210 4508 24220 4564
rect 24276 4508 24286 4564
rect 24658 4508 24668 4564
rect 24724 4508 25452 4564
rect 25508 4508 25518 4564
rect 26898 4508 26908 4564
rect 26964 4508 27916 4564
rect 27972 4508 29260 4564
rect 29316 4508 29326 4564
rect 36082 4508 36092 4564
rect 36148 4508 36876 4564
rect 36932 4508 36942 4564
rect 44594 4508 44604 4564
rect 44660 4508 45724 4564
rect 45780 4508 46956 4564
rect 47012 4508 47022 4564
rect 50372 4508 56364 4564
rect 56420 4508 56430 4564
rect 25452 4452 25508 4508
rect 25452 4396 37436 4452
rect 37492 4396 37502 4452
rect 40226 4396 40236 4452
rect 40292 4396 48076 4452
rect 48132 4396 48142 4452
rect 16930 4284 16940 4340
rect 16996 4284 27916 4340
rect 27972 4284 29596 4340
rect 29652 4284 31948 4340
rect 32004 4284 32014 4340
rect 33394 4284 33404 4340
rect 33460 4284 37548 4340
rect 37604 4284 37614 4340
rect 41346 4284 41356 4340
rect 41412 4284 42700 4340
rect 42756 4284 42766 4340
rect 43138 4284 43148 4340
rect 43204 4284 46732 4340
rect 46788 4284 46798 4340
rect 50372 4228 50428 4508
rect 49298 4172 49308 4228
rect 49364 4172 50428 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 27458 3836 27468 3892
rect 27524 3836 31052 3892
rect 31108 3836 31118 3892
rect 27010 3724 27020 3780
rect 27076 3724 32956 3780
rect 33012 3724 33964 3780
rect 34020 3724 34030 3780
rect 39890 3724 39900 3780
rect 39956 3724 46564 3780
rect 46508 3668 46564 3724
rect 26114 3612 26124 3668
rect 26180 3612 31500 3668
rect 31556 3612 31566 3668
rect 42690 3612 42700 3668
rect 42756 3612 44268 3668
rect 44324 3612 44334 3668
rect 46498 3612 46508 3668
rect 46564 3612 48524 3668
rect 48580 3612 48590 3668
rect 25666 3500 25676 3556
rect 25732 3500 29484 3556
rect 29540 3500 30044 3556
rect 30100 3500 30110 3556
rect 30258 3500 30268 3556
rect 30324 3500 38332 3556
rect 38388 3500 38398 3556
rect 38658 3500 38668 3556
rect 38724 3500 46844 3556
rect 46900 3500 47516 3556
rect 47572 3500 49308 3556
rect 49364 3500 49374 3556
rect 26562 3388 26572 3444
rect 26628 3388 32284 3444
rect 32340 3388 32350 3444
rect 35522 3276 35532 3332
rect 35588 3276 36316 3332
rect 36372 3276 51772 3332
rect 51828 3276 51838 3332
rect 23202 3164 23212 3220
rect 23268 3164 46396 3220
rect 46452 3164 46462 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 13794 2940 13804 2996
rect 13860 2940 39676 2996
rect 39732 2940 39742 2996
<< via3 >>
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 51660 58492 51716 58548
rect 50316 58380 50372 58436
rect 48076 58156 48132 58212
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 52892 56588 52948 56644
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 23772 55356 23828 55412
rect 25452 55020 25508 55076
rect 43932 55020 43988 55076
rect 47180 55020 47236 55076
rect 51212 55020 51268 55076
rect 45052 54908 45108 54964
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 18060 54796 18116 54852
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 34524 54684 34580 54740
rect 11340 54236 11396 54292
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 13580 54012 13636 54068
rect 18060 54012 18116 54068
rect 16044 53676 16100 53732
rect 22876 53564 22932 53620
rect 45052 53564 45108 53620
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 13580 53228 13636 53284
rect 34524 53228 34580 53284
rect 49196 53228 49252 53284
rect 14476 53116 14532 53172
rect 34188 52892 34244 52948
rect 49980 52892 50036 52948
rect 16044 52668 16100 52724
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 14476 52444 14532 52500
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 43820 52444 43876 52500
rect 8428 52220 8484 52276
rect 50316 51996 50372 52052
rect 14476 51884 14532 51940
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 25452 51660 25508 51716
rect 15372 51548 15428 51604
rect 6860 51212 6916 51268
rect 50316 51324 50372 51380
rect 49868 51212 49924 51268
rect 43820 51100 43876 51156
rect 48748 50988 48804 51044
rect 51772 50988 51828 51044
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 43932 50876 43988 50932
rect 51660 50764 51716 50820
rect 50316 50652 50372 50708
rect 34524 50540 34580 50596
rect 42812 50540 42868 50596
rect 4284 50428 4340 50484
rect 51884 50428 51940 50484
rect 61516 50316 61572 50372
rect 49980 50204 50036 50260
rect 51772 50204 51828 50260
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 50204 50092 50260 50148
rect 55804 50092 55860 50148
rect 14140 49644 14196 49700
rect 61516 49644 61572 49700
rect 34188 49420 34244 49476
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 8428 49196 8484 49252
rect 14140 49196 14196 49252
rect 11340 48860 11396 48916
rect 60732 48860 60788 48916
rect 1708 48748 1764 48804
rect 3948 48748 4004 48804
rect 42812 48636 42868 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 49196 48524 49252 48580
rect 45276 48412 45332 48468
rect 57036 48412 57092 48468
rect 50316 48300 50372 48356
rect 51884 48300 51940 48356
rect 62076 48300 62132 48356
rect 57932 48188 57988 48244
rect 1708 48076 1764 48132
rect 51660 47964 51716 48020
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 13020 47516 13076 47572
rect 54236 47516 54292 47572
rect 60620 47404 60676 47460
rect 48748 47068 48804 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 24668 46956 24724 47012
rect 60732 46956 60788 47012
rect 61292 46956 61348 47012
rect 61964 46956 62020 47012
rect 22988 46844 23044 46900
rect 62188 46844 62244 46900
rect 10892 46732 10948 46788
rect 61740 46732 61796 46788
rect 4060 46620 4116 46676
rect 48076 46620 48132 46676
rect 48748 46620 48804 46676
rect 61404 46620 61460 46676
rect 50988 46396 51044 46452
rect 19404 46284 19460 46340
rect 61740 46284 61796 46340
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 27916 46172 27972 46228
rect 53340 46172 53396 46228
rect 62076 46172 62132 46228
rect 33516 46060 33572 46116
rect 42140 45948 42196 46004
rect 20412 45836 20468 45892
rect 33628 45836 33684 45892
rect 53452 45836 53508 45892
rect 61292 45836 61348 45892
rect 62188 45836 62244 45892
rect 50988 45724 51044 45780
rect 20860 45612 20916 45668
rect 50204 45500 50260 45556
rect 53340 45500 53396 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 43932 45388 43988 45444
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 8428 45276 8484 45332
rect 25452 45276 25508 45332
rect 25676 45276 25732 45332
rect 3388 45164 3444 45220
rect 48748 45164 48804 45220
rect 61404 45052 61460 45108
rect 55580 44940 55636 44996
rect 16492 44828 16548 44884
rect 57932 44828 57988 44884
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 25452 44604 25508 44660
rect 43708 44492 43764 44548
rect 10892 44268 10948 44324
rect 54012 44380 54068 44436
rect 28700 44044 28756 44100
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 3836 43820 3892 43876
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 48748 43820 48804 43876
rect 56700 43820 56756 43876
rect 22988 43596 23044 43652
rect 60620 43708 60676 43764
rect 61964 43484 62020 43540
rect 4172 43372 4228 43428
rect 27916 43372 27972 43428
rect 24668 43260 24724 43316
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 13020 43036 13076 43092
rect 15148 42924 15204 42980
rect 19516 42924 19572 42980
rect 14588 42700 14644 42756
rect 17612 42700 17668 42756
rect 21532 42700 21588 42756
rect 4284 42476 4340 42532
rect 3388 42364 3444 42420
rect 61964 42364 62020 42420
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4172 42252 4228 42308
rect 27804 42252 27860 42308
rect 6860 42140 6916 42196
rect 32172 42140 32228 42196
rect 43708 42140 43764 42196
rect 53452 42140 53508 42196
rect 14588 42028 14644 42084
rect 15148 42028 15204 42084
rect 3836 41916 3892 41972
rect 56700 41916 56756 41972
rect 57036 41916 57092 41972
rect 61852 41804 61908 41860
rect 45276 41692 45332 41748
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 32172 41468 32228 41524
rect 51212 41468 51268 41524
rect 44156 41356 44212 41412
rect 55804 41356 55860 41412
rect 25676 41020 25732 41076
rect 52892 41132 52948 41188
rect 34524 40908 34580 40964
rect 61964 40908 62020 40964
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 43932 40572 43988 40628
rect 27580 40460 27636 40516
rect 45276 40460 45332 40516
rect 14588 40348 14644 40404
rect 47180 40460 47236 40516
rect 54236 40460 54292 40516
rect 61516 40348 61572 40404
rect 48636 40236 48692 40292
rect 61964 40124 62020 40180
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 16492 39900 16548 39956
rect 62076 39900 62132 39956
rect 54012 39788 54068 39844
rect 51212 39452 51268 39508
rect 61292 39340 61348 39396
rect 17612 39228 17668 39284
rect 19404 39228 19460 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 49196 39116 49252 39172
rect 3948 39004 4004 39060
rect 41692 39004 41748 39060
rect 42140 39004 42196 39060
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 46732 38892 46788 38948
rect 33404 38780 33460 38836
rect 49868 38780 49924 38836
rect 20860 38556 20916 38612
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19516 38332 19572 38388
rect 46732 38332 46788 38388
rect 48076 38220 48132 38276
rect 21532 37996 21588 38052
rect 33516 37884 33572 37940
rect 20412 37772 20468 37828
rect 28700 37772 28756 37828
rect 50204 37772 50260 37828
rect 3948 37660 4004 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 34524 37660 34580 37716
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 33628 37436 33684 37492
rect 49196 37436 49252 37492
rect 4060 37324 4116 37380
rect 33404 37212 33460 37268
rect 62076 37212 62132 37268
rect 25676 36876 25732 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 61292 36428 61348 36484
rect 48076 36092 48132 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 15148 35980 15204 36036
rect 45164 35868 45220 35924
rect 57596 35756 57652 35812
rect 55580 35532 55636 35588
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 9884 35196 9940 35252
rect 45164 35196 45220 35252
rect 56028 35084 56084 35140
rect 27580 34748 27636 34804
rect 9436 34636 9492 34692
rect 27132 34636 27188 34692
rect 29372 34636 29428 34692
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 15372 34412 15428 34468
rect 29372 34188 29428 34244
rect 7756 34076 7812 34132
rect 50204 34076 50260 34132
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 32508 33628 32564 33684
rect 56140 33628 56196 33684
rect 11340 33516 11396 33572
rect 13356 33516 13412 33572
rect 48636 33516 48692 33572
rect 29372 33404 29428 33460
rect 41692 33404 41748 33460
rect 61404 33292 61460 33348
rect 14252 33068 14308 33124
rect 61628 32956 61684 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 5292 32732 5348 32788
rect 13356 32620 13412 32676
rect 32508 32396 32564 32452
rect 36204 32284 36260 32340
rect 17724 32172 17780 32228
rect 56252 32172 56308 32228
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 23772 32060 23828 32116
rect 34412 31948 34468 32004
rect 14364 31724 14420 31780
rect 6860 31612 6916 31668
rect 7756 31612 7812 31668
rect 34188 31612 34244 31668
rect 9436 31500 9492 31556
rect 15148 31500 15204 31556
rect 31276 31500 31332 31556
rect 50988 31500 51044 31556
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 12012 31276 12068 31332
rect 51100 31164 51156 31220
rect 15148 31052 15204 31108
rect 34412 30828 34468 30884
rect 51436 30716 51492 30772
rect 34188 30604 34244 30660
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 7756 30380 7812 30436
rect 51436 30380 51492 30436
rect 61628 30044 61684 30100
rect 55804 29932 55860 29988
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 3724 29708 3780 29764
rect 9884 29596 9940 29652
rect 38668 29596 38724 29652
rect 44268 29484 44324 29540
rect 57596 29372 57652 29428
rect 35756 29260 35812 29316
rect 40236 29260 40292 29316
rect 43372 29260 43428 29316
rect 35868 29148 35924 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 56364 28924 56420 28980
rect 12684 28812 12740 28868
rect 45164 28812 45220 28868
rect 56252 28700 56308 28756
rect 38556 28588 38612 28644
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 36204 28364 36260 28420
rect 35868 28252 35924 28308
rect 37660 28252 37716 28308
rect 45164 28252 45220 28308
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 40236 28028 40292 28084
rect 56364 28028 56420 28084
rect 11340 27804 11396 27860
rect 35756 27804 35812 27860
rect 31500 27692 31556 27748
rect 46732 27804 46788 27860
rect 35868 27468 35924 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 51436 27580 51492 27636
rect 37660 27468 37716 27524
rect 26796 27356 26852 27412
rect 26796 27132 26852 27188
rect 7868 27020 7924 27076
rect 46172 27020 46228 27076
rect 7084 26908 7140 26964
rect 27132 26908 27188 26964
rect 55804 26908 55860 26964
rect 6748 26796 6804 26852
rect 43372 26796 43428 26852
rect 38556 26684 38612 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 30604 26572 30660 26628
rect 23324 26348 23380 26404
rect 12684 26236 12740 26292
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 56140 26348 56196 26404
rect 56028 26236 56084 26292
rect 22876 26012 22932 26068
rect 4284 25900 4340 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 50316 25788 50372 25844
rect 42812 25676 42868 25732
rect 4284 25564 4340 25620
rect 55692 25564 55748 25620
rect 18396 25452 18452 25508
rect 44268 25452 44324 25508
rect 18060 25340 18116 25396
rect 23212 25340 23268 25396
rect 12012 25228 12068 25284
rect 12460 25228 12516 25284
rect 22876 25228 22932 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 50204 25004 50260 25060
rect 30604 24892 30660 24948
rect 31388 24892 31444 24948
rect 50092 24780 50148 24836
rect 17276 24668 17332 24724
rect 18396 24668 18452 24724
rect 31500 24668 31556 24724
rect 24108 24444 24164 24500
rect 50988 24332 51044 24388
rect 61852 24332 61908 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 44156 24220 44212 24276
rect 45388 24220 45444 24276
rect 50316 24220 50372 24276
rect 12460 24108 12516 24164
rect 17724 24108 17780 24164
rect 23324 23996 23380 24052
rect 50092 23996 50148 24052
rect 6748 23884 6804 23940
rect 7084 23884 7140 23940
rect 33516 23884 33572 23940
rect 50204 23884 50260 23940
rect 23212 23772 23268 23828
rect 9436 23660 9492 23716
rect 3724 23548 3780 23604
rect 5516 23548 5572 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50092 23660 50148 23716
rect 51100 23660 51156 23716
rect 38668 23548 38724 23604
rect 45388 23548 45444 23604
rect 46172 23548 46228 23604
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 7868 23436 7924 23492
rect 24108 23324 24164 23380
rect 24780 23324 24836 23380
rect 60956 23212 61012 23268
rect 36428 23100 36484 23156
rect 6972 22988 7028 23044
rect 23548 22988 23604 23044
rect 27580 22988 27636 23044
rect 48188 22988 48244 23044
rect 16940 22876 16996 22932
rect 18060 22876 18116 22932
rect 46172 22876 46228 22932
rect 14924 22764 14980 22820
rect 34524 22764 34580 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 12012 22540 12068 22596
rect 14476 22540 14532 22596
rect 32732 22428 32788 22484
rect 33292 22428 33348 22484
rect 45500 22428 45556 22484
rect 12348 22204 12404 22260
rect 12908 22204 12964 22260
rect 49084 22204 49140 22260
rect 49644 22204 49700 22260
rect 6636 22092 6692 22148
rect 25004 22092 25060 22148
rect 36428 22092 36484 22148
rect 60956 22092 61012 22148
rect 43372 21980 43428 22036
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 49420 21868 49476 21924
rect 4284 21756 4340 21812
rect 16940 21644 16996 21700
rect 20972 21532 21028 21588
rect 34748 21532 34804 21588
rect 49532 21532 49588 21588
rect 15036 21420 15092 21476
rect 17276 21420 17332 21476
rect 60844 21308 60900 21364
rect 33516 21196 33572 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 6524 20972 6580 21028
rect 33404 20972 33460 21028
rect 51212 20860 51268 20916
rect 49084 20524 49140 20580
rect 14924 20300 14980 20356
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 30940 20412 30996 20468
rect 61180 20412 61236 20468
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 5292 19964 5348 20020
rect 24892 19964 24948 20020
rect 33292 19852 33348 19908
rect 34524 19852 34580 19908
rect 12348 19740 12404 19796
rect 43596 19740 43652 19796
rect 6524 19628 6580 19684
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 49420 19404 49476 19460
rect 12348 19180 12404 19236
rect 25004 18956 25060 19012
rect 49420 18844 49476 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 3612 18732 3668 18788
rect 5292 18620 5348 18676
rect 49644 18620 49700 18676
rect 60956 18620 61012 18676
rect 5516 18396 5572 18452
rect 6972 18396 7028 18452
rect 39788 18396 39844 18452
rect 21756 18284 21812 18340
rect 50092 18284 50148 18340
rect 61852 18284 61908 18340
rect 25004 18172 25060 18228
rect 11900 18060 11956 18116
rect 12908 18060 12964 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 6636 17948 6692 18004
rect 3724 17724 3780 17780
rect 49084 17612 49140 17668
rect 49532 17500 49588 17556
rect 50204 17500 50260 17556
rect 60844 17500 60900 17556
rect 14252 17388 14308 17444
rect 24780 17388 24836 17444
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 49196 17388 49252 17444
rect 24780 17052 24836 17108
rect 14476 16940 14532 16996
rect 4284 16828 4340 16884
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 50204 16940 50260 16996
rect 47740 16716 47796 16772
rect 12012 16604 12068 16660
rect 23548 16492 23604 16548
rect 27468 16492 27524 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 13804 16380 13860 16436
rect 43596 16380 43652 16436
rect 61180 16380 61236 16436
rect 49084 16268 49140 16324
rect 48972 16156 49028 16212
rect 27804 16044 27860 16100
rect 3612 15932 3668 15988
rect 27468 15820 27524 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 23996 15596 24052 15652
rect 36428 15596 36484 15652
rect 44268 15596 44324 15652
rect 61404 15484 61460 15540
rect 49532 15372 49588 15428
rect 3724 15036 3780 15092
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 25004 15148 25060 15204
rect 40908 15148 40964 15204
rect 49308 15036 49364 15092
rect 13804 14924 13860 14980
rect 23436 14812 23492 14868
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 49308 14812 49364 14868
rect 49532 14812 49588 14868
rect 33404 14700 33460 14756
rect 6300 14588 6356 14644
rect 14812 14588 14868 14644
rect 61628 14588 61684 14644
rect 49196 14364 49252 14420
rect 34748 14140 34804 14196
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 32732 13916 32788 13972
rect 39564 13916 39620 13972
rect 54012 13916 54068 13972
rect 30940 13692 30996 13748
rect 48972 13580 49028 13636
rect 39564 13468 39620 13524
rect 50204 13468 50260 13524
rect 54012 13468 54068 13524
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 6300 13356 6356 13412
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 48524 13244 48580 13300
rect 48188 13020 48244 13076
rect 50092 12908 50148 12964
rect 40796 12796 40852 12852
rect 44268 12796 44324 12852
rect 22652 12684 22708 12740
rect 48524 12684 48580 12740
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 55692 12572 55748 12628
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 27468 12460 27524 12516
rect 43372 12236 43428 12292
rect 51212 12236 51268 12292
rect 11900 12124 11956 12180
rect 23996 12012 24052 12068
rect 47740 12012 47796 12068
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 22652 11676 22708 11732
rect 12572 11452 12628 11508
rect 46844 11452 46900 11508
rect 18620 11004 18676 11060
rect 20860 11004 20916 11060
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 27804 10892 27860 10948
rect 31276 10332 31332 10388
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 18620 10108 18676 10164
rect 31388 9884 31444 9940
rect 39900 9884 39956 9940
rect 39788 9548 39844 9604
rect 42812 9436 42868 9492
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 43596 9212 43652 9268
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 27692 8876 27748 8932
rect 31948 8764 32004 8820
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 39900 8540 39956 8596
rect 12572 8316 12628 8372
rect 14812 7980 14868 8036
rect 27804 7980 27860 8036
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 23548 6636 23604 6692
rect 24892 6636 24948 6692
rect 27692 6636 27748 6692
rect 20860 6300 20916 6356
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 23436 6188 23492 6244
rect 20972 6076 21028 6132
rect 21756 6076 21812 6132
rect 24780 6076 24836 6132
rect 23548 5852 23604 5908
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 39788 5292 39844 5348
rect 48524 4956 48580 5012
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 31948 4284 32004 4340
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 39676 2940 39732 2996
<< metal4 >>
rect 4448 60396 4768 60428
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 19808 59612 20128 60428
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 35168 60396 35488 60428
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 50528 59612 50848 60428
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50316 58436 50372 58446
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 18060 54852 18116 54862
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 11340 54292 11396 54302
rect 8428 52276 8484 52286
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4284 50484 4340 50494
rect 1708 48804 1764 48814
rect 1708 48132 1764 48748
rect 1708 48066 1764 48076
rect 3948 48804 4004 48814
rect 3388 45220 3444 45230
rect 3388 42420 3444 45164
rect 3388 42354 3444 42364
rect 3836 43876 3892 43886
rect 3836 41972 3892 43820
rect 3836 41906 3892 41916
rect 3948 39060 4004 48748
rect 3948 37716 4004 39004
rect 3948 37650 4004 37660
rect 4060 46676 4116 46686
rect 4060 37380 4116 46620
rect 4172 43428 4228 43438
rect 4172 42308 4228 43372
rect 4172 42242 4228 42252
rect 4284 42532 4340 50428
rect 4060 37314 4116 37324
rect 3724 29764 3780 29774
rect 3724 23604 3780 29708
rect 4284 25956 4340 42476
rect 4284 25620 4340 25900
rect 4284 25554 4340 25564
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 6860 51268 6916 51278
rect 6860 42196 6916 51212
rect 8428 49252 8484 52220
rect 8428 45332 8484 49196
rect 11340 48916 11396 54236
rect 13580 54068 13636 54078
rect 13580 53284 13636 54012
rect 18060 54068 18116 54796
rect 18060 54002 18116 54012
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 13580 53218 13636 53228
rect 16044 53732 16100 53742
rect 14476 53172 14532 53182
rect 14476 52500 14532 53116
rect 16044 52724 16100 53676
rect 16044 52658 16100 52668
rect 19808 53340 20128 54852
rect 23772 55412 23828 55422
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 14476 52434 14532 52444
rect 14476 51940 14532 51950
rect 14476 50428 14532 51884
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 14364 50372 14532 50428
rect 15372 51604 15428 51614
rect 14140 49700 14196 49710
rect 14140 49252 14196 49644
rect 14140 49186 14196 49196
rect 11340 48850 11396 48860
rect 13020 47572 13076 47582
rect 8428 45266 8484 45276
rect 10892 46788 10948 46798
rect 10892 44324 10948 46732
rect 10892 44258 10948 44268
rect 13020 43092 13076 47516
rect 13020 43026 13076 43036
rect 6860 38668 6916 42140
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 3724 23538 3780 23548
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4284 21812 4340 21822
rect 3612 18788 3668 18798
rect 3612 15988 3668 18732
rect 3612 15922 3668 15932
rect 3724 17780 3780 17790
rect 3724 15092 3780 17724
rect 4284 16884 4340 21756
rect 4284 16818 4340 16828
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 5292 38612 6916 38668
rect 5292 32788 5348 38612
rect 9884 35252 9940 35262
rect 9436 34692 9492 34702
rect 5292 20020 5348 32732
rect 7756 34132 7812 34142
rect 6860 31668 6916 31678
rect 6860 26908 6916 31612
rect 7756 31668 7812 34076
rect 7756 30436 7812 31612
rect 7756 30370 7812 30380
rect 9436 31556 9492 34636
rect 7868 27076 7924 27086
rect 7084 26964 7140 26974
rect 6748 26852 6804 26862
rect 6860 26852 7028 26908
rect 6748 23940 6804 26796
rect 6748 23874 6804 23884
rect 5292 18676 5348 19964
rect 5292 18610 5348 18620
rect 5516 23604 5572 23614
rect 5516 18452 5572 23548
rect 6972 23044 7028 26852
rect 7084 23940 7140 26908
rect 7084 23874 7140 23884
rect 7868 23492 7924 27020
rect 9436 23716 9492 31500
rect 9884 29652 9940 35196
rect 9884 29586 9940 29596
rect 11340 33572 11396 33582
rect 11340 27860 11396 33516
rect 13356 33572 13412 33582
rect 13356 32676 13412 33516
rect 13356 32610 13412 32620
rect 14252 33124 14308 33134
rect 11340 27794 11396 27804
rect 12012 31332 12068 31342
rect 12012 25284 12068 31276
rect 12684 28868 12740 28878
rect 12684 26292 12740 28812
rect 12684 26226 12740 26236
rect 12012 25218 12068 25228
rect 12460 25284 12516 25294
rect 12460 24164 12516 25228
rect 12460 24098 12516 24108
rect 9436 23650 9492 23660
rect 7868 23426 7924 23436
rect 6636 22148 6692 22158
rect 6524 21028 6580 21038
rect 6524 19684 6580 20972
rect 6524 19618 6580 19628
rect 5516 18386 5572 18396
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 3724 15026 3780 15036
rect 4448 16492 4768 18004
rect 6636 18004 6692 22092
rect 6972 18452 7028 22988
rect 6972 18386 7028 18396
rect 12012 22596 12068 22606
rect 6636 17938 6692 17948
rect 11900 18116 11956 18126
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 6300 14644 6356 14654
rect 6300 13412 6356 14588
rect 6300 13346 6356 13356
rect 4448 11788 4768 13300
rect 11900 12180 11956 18060
rect 12012 16660 12068 22540
rect 12348 22260 12404 22270
rect 12348 19796 12404 22204
rect 12348 19236 12404 19740
rect 12348 19170 12404 19180
rect 12908 22260 12964 22270
rect 12908 18116 12964 22204
rect 12908 18050 12964 18060
rect 14252 17444 14308 33068
rect 14364 31780 14420 50372
rect 15148 42980 15204 42990
rect 14588 42756 14644 42766
rect 14588 42084 14644 42700
rect 14588 40404 14644 42028
rect 14588 40338 14644 40348
rect 15148 42084 15204 42924
rect 15148 36036 15204 42028
rect 15148 35970 15204 35980
rect 15372 34468 15428 51548
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19404 46340 19460 46350
rect 16492 44884 16548 44894
rect 16492 39956 16548 44828
rect 16492 39890 16548 39900
rect 17612 42756 17668 42766
rect 17612 39284 17668 42700
rect 17612 39218 17668 39228
rect 19404 39284 19460 46284
rect 19808 45500 20128 47012
rect 22876 53620 22932 53630
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19404 39218 19460 39228
rect 19516 42980 19572 42990
rect 19516 38388 19572 42924
rect 19516 38322 19572 38332
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 15372 34402 15428 34412
rect 19808 37660 20128 39172
rect 20412 45892 20468 45902
rect 20412 37828 20468 45836
rect 20860 45668 20916 45678
rect 20860 38612 20916 45612
rect 20860 38546 20916 38556
rect 21532 42756 21588 42766
rect 21532 38052 21588 42700
rect 21532 37986 21588 37996
rect 20412 37762 20468 37772
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 14364 31714 14420 31724
rect 17724 32228 17780 32238
rect 15148 31556 15204 31566
rect 15148 31108 15204 31500
rect 15148 31042 15204 31052
rect 17276 24724 17332 24734
rect 16940 22932 16996 22942
rect 14924 22820 14980 22830
rect 14252 17378 14308 17388
rect 14476 22596 14532 22606
rect 14476 16996 14532 22540
rect 14924 20356 14980 22764
rect 16940 21700 16996 22876
rect 16940 21634 16996 21644
rect 14924 20290 14980 20300
rect 15036 21476 15092 21486
rect 14476 16930 14532 16940
rect 12012 16594 12068 16604
rect 13804 16436 13860 16446
rect 13804 14980 13860 16380
rect 15036 15148 15092 21420
rect 17276 21476 17332 24668
rect 17724 24164 17780 32172
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 18396 25508 18452 25518
rect 17724 24098 17780 24108
rect 18060 25396 18116 25406
rect 18060 22932 18116 25340
rect 18396 24724 18452 25452
rect 18396 24658 18452 24668
rect 19808 25116 20128 26628
rect 22876 26068 22932 53564
rect 22988 46900 23044 46910
rect 22988 43652 23044 46844
rect 22988 43586 23044 43596
rect 23772 32116 23828 55356
rect 25452 55076 25508 55086
rect 25452 51716 25508 55020
rect 34524 54740 34580 54750
rect 34524 53284 34580 54684
rect 25452 51650 25508 51660
rect 34188 52948 34244 52958
rect 34188 49476 34244 52892
rect 34524 50596 34580 53228
rect 34524 50530 34580 50540
rect 35168 54124 35488 55636
rect 48076 58212 48132 58222
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 43932 55076 43988 55086
rect 35168 50988 35488 52500
rect 43820 52500 43876 52510
rect 43820 51156 43876 52444
rect 43820 51090 43876 51100
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 34188 49410 34244 49420
rect 35168 49420 35488 50932
rect 43932 50932 43988 55020
rect 47180 55076 47236 55086
rect 43932 50866 43988 50876
rect 45052 54964 45108 54974
rect 45052 53620 45108 54908
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 42812 50596 42868 50606
rect 42812 48692 42868 50540
rect 45052 50428 45108 53564
rect 45052 50372 45332 50428
rect 42812 48626 42868 48636
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 24668 47012 24724 47022
rect 24668 43316 24724 46956
rect 35168 46284 35488 47796
rect 27916 46228 27972 46238
rect 25452 45332 25508 45342
rect 25452 44660 25508 45276
rect 25452 44594 25508 44604
rect 25676 45332 25732 45342
rect 24668 43250 24724 43260
rect 25676 41076 25732 45276
rect 27916 43428 27972 46172
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 33516 46116 33572 46126
rect 27916 43362 27972 43372
rect 28700 44100 28756 44110
rect 25676 36932 25732 41020
rect 27804 42308 27860 42318
rect 25676 36866 25732 36876
rect 27580 40516 27636 40526
rect 27580 34804 27636 40460
rect 23772 32050 23828 32060
rect 27132 34692 27188 34702
rect 26796 27412 26852 27422
rect 26796 27188 26852 27356
rect 26796 27122 26852 27132
rect 27132 26964 27188 34636
rect 27132 26898 27188 26908
rect 22876 25284 22932 26012
rect 23324 26404 23380 26414
rect 22876 25218 22932 25228
rect 23212 25396 23268 25406
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 18060 22866 18116 22876
rect 19808 23548 20128 25060
rect 23212 23828 23268 25340
rect 23324 24052 23380 26348
rect 23324 23986 23380 23996
rect 24108 24500 24164 24510
rect 23212 23762 23268 23772
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 17276 21410 17332 21420
rect 19808 21980 20128 23492
rect 24108 23380 24164 24444
rect 24108 23314 24164 23324
rect 24780 23380 24836 23390
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 13804 14914 13860 14924
rect 14812 15092 15092 15148
rect 19808 20412 20128 21924
rect 23548 23044 23604 23054
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 11900 12114 11956 12124
rect 14812 14644 14868 15092
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 12572 11508 12628 11518
rect 12572 8372 12628 11452
rect 12572 8306 12628 8316
rect 14812 8036 14868 14588
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 18620 11060 18676 11070
rect 18620 10164 18676 11004
rect 18620 10098 18676 10108
rect 19808 11004 20128 12516
rect 20972 21588 21028 21598
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 14812 7970 14868 7980
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 20860 11060 20916 11070
rect 20860 6356 20916 11004
rect 20860 6290 20916 6300
rect 19808 4732 20128 6244
rect 20972 6132 21028 21532
rect 20972 6066 21028 6076
rect 21756 18340 21812 18350
rect 21756 6132 21812 18284
rect 23548 16548 23604 22988
rect 24780 17444 24836 23324
rect 27580 23044 27636 34748
rect 27580 22978 27636 22988
rect 25004 22148 25060 22158
rect 24780 17378 24836 17388
rect 24892 20020 24948 20030
rect 23548 16482 23604 16492
rect 24780 17108 24836 17118
rect 23996 15652 24052 15662
rect 23436 14868 23492 14878
rect 22652 12740 22708 12750
rect 22652 11732 22708 12684
rect 22652 11666 22708 11676
rect 23436 6244 23492 14812
rect 23996 12068 24052 15596
rect 23996 12002 24052 12012
rect 23436 6178 23492 6188
rect 23548 6692 23604 6702
rect 21756 6066 21812 6076
rect 23548 5908 23604 6636
rect 24780 6132 24836 17052
rect 24892 6692 24948 19964
rect 25004 19012 25060 22092
rect 25004 18228 25060 18956
rect 25004 15204 25060 18172
rect 25004 15138 25060 15148
rect 27468 16548 27524 16558
rect 27468 15876 27524 16492
rect 27804 16100 27860 42252
rect 28700 37828 28756 44044
rect 32172 42196 32228 42206
rect 32172 41524 32228 42140
rect 32172 41458 32228 41468
rect 28700 37762 28756 37772
rect 33404 38836 33460 38846
rect 33404 37268 33460 38780
rect 33516 37940 33572 46060
rect 33516 37874 33572 37884
rect 33628 45892 33684 45902
rect 33628 37492 33684 45836
rect 35168 44716 35488 46228
rect 45276 48468 45332 50372
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 34524 40964 34580 40974
rect 34524 37716 34580 40908
rect 34524 37650 34580 37660
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 42140 46004 42196 46014
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 33628 37426 33684 37436
rect 33404 37202 33460 37212
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 29372 34692 29428 34702
rect 29372 34244 29428 34636
rect 29372 33460 29428 34188
rect 35168 33740 35488 35252
rect 29372 33394 29428 33404
rect 32508 33684 32564 33694
rect 32508 32452 32564 33628
rect 32508 32386 32564 32396
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 41692 39060 41748 39070
rect 41692 33460 41748 39004
rect 42140 39060 42196 45948
rect 43932 45444 43988 45454
rect 43708 44548 43764 44558
rect 43708 42196 43764 44492
rect 43708 42130 43764 42140
rect 43932 40628 43988 45388
rect 45276 41748 45332 48412
rect 43932 40562 43988 40572
rect 44156 41412 44212 41422
rect 42140 38994 42196 39004
rect 41692 33394 41748 33404
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 34412 32004 34468 32014
rect 34188 31668 34244 31678
rect 31276 31556 31332 31566
rect 30604 26628 30660 26638
rect 30604 24948 30660 26572
rect 30604 24882 30660 24892
rect 27804 16034 27860 16044
rect 30940 20468 30996 20478
rect 27468 12516 27524 15820
rect 30940 13748 30996 20412
rect 30940 13682 30996 13692
rect 27468 12450 27524 12460
rect 27804 10948 27860 10958
rect 24892 6626 24948 6636
rect 27692 8932 27748 8942
rect 27692 6692 27748 8876
rect 27804 8036 27860 10892
rect 31276 10388 31332 31500
rect 34188 30660 34244 31612
rect 34412 30884 34468 31948
rect 34412 30818 34468 30828
rect 34188 30594 34244 30604
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 36204 32340 36260 32350
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 31500 27748 31556 27758
rect 31276 10322 31332 10332
rect 31388 24948 31444 24958
rect 31388 9940 31444 24892
rect 31500 24724 31556 27692
rect 31500 24658 31556 24668
rect 35168 27468 35488 28980
rect 35756 29316 35812 29326
rect 35756 27860 35812 29260
rect 35756 27794 35812 27804
rect 35868 29204 35924 29214
rect 35868 28308 35924 29148
rect 36204 28420 36260 32284
rect 38668 29652 38724 29662
rect 36204 28354 36260 28364
rect 38556 28644 38612 28654
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35868 27524 35924 28252
rect 35868 27458 35924 27468
rect 37660 28308 37716 28318
rect 37660 27524 37716 28252
rect 37660 27458 37716 27468
rect 35168 25900 35488 27412
rect 38556 26740 38612 28588
rect 38556 26674 38612 26684
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 33516 23940 33572 23950
rect 32732 22484 32788 22494
rect 32732 13972 32788 22428
rect 33292 22484 33348 22494
rect 33292 19908 33348 22428
rect 33516 21252 33572 23884
rect 33516 21186 33572 21196
rect 34524 22820 34580 22830
rect 33292 19842 33348 19852
rect 33404 21028 33460 21038
rect 33404 14756 33460 20972
rect 34524 19908 34580 22764
rect 35168 22764 35488 24276
rect 38668 23604 38724 29596
rect 40236 29316 40292 29326
rect 40236 28084 40292 29260
rect 40236 28018 40292 28028
rect 43372 29316 43428 29326
rect 43372 26852 43428 29260
rect 43372 26786 43428 26796
rect 38668 23538 38724 23548
rect 42812 25732 42868 25742
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 34524 19842 34580 19852
rect 34748 21588 34804 21598
rect 33404 14690 33460 14700
rect 34748 14196 34804 21532
rect 34748 14130 34804 14140
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 36428 23156 36484 23166
rect 36428 22148 36484 23100
rect 36428 15652 36484 22092
rect 36428 15586 36484 15596
rect 39788 18452 39844 18462
rect 39788 15148 39844 18396
rect 40908 15204 40964 15214
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 32732 13906 32788 13916
rect 31388 9874 31444 9884
rect 35168 13356 35488 14868
rect 39564 15092 39844 15148
rect 40796 15092 40964 15148
rect 39564 13972 39620 15092
rect 39564 13524 39620 13916
rect 39564 13458 39620 13468
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 40796 12852 40852 15092
rect 40796 12786 40852 12796
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 27804 7970 27860 7980
rect 31948 8820 32004 8830
rect 27692 6626 27748 6636
rect 24780 6066 24836 6076
rect 23548 5842 23604 5852
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 31948 4340 32004 8764
rect 31948 4274 32004 4284
rect 35168 8652 35488 10164
rect 39900 9940 39956 9950
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 39788 9604 39844 9614
rect 39788 5348 39844 9548
rect 39900 8596 39956 9884
rect 42812 9492 42868 25676
rect 44156 24276 44212 41356
rect 45276 40516 45332 41692
rect 45276 40450 45332 40460
rect 47180 40516 47236 55020
rect 48076 46676 48132 58156
rect 49196 53284 49252 53294
rect 48748 51044 48804 51054
rect 48748 47124 48804 50988
rect 49196 48580 49252 53228
rect 49980 52948 50036 52958
rect 49196 48514 49252 48524
rect 49868 51268 49924 51278
rect 48748 47058 48804 47068
rect 48076 46610 48132 46620
rect 48748 46676 48804 46686
rect 48748 45220 48804 46620
rect 48748 43876 48804 45164
rect 48748 43810 48804 43820
rect 47180 40450 47236 40460
rect 48636 40292 48692 40302
rect 46732 38948 46788 38958
rect 46732 38388 46788 38892
rect 46732 38322 46788 38332
rect 48076 38276 48132 38286
rect 48076 36148 48132 38220
rect 48076 36082 48132 36092
rect 45164 35924 45220 35934
rect 45164 35252 45220 35868
rect 45164 35186 45220 35196
rect 48636 33572 48692 40236
rect 49196 39172 49252 39182
rect 49196 37492 49252 39116
rect 49868 38836 49924 51212
rect 49980 50260 50036 52892
rect 50316 52052 50372 58380
rect 50316 51380 50372 51996
rect 50316 51314 50372 51324
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 51660 58548 51716 58558
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 49980 50194 50036 50204
rect 50316 50708 50372 50718
rect 50204 50148 50260 50158
rect 50204 45556 50260 50092
rect 50316 48356 50372 50652
rect 50316 48290 50372 48300
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50204 45490 50260 45500
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 51212 55076 51268 55086
rect 50988 46452 51044 46462
rect 50988 45780 51044 46396
rect 50988 45714 51044 45724
rect 49868 38770 49924 38780
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 51212 41524 51268 55020
rect 51660 50820 51716 58492
rect 52892 56644 52948 56654
rect 51660 48020 51716 50764
rect 51772 51044 51828 51054
rect 51772 50260 51828 50988
rect 51772 50194 51828 50204
rect 51884 50484 51940 50494
rect 51884 48356 51940 50428
rect 51884 48290 51940 48300
rect 51660 47954 51716 47964
rect 51212 39508 51268 41468
rect 52892 41188 52948 56588
rect 61516 50372 61572 50382
rect 55804 50148 55860 50158
rect 54236 47572 54292 47582
rect 53340 46228 53396 46238
rect 53340 45556 53396 46172
rect 53340 45490 53396 45500
rect 53452 45892 53508 45902
rect 53452 42196 53508 45836
rect 53452 42130 53508 42140
rect 54012 44436 54068 44446
rect 52892 41122 52948 41132
rect 54012 39844 54068 44380
rect 54236 40516 54292 47516
rect 54236 40450 54292 40460
rect 55580 44996 55636 45006
rect 54012 39778 54068 39788
rect 51212 39442 51268 39452
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 49196 37426 49252 37436
rect 50204 37828 50260 37838
rect 50204 34132 50260 37772
rect 50204 34066 50260 34076
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 55580 35588 55636 44940
rect 55804 41412 55860 50092
rect 61516 49700 61572 50316
rect 60732 48916 60788 48926
rect 57036 48468 57092 48478
rect 56700 43876 56756 43886
rect 56700 41972 56756 43820
rect 56700 41906 56756 41916
rect 57036 41972 57092 48412
rect 57932 48244 57988 48254
rect 57932 44884 57988 48188
rect 57932 44818 57988 44828
rect 60620 47460 60676 47470
rect 60620 43764 60676 47404
rect 60732 47012 60788 48860
rect 60732 46946 60788 46956
rect 61292 47012 61348 47022
rect 61292 45892 61348 46956
rect 61292 45826 61348 45836
rect 61404 46676 61460 46686
rect 61404 45108 61460 46620
rect 61404 45042 61460 45052
rect 60620 43698 60676 43708
rect 57036 41906 57092 41916
rect 55804 41346 55860 41356
rect 61516 40404 61572 49644
rect 62076 48356 62132 48366
rect 61964 47012 62020 47022
rect 61852 46956 61964 47012
rect 61740 46788 61796 46798
rect 61740 46340 61796 46732
rect 61740 46274 61796 46284
rect 61852 41860 61908 46956
rect 61964 46946 62020 46956
rect 62076 46228 62132 48300
rect 61964 43540 62020 43550
rect 61964 42420 62020 43484
rect 61964 42354 62020 42364
rect 61852 41794 61908 41804
rect 61516 40338 61572 40348
rect 61964 40964 62020 40974
rect 61964 40180 62020 40908
rect 61964 40114 62020 40124
rect 62076 39956 62132 46172
rect 62188 46900 62244 46910
rect 62188 45892 62244 46844
rect 62188 45826 62244 45836
rect 61292 39396 61348 39406
rect 61292 36484 61348 39340
rect 62076 37268 62132 39900
rect 62076 37202 62132 37212
rect 61292 36418 61348 36428
rect 55580 35522 55636 35532
rect 57596 35812 57652 35822
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 48636 33506 48692 33516
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 56028 35140 56084 35150
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 44268 29540 44324 29550
rect 44268 25508 44324 29484
rect 45164 28868 45220 28878
rect 45164 28308 45220 28812
rect 45164 28242 45220 28252
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 46732 27860 46788 27870
rect 44268 25442 44324 25452
rect 46172 27076 46228 27086
rect 44156 24210 44212 24220
rect 45388 24276 45444 24286
rect 45388 23604 45444 24220
rect 46172 23604 46228 27020
rect 46732 26908 46788 27804
rect 46732 26852 46900 26908
rect 45388 23492 45556 23548
rect 45500 22484 45556 23492
rect 46172 22932 46228 23548
rect 46172 22866 46228 22876
rect 45500 22418 45556 22428
rect 43372 22036 43428 22046
rect 43372 12292 43428 21980
rect 43372 12226 43428 12236
rect 43596 19796 43652 19806
rect 43596 16436 43652 19740
rect 42812 9426 42868 9436
rect 43596 9268 43652 16380
rect 44268 15652 44324 15662
rect 44268 12852 44324 15596
rect 44268 12786 44324 12796
rect 46844 11508 46900 26852
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50316 25844 50372 25854
rect 50204 25060 50260 25070
rect 50092 24836 50148 24846
rect 50092 24052 50148 24780
rect 50092 23716 50148 23996
rect 50204 23940 50260 25004
rect 50316 24276 50372 25788
rect 50316 24210 50372 24220
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50204 23874 50260 23884
rect 50092 23650 50148 23660
rect 50528 23548 50848 25060
rect 50988 31556 51044 31566
rect 50988 24388 51044 31500
rect 50988 24322 51044 24332
rect 51100 31220 51156 31230
rect 51100 23716 51156 31164
rect 51436 30772 51492 30782
rect 51436 30436 51492 30716
rect 51436 27636 51492 30380
rect 51436 27570 51492 27580
rect 55804 29988 55860 29998
rect 55804 26964 55860 29932
rect 55804 26898 55860 26908
rect 56028 26292 56084 35084
rect 56140 33684 56196 33694
rect 56140 26404 56196 33628
rect 56252 32228 56308 32238
rect 56252 28756 56308 32172
rect 57596 29428 57652 35756
rect 57596 29362 57652 29372
rect 61404 33348 61460 33358
rect 56252 28690 56308 28700
rect 56364 28980 56420 28990
rect 56364 28084 56420 28924
rect 56364 28018 56420 28028
rect 56140 26338 56196 26348
rect 56028 26226 56084 26236
rect 51100 23650 51156 23660
rect 55692 25620 55748 25630
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 48188 23044 48244 23054
rect 47740 16772 47796 16782
rect 47740 12068 47796 16716
rect 48188 13076 48244 22988
rect 49084 22260 49140 22270
rect 49084 20580 49140 22204
rect 49644 22260 49700 22270
rect 49084 20514 49140 20524
rect 49420 21924 49476 21934
rect 49420 19460 49476 21868
rect 49420 18900 49476 19404
rect 49420 18834 49476 18844
rect 49532 21588 49588 21598
rect 49084 17668 49140 17678
rect 49084 16324 49140 17612
rect 49532 17556 49588 21532
rect 49644 18676 49700 22204
rect 49644 18610 49700 18620
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 49532 17490 49588 17500
rect 50092 18340 50148 18350
rect 49084 16258 49140 16268
rect 49196 17444 49252 17454
rect 48972 16212 49028 16222
rect 48972 13636 49028 16156
rect 49196 14420 49252 17388
rect 49532 15428 49588 15438
rect 49308 15092 49364 15102
rect 49308 14868 49364 15036
rect 49308 14802 49364 14812
rect 49532 14868 49588 15372
rect 49532 14802 49588 14812
rect 49196 14354 49252 14364
rect 48972 13570 49028 13580
rect 48188 13010 48244 13020
rect 48524 13300 48580 13310
rect 47740 12002 47796 12012
rect 48524 12740 48580 13244
rect 50092 12964 50148 18284
rect 50204 17556 50260 17566
rect 50204 16996 50260 17500
rect 50204 13524 50260 16940
rect 50204 13458 50260 13468
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50092 12898 50148 12908
rect 46844 11442 46900 11452
rect 43596 9202 43652 9212
rect 39900 8530 39956 8540
rect 39788 3388 39844 5292
rect 48524 5012 48580 12684
rect 48524 4946 48580 4956
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 51212 20916 51268 20926
rect 51212 12292 51268 20860
rect 54012 13972 54068 13982
rect 54012 13524 54068 13916
rect 54012 13458 54068 13468
rect 55692 12628 55748 25564
rect 60956 23268 61012 23278
rect 60956 22148 61012 23212
rect 60844 21364 60900 21374
rect 60844 17556 60900 21308
rect 60956 18676 61012 22092
rect 60956 18610 61012 18620
rect 61180 20468 61236 20478
rect 60844 17490 60900 17500
rect 61180 16436 61236 20412
rect 61180 16370 61236 16380
rect 61404 15540 61460 33292
rect 61404 15474 61460 15484
rect 61628 33012 61684 33022
rect 61628 30100 61684 32956
rect 61628 14644 61684 30044
rect 61852 24388 61908 24398
rect 61852 18340 61908 24332
rect 61852 18274 61908 18284
rect 61628 14578 61684 14588
rect 55692 12562 55748 12572
rect 51212 12226 51268 12236
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 39676 3332 39844 3388
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 39676 2996 39732 3332
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 39676 2930 39732 2940
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1801_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1802_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35392 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1803_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37072 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1804_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 49504 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1805_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1806_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48384 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1807_
timestamp 1698431365
transform -1 0 50288 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1808_
timestamp 1698431365
transform 1 0 46592 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1809_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46592 0 -1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1810_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1811_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48720 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1812_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 49504 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1813_
timestamp 1698431365
transform 1 0 46704 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1814_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1815_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47488 0 1 29792
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1816_
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1817_
timestamp 1698431365
transform -1 0 51184 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1818_
timestamp 1698431365
transform -1 0 60032 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1819_
timestamp 1698431365
transform -1 0 61600 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1820_
timestamp 1698431365
transform 1 0 60368 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1821_
timestamp 1698431365
transform -1 0 60032 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1822_
timestamp 1698431365
transform -1 0 62160 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1823_
timestamp 1698431365
transform 1 0 54432 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1824_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1825_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1826_
timestamp 1698431365
transform -1 0 35728 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1827_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37184 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1828_
timestamp 1698431365
transform 1 0 37856 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1829_
timestamp 1698431365
transform 1 0 38752 0 1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1830_
timestamp 1698431365
transform 1 0 55328 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1831_
timestamp 1698431365
transform 1 0 50624 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1832_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 53424 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1833_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 49168 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1834_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 53536 0 -1 43904
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1835_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48608 0 1 51744
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1836_
timestamp 1698431365
transform -1 0 52864 0 -1 45472
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1837_
timestamp 1698431365
transform 1 0 53872 0 1 43904
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1838_
timestamp 1698431365
transform -1 0 52192 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1839_
timestamp 1698431365
transform -1 0 56224 0 1 42336
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1840_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48720 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1841_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 50624 0 -1 53312
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1842_
timestamp 1698431365
transform -1 0 18144 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1843_
timestamp 1698431365
transform -1 0 20944 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1844_
timestamp 1698431365
transform -1 0 22736 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1845_
timestamp 1698431365
transform -1 0 15680 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1846_
timestamp 1698431365
transform -1 0 15008 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1847_
timestamp 1698431365
transform -1 0 17472 0 1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1848_
timestamp 1698431365
transform -1 0 14224 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1849_
timestamp 1698431365
transform -1 0 16576 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1850_
timestamp 1698431365
transform -1 0 49504 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1851_
timestamp 1698431365
transform -1 0 50848 0 1 54880
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1852_
timestamp 1698431365
transform -1 0 23408 0 1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1853_
timestamp 1698431365
transform 1 0 32928 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1854_
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1855_
timestamp 1698431365
transform -1 0 32928 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1856_
timestamp 1698431365
transform 1 0 32032 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1857_
timestamp 1698431365
transform 1 0 3920 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1858_
timestamp 1698431365
transform -1 0 6384 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1859_
timestamp 1698431365
transform -1 0 4480 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1860_
timestamp 1698431365
transform 1 0 4368 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1861_
timestamp 1698431365
transform -1 0 7840 0 -1 48608
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1862_
timestamp 1698431365
transform 1 0 25424 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1863_
timestamp 1698431365
transform 1 0 26432 0 1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1864_
timestamp 1698431365
transform 1 0 24416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1865_
timestamp 1698431365
transform 1 0 19824 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1866_
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1867_
timestamp 1698431365
transform -1 0 14224 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1868_
timestamp 1698431365
transform 1 0 19824 0 -1 58016
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1869_
timestamp 1698431365
transform 1 0 22736 0 1 58016
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1870_
timestamp 1698431365
transform -1 0 30240 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1871_
timestamp 1698431365
transform -1 0 32928 0 1 58016
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1872_
timestamp 1698431365
transform 1 0 27216 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1873_
timestamp 1698431365
transform 1 0 25088 0 1 56448
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1874_
timestamp 1698431365
transform -1 0 29232 0 -1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1875_
timestamp 1698431365
transform 1 0 41104 0 1 56448
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1876_
timestamp 1698431365
transform -1 0 48384 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1877_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46032 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1878_
timestamp 1698431365
transform -1 0 51744 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1879_
timestamp 1698431365
transform -1 0 30128 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1880_
timestamp 1698431365
transform -1 0 28784 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1881_
timestamp 1698431365
transform -1 0 25872 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1882_
timestamp 1698431365
transform -1 0 33600 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1883_
timestamp 1698431365
transform -1 0 32704 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1884_
timestamp 1698431365
transform 1 0 34496 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1885_
timestamp 1698431365
transform 1 0 33600 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1886_
timestamp 1698431365
transform -1 0 36512 0 -1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1887_
timestamp 1698431365
transform 1 0 27216 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1888_
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1889_
timestamp 1698431365
transform 1 0 5824 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1890_
timestamp 1698431365
transform 1 0 1680 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1891_
timestamp 1698431365
transform -1 0 4032 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1892_
timestamp 1698431365
transform 1 0 4032 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1893_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3248 0 -1 37632
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1894_
timestamp 1698431365
transform -1 0 29120 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1895_
timestamp 1698431365
transform 1 0 30912 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1896_
timestamp 1698431365
transform -1 0 32256 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1897_
timestamp 1698431365
transform -1 0 28784 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1898_
timestamp 1698431365
transform -1 0 28224 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1899_
timestamp 1698431365
transform 1 0 29008 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1900_
timestamp 1698431365
transform 1 0 26656 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1901_
timestamp 1698431365
transform 1 0 27552 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1902_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28448 0 -1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1903_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1904_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 33712 0 1 37632
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1905_
timestamp 1698431365
transform 1 0 29792 0 1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1906_
timestamp 1698431365
transform -1 0 33712 0 1 36064
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1907_
timestamp 1698431365
transform -1 0 29344 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1908_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30464 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1909_
timestamp 1698431365
transform -1 0 53424 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1910_
timestamp 1698431365
transform 1 0 56224 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1911_
timestamp 1698431365
transform 1 0 61488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1912_
timestamp 1698431365
transform 1 0 60368 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1913_
timestamp 1698431365
transform 1 0 60368 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1914_
timestamp 1698431365
transform 1 0 59248 0 -1 45472
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1915_
timestamp 1698431365
transform -1 0 36400 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1916_
timestamp 1698431365
transform 1 0 36960 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1917_
timestamp 1698431365
transform -1 0 34944 0 -1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1918_
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1919_
timestamp 1698431365
transform 1 0 37072 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1920_
timestamp 1698431365
transform -1 0 38752 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1921_
timestamp 1698431365
transform 1 0 56448 0 -1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1922_
timestamp 1698431365
transform -1 0 50736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1923_
timestamp 1698431365
transform -1 0 46816 0 1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1924_
timestamp 1698431365
transform -1 0 48160 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1925_
timestamp 1698431365
transform 1 0 49728 0 -1 54880
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1926_
timestamp 1698431365
transform 1 0 58576 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1927_
timestamp 1698431365
transform 1 0 54544 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1928_
timestamp 1698431365
transform -1 0 54320 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1929_
timestamp 1698431365
transform -1 0 52304 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1930_
timestamp 1698431365
transform -1 0 54096 0 -1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1931_
timestamp 1698431365
transform -1 0 56112 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1932_
timestamp 1698431365
transform -1 0 55216 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1933_
timestamp 1698431365
transform 1 0 54096 0 -1 54880
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1934_
timestamp 1698431365
transform 1 0 58128 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1935_
timestamp 1698431365
transform 1 0 37632 0 1 54880
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1936_
timestamp 1698431365
transform -1 0 58352 0 1 54880
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1937_
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1938_
timestamp 1698431365
transform -1 0 56224 0 -1 51744
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1939_
timestamp 1698431365
transform 1 0 53536 0 1 53312
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1940_
timestamp 1698431365
transform 1 0 53424 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1941_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 52192 0 1 53312
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1942_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46144 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1943_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47264 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1944_
timestamp 1698431365
transform -1 0 35392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1945_
timestamp 1698431365
transform 1 0 34720 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1946_
timestamp 1698431365
transform -1 0 35616 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1947_
timestamp 1698431365
transform 1 0 37632 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1948_
timestamp 1698431365
transform 1 0 43568 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1949_
timestamp 1698431365
transform 1 0 44912 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1950_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1951_
timestamp 1698431365
transform 1 0 36960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1952_
timestamp 1698431365
transform 1 0 44464 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1953_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1954_
timestamp 1698431365
transform 1 0 48608 0 -1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1955_
timestamp 1698431365
transform 1 0 47712 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1956_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 53424 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1957_
timestamp 1698431365
transform -1 0 55776 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1958_
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1959_
timestamp 1698431365
transform 1 0 36400 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1960_
timestamp 1698431365
transform -1 0 42560 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1961_
timestamp 1698431365
transform -1 0 56224 0 -1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1962_
timestamp 1698431365
transform -1 0 59696 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1963_
timestamp 1698431365
transform -1 0 56112 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1964_
timestamp 1698431365
transform 1 0 61264 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1965_
timestamp 1698431365
transform 1 0 59472 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1966_
timestamp 1698431365
transform -1 0 58352 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1967_
timestamp 1698431365
transform -1 0 55216 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1968_
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1969_
timestamp 1698431365
transform 1 0 58128 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1970_
timestamp 1698431365
transform -1 0 56112 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1971_
timestamp 1698431365
transform 1 0 60368 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1972_
timestamp 1698431365
transform -1 0 56224 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1973_
timestamp 1698431365
transform 1 0 53536 0 -1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1974_
timestamp 1698431365
transform 1 0 61488 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1975_
timestamp 1698431365
transform -1 0 55440 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1976_
timestamp 1698431365
transform -1 0 57344 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1977_
timestamp 1698431365
transform -1 0 61040 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1978_
timestamp 1698431365
transform -1 0 58688 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1979_
timestamp 1698431365
transform -1 0 60144 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1980_
timestamp 1698431365
transform 1 0 60368 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1981_
timestamp 1698431365
transform 1 0 60368 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1982_
timestamp 1698431365
transform -1 0 62384 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1983_
timestamp 1698431365
transform 1 0 56672 0 1 42336
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1984_
timestamp 1698431365
transform -1 0 62384 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1985_
timestamp 1698431365
transform 1 0 58240 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1986_
timestamp 1698431365
transform -1 0 62384 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1987_
timestamp 1698431365
transform -1 0 57008 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1988_
timestamp 1698431365
transform -1 0 59248 0 1 39200
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1989_
timestamp 1698431365
transform -1 0 58240 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1990_
timestamp 1698431365
transform 1 0 54208 0 1 45472
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1991_
timestamp 1698431365
transform 1 0 54544 0 1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1992_
timestamp 1698431365
transform 1 0 57120 0 -1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1993_
timestamp 1698431365
transform -1 0 61264 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1994_
timestamp 1698431365
transform -1 0 60368 0 -1 40768
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1995_
timestamp 1698431365
transform 1 0 54768 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1996_
timestamp 1698431365
transform 1 0 54096 0 -1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1997_
timestamp 1698431365
transform -1 0 30128 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1998_
timestamp 1698431365
transform 1 0 29344 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1999_
timestamp 1698431365
transform -1 0 28784 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2000_
timestamp 1698431365
transform -1 0 23856 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2001_
timestamp 1698431365
transform 1 0 23520 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2002_
timestamp 1698431365
transform -1 0 27216 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2003_
timestamp 1698431365
transform 1 0 27888 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2004_
timestamp 1698431365
transform -1 0 29904 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2005_
timestamp 1698431365
transform -1 0 59472 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2006_
timestamp 1698431365
transform 1 0 53872 0 1 47040
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2007_
timestamp 1698431365
transform -1 0 31920 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2008_
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2009_
timestamp 1698431365
transform 1 0 38192 0 -1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2010_
timestamp 1698431365
transform -1 0 36512 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2011_
timestamp 1698431365
transform 1 0 33152 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2012_
timestamp 1698431365
transform -1 0 30016 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2013_
timestamp 1698431365
transform -1 0 32704 0 -1 58016
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2014_
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2015_
timestamp 1698431365
transform 1 0 31024 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2016_
timestamp 1698431365
transform 1 0 32256 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2017_
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2018_
timestamp 1698431365
transform 1 0 30128 0 1 50176
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2019_
timestamp 1698431365
transform 1 0 27552 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2020_
timestamp 1698431365
transform 1 0 29232 0 1 47040
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2021_
timestamp 1698431365
transform -1 0 33936 0 1 48608
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2022_
timestamp 1698431365
transform -1 0 36624 0 -1 51744
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2023_
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2024_
timestamp 1698431365
transform -1 0 34496 0 1 51744
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2025_
timestamp 1698431365
transform -1 0 32592 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2026_
timestamp 1698431365
transform 1 0 49056 0 -1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2027_
timestamp 1698431365
transform -1 0 53872 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2028_
timestamp 1698431365
transform 1 0 53424 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2029_
timestamp 1698431365
transform -1 0 53424 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2030_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 52528 0 -1 58016
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2031_
timestamp 1698431365
transform 1 0 51744 0 -1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2032_
timestamp 1698431365
transform -1 0 47936 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2033_
timestamp 1698431365
transform 1 0 44128 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2034_
timestamp 1698431365
transform -1 0 54768 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2035_
timestamp 1698431365
transform 1 0 57344 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2036_
timestamp 1698431365
transform 1 0 55328 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2037_
timestamp 1698431365
transform 1 0 54880 0 1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2038_
timestamp 1698431365
transform -1 0 40544 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2039_
timestamp 1698431365
transform -1 0 39984 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2040_
timestamp 1698431365
transform -1 0 39760 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2041_
timestamp 1698431365
transform -1 0 39312 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2042_
timestamp 1698431365
transform 1 0 39648 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2043_
timestamp 1698431365
transform -1 0 41440 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2044_
timestamp 1698431365
transform 1 0 43568 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2045_
timestamp 1698431365
transform 1 0 42112 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2046_
timestamp 1698431365
transform -1 0 57344 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2047_
timestamp 1698431365
transform 1 0 52752 0 1 50176
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2048_
timestamp 1698431365
transform 1 0 50176 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2049_
timestamp 1698431365
transform -1 0 45696 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2050_
timestamp 1698431365
transform -1 0 46368 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2051_
timestamp 1698431365
transform 1 0 45696 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2052_
timestamp 1698431365
transform 1 0 51072 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2053_
timestamp 1698431365
transform 1 0 46144 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2054_
timestamp 1698431365
transform 1 0 43568 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2055_
timestamp 1698431365
transform 1 0 45584 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2056_
timestamp 1698431365
transform -1 0 47600 0 1 48608
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2057_
timestamp 1698431365
transform -1 0 44016 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2058_
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2059_
timestamp 1698431365
transform -1 0 46928 0 -1 48608
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2060_
timestamp 1698431365
transform -1 0 48944 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2061_
timestamp 1698431365
transform -1 0 49504 0 1 45472
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2062_
timestamp 1698431365
transform -1 0 49168 0 1 47040
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2063_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 50064 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2064_
timestamp 1698431365
transform 1 0 48496 0 1 48608
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2065_
timestamp 1698431365
transform 1 0 50288 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2066_
timestamp 1698431365
transform 1 0 51632 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2067_
timestamp 1698431365
transform 1 0 28896 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2068_
timestamp 1698431365
transform 1 0 50848 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2069_
timestamp 1698431365
transform 1 0 50176 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2070_
timestamp 1698431365
transform -1 0 51968 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2071_
timestamp 1698431365
transform -1 0 50176 0 1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2072_
timestamp 1698431365
transform -1 0 46144 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2073_
timestamp 1698431365
transform -1 0 44016 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2074_
timestamp 1698431365
transform -1 0 42896 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2075_
timestamp 1698431365
transform 1 0 42672 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2076_
timestamp 1698431365
transform 1 0 41216 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2077_
timestamp 1698431365
transform 1 0 42000 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2078_
timestamp 1698431365
transform -1 0 43568 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2079_
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2080_
timestamp 1698431365
transform -1 0 48048 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2081_
timestamp 1698431365
transform -1 0 44464 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2082_
timestamp 1698431365
transform -1 0 46368 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2083_
timestamp 1698431365
transform -1 0 49504 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2084_
timestamp 1698431365
transform 1 0 47152 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2085_
timestamp 1698431365
transform -1 0 52192 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2086_
timestamp 1698431365
transform 1 0 52752 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2087_
timestamp 1698431365
transform -1 0 52192 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2088_
timestamp 1698431365
transform -1 0 51296 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2089_
timestamp 1698431365
transform -1 0 52864 0 -1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2090_
timestamp 1698431365
transform 1 0 52416 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2091_
timestamp 1698431365
transform 1 0 50624 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2092_
timestamp 1698431365
transform 1 0 47040 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2093_
timestamp 1698431365
transform 1 0 46368 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2094_
timestamp 1698431365
transform -1 0 46368 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2095_
timestamp 1698431365
transform -1 0 44800 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2096_
timestamp 1698431365
transform 1 0 46144 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2097_
timestamp 1698431365
transform 1 0 47488 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2098_
timestamp 1698431365
transform 1 0 55328 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2099_
timestamp 1698431365
transform -1 0 59472 0 1 34496
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2100_
timestamp 1698431365
transform -1 0 52080 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2101_
timestamp 1698431365
transform 1 0 49840 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2102_
timestamp 1698431365
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2103_
timestamp 1698431365
transform 1 0 48720 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2104_
timestamp 1698431365
transform 1 0 49168 0 -1 36064
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2105_
timestamp 1698431365
transform 1 0 50624 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2106_
timestamp 1698431365
transform -1 0 51856 0 1 39200
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2107_
timestamp 1698431365
transform -1 0 52304 0 1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2108_
timestamp 1698431365
transform 1 0 46144 0 1 34496
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2109_
timestamp 1698431365
transform 1 0 51520 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2110_
timestamp 1698431365
transform -1 0 52080 0 1 36064
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2111_
timestamp 1698431365
transform -1 0 46816 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2112_
timestamp 1698431365
transform -1 0 50624 0 -1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2113_
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2114_
timestamp 1698431365
transform -1 0 20944 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2115_
timestamp 1698431365
transform 1 0 19936 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2116_
timestamp 1698431365
transform -1 0 17024 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2117_
timestamp 1698431365
transform -1 0 20384 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2118_
timestamp 1698431365
transform 1 0 19152 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2119_
timestamp 1698431365
transform 1 0 22624 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2120_
timestamp 1698431365
transform 1 0 46592 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2121_
timestamp 1698431365
transform 1 0 45696 0 -1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2122_
timestamp 1698431365
transform -1 0 18928 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2123_
timestamp 1698431365
transform 1 0 12544 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2124_
timestamp 1698431365
transform 1 0 12656 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2125_
timestamp 1698431365
transform -1 0 15008 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2126_
timestamp 1698431365
transform 1 0 10304 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2127_
timestamp 1698431365
transform -1 0 14784 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2128_
timestamp 1698431365
transform -1 0 34944 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2129_
timestamp 1698431365
transform -1 0 36176 0 -1 50176
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2130_
timestamp 1698431365
transform -1 0 20720 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2131_
timestamp 1698431365
transform -1 0 16240 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2132_
timestamp 1698431365
transform -1 0 21616 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2133_
timestamp 1698431365
transform -1 0 17024 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2134_
timestamp 1698431365
transform -1 0 20944 0 1 47040
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2135_
timestamp 1698431365
transform 1 0 17360 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2136_
timestamp 1698431365
transform 1 0 18816 0 -1 45472
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2137_
timestamp 1698431365
transform -1 0 22624 0 -1 47040
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2138_
timestamp 1698431365
transform 1 0 13328 0 -1 48608
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2139_
timestamp 1698431365
transform -1 0 15904 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2140_
timestamp 1698431365
transform -1 0 19936 0 1 48608
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2141_
timestamp 1698431365
transform -1 0 22624 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2142_
timestamp 1698431365
transform 1 0 41552 0 -1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2143_
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2144_
timestamp 1698431365
transform 1 0 47152 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2145_
timestamp 1698431365
transform -1 0 45360 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2146_
timestamp 1698431365
transform -1 0 48384 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2147_
timestamp 1698431365
transform -1 0 48272 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2148_
timestamp 1698431365
transform -1 0 44016 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2149_
timestamp 1698431365
transform 1 0 38304 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2150_
timestamp 1698431365
transform 1 0 42560 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2151_
timestamp 1698431365
transform -1 0 46816 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2152_
timestamp 1698431365
transform -1 0 43120 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2153_
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2154_
timestamp 1698431365
transform -1 0 13104 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2155_
timestamp 1698431365
transform -1 0 13104 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2156_
timestamp 1698431365
transform -1 0 13888 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2157_
timestamp 1698431365
transform -1 0 13328 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2158_
timestamp 1698431365
transform 1 0 11648 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2159_
timestamp 1698431365
transform -1 0 15008 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2160_
timestamp 1698431365
transform 1 0 40768 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2161_
timestamp 1698431365
transform 1 0 51184 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2162_
timestamp 1698431365
transform 1 0 45808 0 1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2163_
timestamp 1698431365
transform 1 0 34496 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2164_
timestamp 1698431365
transform -1 0 34048 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2165_
timestamp 1698431365
transform 1 0 39088 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2166_
timestamp 1698431365
transform 1 0 37408 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2167_
timestamp 1698431365
transform -1 0 39536 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2168_
timestamp 1698431365
transform 1 0 38640 0 1 43904
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2169_
timestamp 1698431365
transform -1 0 42336 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2170_
timestamp 1698431365
transform 1 0 13328 0 -1 45472
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2171_
timestamp 1698431365
transform -1 0 40544 0 1 42336
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2172_
timestamp 1698431365
transform 1 0 43680 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2173_
timestamp 1698431365
transform 1 0 32928 0 1 43904
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2174_
timestamp 1698431365
transform -1 0 39536 0 -1 45472
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2175_
timestamp 1698431365
transform -1 0 42224 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2176_
timestamp 1698431365
transform 1 0 41552 0 -1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2177_
timestamp 1698431365
transform 1 0 43680 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2178_
timestamp 1698431365
transform 1 0 44016 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2179_
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2180_
timestamp 1698431365
transform 1 0 43568 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2181_
timestamp 1698431365
transform -1 0 42896 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2182_
timestamp 1698431365
transform 1 0 42448 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2183_
timestamp 1698431365
transform 1 0 36960 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2184_
timestamp 1698431365
transform -1 0 38304 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2185_
timestamp 1698431365
transform 1 0 39536 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2186_
timestamp 1698431365
transform -1 0 36176 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2187_
timestamp 1698431365
transform -1 0 41440 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2188_
timestamp 1698431365
transform -1 0 41664 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2189_
timestamp 1698431365
transform -1 0 34496 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2190_
timestamp 1698431365
transform -1 0 36176 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2191_
timestamp 1698431365
transform 1 0 36512 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2192_
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2193_
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2194_
timestamp 1698431365
transform -1 0 36624 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2195_
timestamp 1698431365
transform 1 0 35840 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2196_
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2197_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2198_
timestamp 1698431365
transform 1 0 35952 0 -1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2199_
timestamp 1698431365
transform -1 0 36624 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2200_
timestamp 1698431365
transform -1 0 35728 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2201_
timestamp 1698431365
transform 1 0 39536 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2202_
timestamp 1698431365
transform 1 0 39088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2203_
timestamp 1698431365
transform 1 0 38192 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2204_
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2205_
timestamp 1698431365
transform -1 0 47488 0 -1 36064
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2206_
timestamp 1698431365
transform 1 0 43344 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2207_
timestamp 1698431365
transform 1 0 37408 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2208_
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2209_
timestamp 1698431365
transform -1 0 37408 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2210_
timestamp 1698431365
transform -1 0 39424 0 -1 36064
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2211_
timestamp 1698431365
transform 1 0 34160 0 -1 39200
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2212_
timestamp 1698431365
transform 1 0 34832 0 -1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2213_
timestamp 1698431365
transform 1 0 38080 0 1 32928
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2214_
timestamp 1698431365
transform 1 0 44128 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2215_
timestamp 1698431365
transform 1 0 37968 0 1 34496
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2216_
timestamp 1698431365
transform 1 0 35392 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2217_
timestamp 1698431365
transform 1 0 33712 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2218_
timestamp 1698431365
transform 1 0 6608 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2219_
timestamp 1698431365
transform -1 0 7280 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2220_
timestamp 1698431365
transform -1 0 5264 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2221_
timestamp 1698431365
transform 1 0 6160 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2222_
timestamp 1698431365
transform 1 0 6608 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2223_
timestamp 1698431365
transform -1 0 8624 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2224_
timestamp 1698431365
transform 1 0 8176 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2225_
timestamp 1698431365
transform -1 0 10416 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2226_
timestamp 1698431365
transform -1 0 34496 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2227_
timestamp 1698431365
transform -1 0 36288 0 1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2228_
timestamp 1698431365
transform -1 0 8960 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2229_
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2230_
timestamp 1698431365
transform -1 0 2912 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2231_
timestamp 1698431365
transform 1 0 9744 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2232_
timestamp 1698431365
transform 1 0 11648 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2233_
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2234_
timestamp 1698431365
transform -1 0 8064 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2235_
timestamp 1698431365
transform 1 0 4816 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2236_
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2237_
timestamp 1698431365
transform 1 0 7504 0 1 42336
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2238_
timestamp 1698431365
transform 1 0 7504 0 1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2239_
timestamp 1698431365
transform 1 0 6608 0 -1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2240_
timestamp 1698431365
transform -1 0 6384 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2241_
timestamp 1698431365
transform 1 0 5712 0 -1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2242_
timestamp 1698431365
transform 1 0 8512 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2243_
timestamp 1698431365
transform 1 0 4928 0 -1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2244_
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2245_
timestamp 1698431365
transform -1 0 10864 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2246_
timestamp 1698431365
transform 1 0 26768 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2247_
timestamp 1698431365
transform -1 0 32816 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2248_
timestamp 1698431365
transform 1 0 31472 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2249_
timestamp 1698431365
transform -1 0 33600 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2250_
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2251_
timestamp 1698431365
transform -1 0 42224 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2252_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30688 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2253_
timestamp 1698431365
transform -1 0 32032 0 1 40768
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2254_
timestamp 1698431365
transform 1 0 30352 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2255_
timestamp 1698431365
transform 1 0 31248 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2256_
timestamp 1698431365
transform 1 0 30128 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2257_
timestamp 1698431365
transform 1 0 29232 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2258_
timestamp 1698431365
transform -1 0 23856 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2259_
timestamp 1698431365
transform -1 0 20160 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2260_
timestamp 1698431365
transform 1 0 27328 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2261_
timestamp 1698431365
transform 1 0 29120 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2262_
timestamp 1698431365
transform -1 0 34720 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2263_
timestamp 1698431365
transform 1 0 26880 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2264_
timestamp 1698431365
transform 1 0 19376 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2265_
timestamp 1698431365
transform 1 0 27664 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2266_
timestamp 1698431365
transform -1 0 30464 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2267_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27328 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2268_
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2269_
timestamp 1698431365
transform 1 0 16128 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2270_
timestamp 1698431365
transform -1 0 28896 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2271_
timestamp 1698431365
transform -1 0 24864 0 -1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2272_
timestamp 1698431365
transform -1 0 24752 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2273_
timestamp 1698431365
transform -1 0 30688 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2274_
timestamp 1698431365
transform 1 0 20272 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2275_
timestamp 1698431365
transform 1 0 22064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2276_
timestamp 1698431365
transform -1 0 28784 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2277_
timestamp 1698431365
transform 1 0 25648 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2278_
timestamp 1698431365
transform 1 0 23632 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2279_
timestamp 1698431365
transform 1 0 20720 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2280_
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2281_
timestamp 1698431365
transform 1 0 23184 0 -1 59584
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2282_
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2283_
timestamp 1698431365
transform -1 0 32928 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2284_
timestamp 1698431365
transform -1 0 59808 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2285_
timestamp 1698431365
transform 1 0 55328 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2286_
timestamp 1698431365
transform 1 0 54656 0 1 51744
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2287_
timestamp 1698431365
transform -1 0 59136 0 1 54880
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2288_
timestamp 1698431365
transform -1 0 58912 0 1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2289_
timestamp 1698431365
transform 1 0 32928 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2290_
timestamp 1698431365
transform -1 0 28784 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2291_
timestamp 1698431365
transform 1 0 20048 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2292_
timestamp 1698431365
transform -1 0 28672 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2293_
timestamp 1698431365
transform -1 0 26320 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2294_
timestamp 1698431365
transform -1 0 22848 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2295_
timestamp 1698431365
transform 1 0 27776 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2296_
timestamp 1698431365
transform 1 0 23968 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2297_
timestamp 1698431365
transform -1 0 25984 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2298_
timestamp 1698431365
transform -1 0 37072 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2299_
timestamp 1698431365
transform 1 0 34272 0 -1 56448
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2300_
timestamp 1698431365
transform -1 0 25984 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2301_
timestamp 1698431365
transform 1 0 23184 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2302_
timestamp 1698431365
transform -1 0 23184 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2303_
timestamp 1698431365
transform 1 0 23856 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2304_
timestamp 1698431365
transform -1 0 22512 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2305_
timestamp 1698431365
transform -1 0 20944 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2306_
timestamp 1698431365
transform -1 0 21168 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2307_
timestamp 1698431365
transform -1 0 17024 0 -1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2308_
timestamp 1698431365
transform -1 0 18368 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2309_
timestamp 1698431365
transform -1 0 19936 0 -1 56448
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2310_
timestamp 1698431365
transform -1 0 20048 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2311_
timestamp 1698431365
transform -1 0 23184 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2312_
timestamp 1698431365
transform 1 0 18368 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2313_
timestamp 1698431365
transform -1 0 27776 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2314_
timestamp 1698431365
transform -1 0 24416 0 -1 54880
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2315_
timestamp 1698431365
transform -1 0 27664 0 1 50176
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2316_
timestamp 1698431365
transform 1 0 23408 0 1 53312
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2317_
timestamp 1698431365
transform -1 0 24416 0 -1 50176
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2318_
timestamp 1698431365
transform -1 0 18032 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2319_
timestamp 1698431365
transform -1 0 24864 0 -1 53312
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2320_
timestamp 1698431365
transform 1 0 25088 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2321_
timestamp 1698431365
transform -1 0 27216 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2322_
timestamp 1698431365
transform 1 0 33600 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2323_
timestamp 1698431365
transform 1 0 29568 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2324_
timestamp 1698431365
transform -1 0 32704 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2325_
timestamp 1698431365
transform -1 0 32144 0 -1 51744
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2326_
timestamp 1698431365
transform -1 0 29904 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2327_
timestamp 1698431365
transform -1 0 31920 0 -1 54880
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2328_
timestamp 1698431365
transform -1 0 28672 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2329_
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2330_
timestamp 1698431365
transform 1 0 29904 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2331_
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2332_
timestamp 1698431365
transform -1 0 32704 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2333_
timestamp 1698431365
transform 1 0 27104 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2334_
timestamp 1698431365
transform -1 0 31808 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2335_
timestamp 1698431365
transform -1 0 41664 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2336_
timestamp 1698431365
transform -1 0 31136 0 1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2337_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31136 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2338_
timestamp 1698431365
transform -1 0 30800 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2339_
timestamp 1698431365
transform -1 0 31024 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2340_
timestamp 1698431365
transform -1 0 32704 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2341_
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2342_
timestamp 1698431365
transform -1 0 26992 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2343_
timestamp 1698431365
transform -1 0 45584 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2344_
timestamp 1698431365
transform -1 0 45584 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2345_
timestamp 1698431365
transform -1 0 48384 0 -1 50176
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2346_
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2347_
timestamp 1698431365
transform -1 0 42784 0 -1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2348_
timestamp 1698431365
transform -1 0 20944 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2349_
timestamp 1698431365
transform -1 0 25984 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2350_
timestamp 1698431365
transform -1 0 22176 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2351_
timestamp 1698431365
transform -1 0 21840 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2352_
timestamp 1698431365
transform 1 0 22736 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2353_
timestamp 1698431365
transform -1 0 11088 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2354_
timestamp 1698431365
transform 1 0 11088 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2355_
timestamp 1698431365
transform -1 0 22736 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2356_
timestamp 1698431365
transform 1 0 20048 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2357_
timestamp 1698431365
transform -1 0 40096 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2358_
timestamp 1698431365
transform -1 0 41776 0 1 48608
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2359_
timestamp 1698431365
transform -1 0 24864 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2360_
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2361_
timestamp 1698431365
transform -1 0 21056 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2362_
timestamp 1698431365
transform 1 0 18592 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2363_
timestamp 1698431365
transform 1 0 16128 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2364_
timestamp 1698431365
transform -1 0 18592 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2365_
timestamp 1698431365
transform 1 0 23632 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2366_
timestamp 1698431365
transform 1 0 22512 0 1 48608
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2367_
timestamp 1698431365
transform -1 0 23296 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2368_
timestamp 1698431365
transform -1 0 22736 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2369_
timestamp 1698431365
transform 1 0 22400 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2370_
timestamp 1698431365
transform 1 0 23408 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2371_
timestamp 1698431365
transform 1 0 23296 0 1 39200
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2372_
timestamp 1698431365
transform -1 0 27328 0 1 36064
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2373_
timestamp 1698431365
transform -1 0 27440 0 1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2374_
timestamp 1698431365
transform 1 0 20048 0 -1 40768
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2375_
timestamp 1698431365
transform -1 0 20944 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2376_
timestamp 1698431365
transform -1 0 25984 0 1 40768
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2377_
timestamp 1698431365
transform -1 0 26880 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2378_
timestamp 1698431365
transform 1 0 32928 0 1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2379_
timestamp 1698431365
transform -1 0 39088 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2380_
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2381_
timestamp 1698431365
transform -1 0 36512 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2382_
timestamp 1698431365
transform -1 0 30016 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2383_
timestamp 1698431365
transform 1 0 30464 0 -1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2384_
timestamp 1698431365
transform 1 0 17472 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2385_
timestamp 1698431365
transform 1 0 17472 0 -1 48608
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2386_
timestamp 1698431365
transform -1 0 19264 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2387_
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2388_
timestamp 1698431365
transform 1 0 34496 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2389_
timestamp 1698431365
transform 1 0 36624 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2390_
timestamp 1698431365
transform 1 0 35616 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2391_
timestamp 1698431365
transform 1 0 34944 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2392_
timestamp 1698431365
transform 1 0 13216 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2393_
timestamp 1698431365
transform 1 0 34384 0 1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2394_
timestamp 1698431365
transform 1 0 12432 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2395_
timestamp 1698431365
transform 1 0 15904 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2396_
timestamp 1698431365
transform -1 0 17024 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2397_
timestamp 1698431365
transform 1 0 8512 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2398_
timestamp 1698431365
transform -1 0 21280 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2399_
timestamp 1698431365
transform 1 0 13552 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2400_
timestamp 1698431365
transform 1 0 15568 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2401_
timestamp 1698431365
transform -1 0 13776 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2402_
timestamp 1698431365
transform -1 0 43232 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2403_
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2404_
timestamp 1698431365
transform -1 0 40544 0 -1 43904
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2405_
timestamp 1698431365
transform -1 0 41552 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2406_
timestamp 1698431365
transform -1 0 40544 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2407_
timestamp 1698431365
transform -1 0 10976 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2408_
timestamp 1698431365
transform 1 0 13552 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2409_
timestamp 1698431365
transform 1 0 12096 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2410_
timestamp 1698431365
transform -1 0 16576 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2411_
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2412_
timestamp 1698431365
transform 1 0 11424 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2413_
timestamp 1698431365
transform -1 0 14784 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2414_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16128 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2415_
timestamp 1698431365
transform -1 0 14448 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2416_
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2417_
timestamp 1698431365
transform -1 0 16016 0 1 45472
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2418_
timestamp 1698431365
transform 1 0 13216 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2419_
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2420_
timestamp 1698431365
transform 1 0 9632 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2421_
timestamp 1698431365
transform -1 0 9184 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2422_
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2423_
timestamp 1698431365
transform 1 0 11200 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2424_
timestamp 1698431365
transform 1 0 16128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2425_
timestamp 1698431365
transform -1 0 20944 0 1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2426_
timestamp 1698431365
transform 1 0 10080 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2427_
timestamp 1698431365
transform -1 0 12320 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2428_
timestamp 1698431365
transform -1 0 9968 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2429_
timestamp 1698431365
transform 1 0 8848 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2430_
timestamp 1698431365
transform 1 0 11648 0 -1 37632
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2431_
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2432_
timestamp 1698431365
transform -1 0 17024 0 1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2433_
timestamp 1698431365
transform 1 0 9408 0 1 36064
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2434_
timestamp 1698431365
transform -1 0 9408 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2435_
timestamp 1698431365
transform -1 0 16016 0 -1 39200
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2436_
timestamp 1698431365
transform 1 0 12208 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2437_
timestamp 1698431365
transform -1 0 12544 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2438_
timestamp 1698431365
transform -1 0 11536 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2439_
timestamp 1698431365
transform -1 0 11424 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2440_
timestamp 1698431365
transform 1 0 7392 0 1 43904
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2441_
timestamp 1698431365
transform -1 0 9520 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2442_
timestamp 1698431365
transform 1 0 8960 0 1 47040
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2443_
timestamp 1698431365
transform 1 0 13440 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2444_
timestamp 1698431365
transform -1 0 15680 0 1 47040
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2445_
timestamp 1698431365
transform -1 0 9184 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2446_
timestamp 1698431365
transform 1 0 10304 0 -1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2447_
timestamp 1698431365
transform -1 0 12656 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2448_
timestamp 1698431365
transform 1 0 11088 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2449_
timestamp 1698431365
transform -1 0 10752 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2450_
timestamp 1698431365
transform -1 0 9184 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2451_
timestamp 1698431365
transform 1 0 45024 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2452_
timestamp 1698431365
transform -1 0 5488 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2453_
timestamp 1698431365
transform 1 0 6944 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2454_
timestamp 1698431365
transform 1 0 23968 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2455_
timestamp 1698431365
transform -1 0 8512 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2456_
timestamp 1698431365
transform -1 0 7392 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2457_
timestamp 1698431365
transform 1 0 3136 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2458_
timestamp 1698431365
transform 1 0 3696 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2459_
timestamp 1698431365
transform 1 0 33824 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2460_
timestamp 1698431365
transform 1 0 25536 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2461_
timestamp 1698431365
transform -1 0 32144 0 -1 37632
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2462_
timestamp 1698431365
transform -1 0 32256 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2463_
timestamp 1698431365
transform -1 0 5264 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2464_
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2465_
timestamp 1698431365
transform -1 0 6160 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2466_
timestamp 1698431365
transform -1 0 3248 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2467_
timestamp 1698431365
transform 1 0 8960 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2468_
timestamp 1698431365
transform -1 0 12544 0 1 34496
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2469_
timestamp 1698431365
transform -1 0 7616 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2470_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2471_
timestamp 1698431365
transform -1 0 2912 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2472_
timestamp 1698431365
transform -1 0 9072 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2473_
timestamp 1698431365
transform -1 0 6496 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2474_
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2475_
timestamp 1698431365
transform -1 0 6384 0 -1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2476_
timestamp 1698431365
transform -1 0 6944 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2477_
timestamp 1698431365
transform -1 0 5824 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2478_
timestamp 1698431365
transform 1 0 4032 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2479_
timestamp 1698431365
transform -1 0 3696 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2480_
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2481_
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2482_
timestamp 1698431365
transform 1 0 2800 0 -1 31360
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2483_
timestamp 1698431365
transform -1 0 3360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2484_
timestamp 1698431365
transform 1 0 4144 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2485_
timestamp 1698431365
transform 1 0 4256 0 -1 32928
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2486_
timestamp 1698431365
transform 1 0 2688 0 -1 36064
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2487_
timestamp 1698431365
transform 1 0 6720 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2488_
timestamp 1698431365
transform 1 0 2800 0 -1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2489_
timestamp 1698431365
transform 1 0 1792 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2490_
timestamp 1698431365
transform -1 0 4816 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2491_
timestamp 1698431365
transform 1 0 3920 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2492_
timestamp 1698431365
transform 1 0 3024 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2493_
timestamp 1698431365
transform 1 0 2128 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2494_
timestamp 1698431365
transform -1 0 8960 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2495_
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2496_
timestamp 1698431365
transform 1 0 2912 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2497_
timestamp 1698431365
transform -1 0 3024 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2498_
timestamp 1698431365
transform -1 0 26320 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2499_
timestamp 1698431365
transform 1 0 4032 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2500_
timestamp 1698431365
transform 1 0 4032 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2501_
timestamp 1698431365
transform -1 0 12992 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2502_
timestamp 1698431365
transform -1 0 4144 0 -1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2503_
timestamp 1698431365
transform 1 0 23184 0 -1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2504_
timestamp 1698431365
transform -1 0 20944 0 1 56448
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2505_
timestamp 1698431365
transform 1 0 13664 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2506_
timestamp 1698431365
transform -1 0 14560 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2507_
timestamp 1698431365
transform 1 0 11984 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2508_
timestamp 1698431365
transform 1 0 13216 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2509_
timestamp 1698431365
transform -1 0 19936 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2510_
timestamp 1698431365
transform 1 0 18480 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2511_
timestamp 1698431365
transform -1 0 12992 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2512_
timestamp 1698431365
transform -1 0 15232 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2513_
timestamp 1698431365
transform 1 0 14896 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2514_
timestamp 1698431365
transform -1 0 20832 0 1 58016
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2515_
timestamp 1698431365
transform 1 0 13888 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2516_
timestamp 1698431365
transform -1 0 21840 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2517_
timestamp 1698431365
transform 1 0 20944 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2518_
timestamp 1698431365
transform -1 0 18256 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2519_
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2520_
timestamp 1698431365
transform -1 0 5936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2521_
timestamp 1698431365
transform -1 0 5264 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2522_
timestamp 1698431365
transform 1 0 4480 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2523_
timestamp 1698431365
transform 1 0 3920 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2524_
timestamp 1698431365
transform -1 0 8176 0 1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2525_
timestamp 1698431365
transform 1 0 12880 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2526_
timestamp 1698431365
transform 1 0 14224 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2527_
timestamp 1698431365
transform 1 0 11200 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2528_
timestamp 1698431365
transform 1 0 12320 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2529_
timestamp 1698431365
transform -1 0 17248 0 1 31360
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2530_
timestamp 1698431365
transform -1 0 16128 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2531_
timestamp 1698431365
transform -1 0 18704 0 1 28224
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2532_
timestamp 1698431365
transform -1 0 18256 0 1 29792
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2533_
timestamp 1698431365
transform 1 0 16128 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2534_
timestamp 1698431365
transform -1 0 20944 0 -1 32928
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2535_
timestamp 1698431365
transform -1 0 11312 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2536_
timestamp 1698431365
transform 1 0 14448 0 1 32928
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2537_
timestamp 1698431365
transform -1 0 16016 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2538_
timestamp 1698431365
transform 1 0 14672 0 1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2539_
timestamp 1698431365
transform 1 0 11984 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2540_
timestamp 1698431365
transform 1 0 16688 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2541_
timestamp 1698431365
transform -1 0 15344 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2542_
timestamp 1698431365
transform 1 0 3360 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2543_
timestamp 1698431365
transform -1 0 9072 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2544_
timestamp 1698431365
transform -1 0 5264 0 1 31360
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2545_
timestamp 1698431365
transform 1 0 1904 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2546_
timestamp 1698431365
transform 1 0 6832 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2547_
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2548_
timestamp 1698431365
transform 1 0 15008 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2549_
timestamp 1698431365
transform 1 0 21728 0 1 51744
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2550_
timestamp 1698431365
transform 1 0 20944 0 -1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2551_
timestamp 1698431365
transform -1 0 20720 0 -1 54880
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2552_
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2553_
timestamp 1698431365
transform -1 0 14000 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2554_
timestamp 1698431365
transform -1 0 15568 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2555_
timestamp 1698431365
transform 1 0 15568 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2556_
timestamp 1698431365
transform 1 0 12992 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2557_
timestamp 1698431365
transform 1 0 14896 0 -1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2558_
timestamp 1698431365
transform 1 0 15344 0 -1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2559_
timestamp 1698431365
transform 1 0 14224 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2560_
timestamp 1698431365
transform -1 0 22288 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2561_
timestamp 1698431365
transform -1 0 24976 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2562_
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2563_
timestamp 1698431365
transform -1 0 21728 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2564_
timestamp 1698431365
transform 1 0 20272 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2565_
timestamp 1698431365
transform 1 0 34832 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2566_
timestamp 1698431365
transform -1 0 30240 0 -1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2567_
timestamp 1698431365
transform -1 0 30800 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2568_
timestamp 1698431365
transform -1 0 29904 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2569_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2570_
timestamp 1698431365
transform 1 0 31920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2571_
timestamp 1698431365
transform -1 0 36400 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2572_
timestamp 1698431365
transform 1 0 32928 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2573_
timestamp 1698431365
transform 1 0 31024 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2574_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2575_
timestamp 1698431365
transform 1 0 27888 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2576_
timestamp 1698431365
transform -1 0 31136 0 -1 47040
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2577_
timestamp 1698431365
transform 1 0 29904 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2578_
timestamp 1698431365
transform 1 0 17472 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2579_
timestamp 1698431365
transform -1 0 13664 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2580_
timestamp 1698431365
transform 1 0 19600 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2581_
timestamp 1698431365
transform 1 0 18704 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2582_
timestamp 1698431365
transform -1 0 20944 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2583_
timestamp 1698431365
transform 1 0 18256 0 1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2584_
timestamp 1698431365
transform -1 0 24752 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2585_
timestamp 1698431365
transform -1 0 20160 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2586_
timestamp 1698431365
transform -1 0 28000 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2587_
timestamp 1698431365
transform 1 0 25872 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2588_
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2589_
timestamp 1698431365
transform 1 0 32704 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2590_
timestamp 1698431365
transform -1 0 34496 0 1 28224
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2591_
timestamp 1698431365
transform -1 0 32704 0 1 29792
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2592_
timestamp 1698431365
transform 1 0 18480 0 -1 29792
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2593_
timestamp 1698431365
transform -1 0 27888 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2594_
timestamp 1698431365
transform 1 0 21280 0 1 29792
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2595_
timestamp 1698431365
transform -1 0 28784 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2596_
timestamp 1698431365
transform -1 0 29232 0 -1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2597_
timestamp 1698431365
transform 1 0 26768 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2598_
timestamp 1698431365
transform 1 0 26432 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2599_
timestamp 1698431365
transform 1 0 23184 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2600_
timestamp 1698431365
transform -1 0 19152 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2601_
timestamp 1698431365
transform 1 0 21504 0 1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2602_
timestamp 1698431365
transform -1 0 23296 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2603_
timestamp 1698431365
transform 1 0 14784 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2604_
timestamp 1698431365
transform 1 0 22736 0 -1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2605_
timestamp 1698431365
transform 1 0 24976 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2606_
timestamp 1698431365
transform 1 0 23520 0 1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2607_
timestamp 1698431365
transform -1 0 25536 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2608_
timestamp 1698431365
transform -1 0 24864 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2609_
timestamp 1698431365
transform -1 0 26432 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2610_
timestamp 1698431365
transform 1 0 23744 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2611_
timestamp 1698431365
transform -1 0 20048 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2612_
timestamp 1698431365
transform 1 0 15120 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2613_
timestamp 1698431365
transform 1 0 22512 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2614_
timestamp 1698431365
transform -1 0 36064 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2615_
timestamp 1698431365
transform -1 0 20160 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2616_
timestamp 1698431365
transform -1 0 22288 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2617_
timestamp 1698431365
transform -1 0 24864 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2618_
timestamp 1698431365
transform 1 0 18144 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2619_
timestamp 1698431365
transform -1 0 21728 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2620_
timestamp 1698431365
transform 1 0 18368 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2621_
timestamp 1698431365
transform -1 0 16352 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2622_
timestamp 1698431365
transform -1 0 20496 0 1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2623_
timestamp 1698431365
transform 1 0 18032 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2624_
timestamp 1698431365
transform -1 0 18256 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2625_
timestamp 1698431365
transform 1 0 15792 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2626_
timestamp 1698431365
transform -1 0 18368 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2627_
timestamp 1698431365
transform -1 0 22848 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2628_
timestamp 1698431365
transform -1 0 22512 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2629_
timestamp 1698431365
transform -1 0 18592 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2630_
timestamp 1698431365
transform 1 0 18256 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2631_
timestamp 1698431365
transform -1 0 20944 0 1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2632_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2633_
timestamp 1698431365
transform 1 0 12320 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2634_
timestamp 1698431365
transform 1 0 11536 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2635_
timestamp 1698431365
transform -1 0 15008 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2636_
timestamp 1698431365
transform 1 0 12432 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2637_
timestamp 1698431365
transform 1 0 12208 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2638_
timestamp 1698431365
transform 1 0 16128 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2639_
timestamp 1698431365
transform -1 0 20048 0 -1 28224
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2640_
timestamp 1698431365
transform 1 0 15568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2641_
timestamp 1698431365
transform -1 0 16912 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2642_
timestamp 1698431365
transform -1 0 16912 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2643_
timestamp 1698431365
transform -1 0 15568 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2644_
timestamp 1698431365
transform -1 0 21168 0 -1 20384
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2645_
timestamp 1698431365
transform 1 0 20048 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2646_
timestamp 1698431365
transform -1 0 23408 0 -1 17248
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2647_
timestamp 1698431365
transform -1 0 21952 0 -1 18816
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2648_
timestamp 1698431365
transform 1 0 13328 0 -1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2649_
timestamp 1698431365
transform -1 0 15568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2650_
timestamp 1698431365
transform -1 0 19600 0 1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2651_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2652_
timestamp 1698431365
transform -1 0 19152 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2653_
timestamp 1698431365
transform -1 0 17360 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2654_
timestamp 1698431365
transform -1 0 17360 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2655_
timestamp 1698431365
transform -1 0 18144 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2656_
timestamp 1698431365
transform -1 0 26768 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2657_
timestamp 1698431365
transform -1 0 24976 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2658_
timestamp 1698431365
transform -1 0 10528 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2659_
timestamp 1698431365
transform 1 0 9520 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2660_
timestamp 1698431365
transform 1 0 10976 0 1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2661_
timestamp 1698431365
transform -1 0 14672 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2662_
timestamp 1698431365
transform 1 0 13888 0 1 39200
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2663_
timestamp 1698431365
transform 1 0 15344 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2664_
timestamp 1698431365
transform 1 0 16352 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2665_
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2666_
timestamp 1698431365
transform 1 0 15232 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2667_
timestamp 1698431365
transform -1 0 15232 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2668_
timestamp 1698431365
transform 1 0 14448 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2669_
timestamp 1698431365
transform -1 0 13328 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2670_
timestamp 1698431365
transform 1 0 15568 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2671_
timestamp 1698431365
transform -1 0 15904 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2672_
timestamp 1698431365
transform 1 0 15120 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2673_
timestamp 1698431365
transform 1 0 18144 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2674_
timestamp 1698431365
transform 1 0 6832 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2675_
timestamp 1698431365
transform 1 0 6160 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2676_
timestamp 1698431365
transform -1 0 12880 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2677_
timestamp 1698431365
transform -1 0 11536 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2678_
timestamp 1698431365
transform 1 0 10304 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2679_
timestamp 1698431365
transform -1 0 11984 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2680_
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2681_
timestamp 1698431365
transform 1 0 7952 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2682_
timestamp 1698431365
transform -1 0 12096 0 1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2683_
timestamp 1698431365
transform -1 0 6160 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2684_
timestamp 1698431365
transform -1 0 9184 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2685_
timestamp 1698431365
transform 1 0 3808 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2686_
timestamp 1698431365
transform -1 0 5040 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2687_
timestamp 1698431365
transform -1 0 10976 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2688_
timestamp 1698431365
transform 1 0 11648 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2689_
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2690_
timestamp 1698431365
transform -1 0 7616 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2691_
timestamp 1698431365
transform 1 0 4928 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2692_
timestamp 1698431365
transform 1 0 5376 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2693_
timestamp 1698431365
transform 1 0 7056 0 1 17248
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2694_
timestamp 1698431365
transform -1 0 11536 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2695_
timestamp 1698431365
transform -1 0 11424 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2696_
timestamp 1698431365
transform 1 0 9856 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2697_
timestamp 1698431365
transform 1 0 5040 0 -1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2698_
timestamp 1698431365
transform 1 0 5936 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2699_
timestamp 1698431365
transform -1 0 7952 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2700_
timestamp 1698431365
transform 1 0 7392 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2701_
timestamp 1698431365
transform 1 0 10080 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2702_
timestamp 1698431365
transform 1 0 7280 0 -1 29792
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2703_
timestamp 1698431365
transform -1 0 7504 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2704_
timestamp 1698431365
transform 1 0 7280 0 -1 40768
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2705_
timestamp 1698431365
transform 1 0 9744 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2706_
timestamp 1698431365
transform -1 0 9184 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2707_
timestamp 1698431365
transform -1 0 13104 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2708_
timestamp 1698431365
transform -1 0 12208 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2709_
timestamp 1698431365
transform 1 0 3696 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2710_
timestamp 1698431365
transform -1 0 7392 0 1 32928
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2711_
timestamp 1698431365
transform 1 0 7392 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2712_
timestamp 1698431365
transform -1 0 10304 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2713_
timestamp 1698431365
transform 1 0 8512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2714_
timestamp 1698431365
transform -1 0 11200 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2715_
timestamp 1698431365
transform 1 0 7616 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2716_
timestamp 1698431365
transform -1 0 8512 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2717_
timestamp 1698431365
transform 1 0 2016 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2718_
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2719_
timestamp 1698431365
transform 1 0 8848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2720_
timestamp 1698431365
transform 1 0 6720 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2721_
timestamp 1698431365
transform 1 0 11312 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2722_
timestamp 1698431365
transform 1 0 15904 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2723_
timestamp 1698431365
transform 1 0 15008 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2724_
timestamp 1698431365
transform 1 0 15568 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2725_
timestamp 1698431365
transform -1 0 25760 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2726_
timestamp 1698431365
transform -1 0 24864 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2727_
timestamp 1698431365
transform 1 0 16128 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2728_
timestamp 1698431365
transform -1 0 17808 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2729_
timestamp 1698431365
transform 1 0 11088 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2730_
timestamp 1698431365
transform 1 0 12880 0 -1 31360
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2731_
timestamp 1698431365
transform 1 0 12656 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2732_
timestamp 1698431365
transform -1 0 12992 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2733_
timestamp 1698431365
transform -1 0 23072 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2734_
timestamp 1698431365
transform 1 0 22400 0 -1 56448
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2735_
timestamp 1698431365
transform 1 0 23408 0 1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2736_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2737_
timestamp 1698431365
transform 1 0 23856 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2738_
timestamp 1698431365
transform -1 0 24864 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2739_
timestamp 1698431365
transform 1 0 41776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2740_
timestamp 1698431365
transform 1 0 44016 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2741_
timestamp 1698431365
transform 1 0 45248 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2742_
timestamp 1698431365
transform -1 0 45584 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2743_
timestamp 1698431365
transform 1 0 30240 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2744_
timestamp 1698431365
transform 1 0 26320 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2745_
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2746_
timestamp 1698431365
transform 1 0 23968 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2747_
timestamp 1698431365
transform 1 0 27104 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2748_
timestamp 1698431365
transform -1 0 29680 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2749_
timestamp 1698431365
transform 1 0 34608 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2750_
timestamp 1698431365
transform -1 0 30464 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2751_
timestamp 1698431365
transform -1 0 31024 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2752_
timestamp 1698431365
transform -1 0 21616 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2753_
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2754_
timestamp 1698431365
transform -1 0 23856 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2755_
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2756_
timestamp 1698431365
transform -1 0 24864 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2757_
timestamp 1698431365
transform 1 0 26880 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2758_
timestamp 1698431365
transform -1 0 24528 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2759_
timestamp 1698431365
transform 1 0 22064 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2760_
timestamp 1698431365
transform 1 0 26208 0 1 25088
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2761_
timestamp 1698431365
transform -1 0 30688 0 -1 26656
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2762_
timestamp 1698431365
transform 1 0 26544 0 -1 25088
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2763_
timestamp 1698431365
transform -1 0 29904 0 -1 23520
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2764_
timestamp 1698431365
transform -1 0 22512 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2765_
timestamp 1698431365
transform 1 0 25088 0 1 21952
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2766_
timestamp 1698431365
transform -1 0 25424 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2767_
timestamp 1698431365
transform -1 0 24864 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2768_
timestamp 1698431365
transform 1 0 27888 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2769_
timestamp 1698431365
transform -1 0 25872 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2770_
timestamp 1698431365
transform 1 0 25312 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2771_
timestamp 1698431365
transform 1 0 25424 0 -1 31360
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2772_
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2773_
timestamp 1698431365
transform -1 0 23408 0 -1 31360
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2774_
timestamp 1698431365
transform 1 0 11648 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2775_
timestamp 1698431365
transform 1 0 18144 0 1 32928
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2776_
timestamp 1698431365
transform 1 0 21728 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2777_
timestamp 1698431365
transform 1 0 22736 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2778_
timestamp 1698431365
transform -1 0 26208 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2779_
timestamp 1698431365
transform -1 0 26208 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2780_
timestamp 1698431365
transform 1 0 37856 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2781_
timestamp 1698431365
transform -1 0 23296 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2782_
timestamp 1698431365
transform 1 0 23856 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2783_
timestamp 1698431365
transform 1 0 21280 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2784_
timestamp 1698431365
transform 1 0 28224 0 -1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2785_
timestamp 1698431365
transform -1 0 22624 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2786_
timestamp 1698431365
transform -1 0 23856 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2787_
timestamp 1698431365
transform 1 0 22400 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2788_
timestamp 1698431365
transform -1 0 23296 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2789_
timestamp 1698431365
transform -1 0 24864 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2790_
timestamp 1698431365
transform -1 0 33824 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2791_
timestamp 1698431365
transform -1 0 28448 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2792_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2793_
timestamp 1698431365
transform -1 0 37520 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2794_
timestamp 1698431365
transform -1 0 37744 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2795_
timestamp 1698431365
transform 1 0 43680 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2796_
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2797_
timestamp 1698431365
transform -1 0 38640 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2798_
timestamp 1698431365
transform 1 0 35504 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2799_
timestamp 1698431365
transform 1 0 22960 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2800_
timestamp 1698431365
transform -1 0 26544 0 1 34496
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2801_
timestamp 1698431365
transform 1 0 28448 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2802_
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2803_
timestamp 1698431365
transform 1 0 18480 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2804_
timestamp 1698431365
transform -1 0 24304 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2805_
timestamp 1698431365
transform 1 0 23968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2806_
timestamp 1698431365
transform -1 0 26992 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2807_
timestamp 1698431365
transform -1 0 34720 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2808_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2809_
timestamp 1698431365
transform -1 0 31136 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2810_
timestamp 1698431365
transform -1 0 27888 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2811_
timestamp 1698431365
transform 1 0 27104 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2812_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2813_
timestamp 1698431365
transform 1 0 27664 0 -1 18816
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2814_
timestamp 1698431365
transform -1 0 37520 0 -1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2815_
timestamp 1698431365
transform -1 0 28784 0 1 18816
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2816_
timestamp 1698431365
transform 1 0 26096 0 -1 15680
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2817_
timestamp 1698431365
transform -1 0 23968 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2818_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2819_
timestamp 1698431365
transform 1 0 25424 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2820_
timestamp 1698431365
transform -1 0 27104 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2821_
timestamp 1698431365
transform 1 0 10528 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2822_
timestamp 1698431365
transform -1 0 13664 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2823_
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2824_
timestamp 1698431365
transform 1 0 20160 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2825_
timestamp 1698431365
transform 1 0 22176 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2826_
timestamp 1698431365
transform 1 0 15232 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2827_
timestamp 1698431365
transform -1 0 20608 0 1 18816
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2828_
timestamp 1698431365
transform 1 0 14672 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2829_
timestamp 1698431365
transform -1 0 15792 0 -1 23520
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2830_
timestamp 1698431365
transform -1 0 14448 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2831_
timestamp 1698431365
transform 1 0 16352 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2832_
timestamp 1698431365
transform -1 0 30688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2833_
timestamp 1698431365
transform 1 0 12208 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2834_
timestamp 1698431365
transform -1 0 14112 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2835_
timestamp 1698431365
transform 1 0 10976 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2836_
timestamp 1698431365
transform 1 0 11536 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2837_
timestamp 1698431365
transform 1 0 20496 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2838_
timestamp 1698431365
transform -1 0 15344 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2839_
timestamp 1698431365
transform -1 0 15904 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2840_
timestamp 1698431365
transform -1 0 19824 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2841_
timestamp 1698431365
transform -1 0 16352 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2842_
timestamp 1698431365
transform 1 0 16912 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2843_
timestamp 1698431365
transform -1 0 20832 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2844_
timestamp 1698431365
transform -1 0 13776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2845_
timestamp 1698431365
transform 1 0 12320 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2846_
timestamp 1698431365
transform -1 0 15232 0 -1 40768
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2847_
timestamp 1698431365
transform 1 0 13440 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2848_
timestamp 1698431365
transform 1 0 14784 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2849_
timestamp 1698431365
transform -1 0 20608 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2850_
timestamp 1698431365
transform -1 0 42896 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2851_
timestamp 1698431365
transform -1 0 42560 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2852_
timestamp 1698431365
transform 1 0 42784 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2853_
timestamp 1698431365
transform -1 0 40544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2854_
timestamp 1698431365
transform 1 0 23072 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2855_
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2856_
timestamp 1698431365
transform 1 0 15456 0 1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2857_
timestamp 1698431365
transform 1 0 19936 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2858_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2859_
timestamp 1698431365
transform 1 0 15792 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2860_
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2861_
timestamp 1698431365
transform 1 0 13664 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2862_
timestamp 1698431365
transform -1 0 16352 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2863_
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2864_
timestamp 1698431365
transform -1 0 27776 0 1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2865_
timestamp 1698431365
transform -1 0 17248 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2866_
timestamp 1698431365
transform -1 0 18928 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2867_
timestamp 1698431365
transform -1 0 20944 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2868_
timestamp 1698431365
transform 1 0 16464 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2869_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2870_
timestamp 1698431365
transform -1 0 24528 0 -1 7840
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2871_
timestamp 1698431365
transform -1 0 23072 0 -1 9408
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2872_
timestamp 1698431365
transform 1 0 16016 0 1 7840
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2873_
timestamp 1698431365
transform 1 0 21840 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2874_
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2875_
timestamp 1698431365
transform 1 0 17360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2876_
timestamp 1698431365
transform 1 0 16128 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2877_
timestamp 1698431365
transform -1 0 14224 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2878_
timestamp 1698431365
transform 1 0 4704 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2879_
timestamp 1698431365
transform 1 0 7056 0 1 18816
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2880_
timestamp 1698431365
transform 1 0 8288 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2881_
timestamp 1698431365
transform 1 0 11424 0 -1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2882_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2883_
timestamp 1698431365
transform -1 0 15232 0 1 18816
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2884_
timestamp 1698431365
transform -1 0 10752 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2885_
timestamp 1698431365
transform 1 0 13776 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2886_
timestamp 1698431365
transform -1 0 44016 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2887_
timestamp 1698431365
transform -1 0 17584 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2888_
timestamp 1698431365
transform -1 0 16464 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2889_
timestamp 1698431365
transform -1 0 13104 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2890_
timestamp 1698431365
transform 1 0 12432 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2891_
timestamp 1698431365
transform 1 0 8288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2892_
timestamp 1698431365
transform -1 0 8736 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2893_
timestamp 1698431365
transform -1 0 9184 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2894_
timestamp 1698431365
transform -1 0 8848 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2895_
timestamp 1698431365
transform -1 0 5936 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2896_
timestamp 1698431365
transform -1 0 4592 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2897_
timestamp 1698431365
transform 1 0 1680 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2898_
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2899_
timestamp 1698431365
transform -1 0 5264 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2900_
timestamp 1698431365
transform -1 0 5264 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2901_
timestamp 1698431365
transform -1 0 5040 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2902_
timestamp 1698431365
transform 1 0 4368 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2903_
timestamp 1698431365
transform 1 0 13776 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2904_
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2905_
timestamp 1698431365
transform -1 0 9184 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2906_
timestamp 1698431365
transform -1 0 7168 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2907_
timestamp 1698431365
transform 1 0 25424 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2908_
timestamp 1698431365
transform -1 0 27888 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2909_
timestamp 1698431365
transform 1 0 26208 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2910_
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2911_
timestamp 1698431365
transform -1 0 28784 0 1 9408
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2912_
timestamp 1698431365
transform 1 0 3696 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2913_
timestamp 1698431365
transform 1 0 2912 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2914_
timestamp 1698431365
transform -1 0 5264 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2915_
timestamp 1698431365
transform -1 0 6944 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2916_
timestamp 1698431365
transform 1 0 3920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2917_
timestamp 1698431365
transform 1 0 5824 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2918_
timestamp 1698431365
transform -1 0 9184 0 -1 12544
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2919_
timestamp 1698431365
transform 1 0 6944 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2920_
timestamp 1698431365
transform 1 0 6496 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2921_
timestamp 1698431365
transform -1 0 11200 0 1 10976
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2922_
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2923_
timestamp 1698431365
transform -1 0 4368 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2924_
timestamp 1698431365
transform -1 0 10640 0 1 14112
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2925_
timestamp 1698431365
transform -1 0 5264 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2926_
timestamp 1698431365
transform -1 0 7952 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2927_
timestamp 1698431365
transform 1 0 6608 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2928_
timestamp 1698431365
transform 1 0 6608 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2929_
timestamp 1698431365
transform -1 0 7392 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2930_
timestamp 1698431365
transform 1 0 8960 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2931_
timestamp 1698431365
transform -1 0 10080 0 1 21952
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2932_
timestamp 1698431365
transform -1 0 7392 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2933_
timestamp 1698431365
transform -1 0 6720 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2934_
timestamp 1698431365
transform -1 0 8176 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2935_
timestamp 1698431365
transform 1 0 6720 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2936_
timestamp 1698431365
transform -1 0 11536 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2937_
timestamp 1698431365
transform -1 0 8624 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2938_
timestamp 1698431365
transform -1 0 13104 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2939_
timestamp 1698431365
transform 1 0 14560 0 -1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2940_
timestamp 1698431365
transform 1 0 37968 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2941_
timestamp 1698431365
transform -1 0 40320 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2942_
timestamp 1698431365
transform 1 0 37520 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2943_
timestamp 1698431365
transform -1 0 47824 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2944_
timestamp 1698431365
transform -1 0 46704 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2945_
timestamp 1698431365
transform -1 0 40544 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2946_
timestamp 1698431365
transform 1 0 15456 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2947_
timestamp 1698431365
transform -1 0 18480 0 1 26656
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2948_
timestamp 1698431365
transform 1 0 38864 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2949_
timestamp 1698431365
transform 1 0 45584 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2950_
timestamp 1698431365
transform -1 0 44688 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2951_
timestamp 1698431365
transform 1 0 46144 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2952_
timestamp 1698431365
transform -1 0 44016 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2953_
timestamp 1698431365
transform -1 0 45584 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2954_
timestamp 1698431365
transform 1 0 31472 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2955_
timestamp 1698431365
transform -1 0 32704 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2956_
timestamp 1698431365
transform -1 0 29456 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2957_
timestamp 1698431365
transform 1 0 30016 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2958_
timestamp 1698431365
transform -1 0 34608 0 1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2959_
timestamp 1698431365
transform 1 0 39312 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2960_
timestamp 1698431365
transform 1 0 42336 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2961_
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2962_
timestamp 1698431365
transform 1 0 37856 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _2963_
timestamp 1698431365
transform -1 0 42336 0 1 25088
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2964_
timestamp 1698431365
transform -1 0 44128 0 1 28224
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2965_
timestamp 1698431365
transform -1 0 43008 0 1 26656
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2966_
timestamp 1698431365
transform -1 0 44464 0 -1 23520
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2967_
timestamp 1698431365
transform -1 0 37744 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2968_
timestamp 1698431365
transform -1 0 41440 0 1 23520
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2969_
timestamp 1698431365
transform 1 0 37184 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2970_
timestamp 1698431365
transform -1 0 39312 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2971_
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2972_
timestamp 1698431365
transform 1 0 17360 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2973_
timestamp 1698431365
transform -1 0 22064 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2974_
timestamp 1698431365
transform 1 0 11536 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2975_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2976_
timestamp 1698431365
transform 1 0 6048 0 1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2977_
timestamp 1698431365
transform -1 0 8624 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2978_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2979_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2980_
timestamp 1698431365
transform 1 0 23408 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2981_
timestamp 1698431365
transform 1 0 26096 0 1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2982_
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2983_
timestamp 1698431365
transform -1 0 25312 0 1 23520
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2984_
timestamp 1698431365
transform 1 0 19488 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2985_
timestamp 1698431365
transform -1 0 18032 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2986_
timestamp 1698431365
transform 1 0 18144 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2987_
timestamp 1698431365
transform -1 0 19376 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2988_
timestamp 1698431365
transform 1 0 22288 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2989_
timestamp 1698431365
transform -1 0 25424 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2990_
timestamp 1698431365
transform -1 0 19264 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2991_
timestamp 1698431365
transform 1 0 20160 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2992_
timestamp 1698431365
transform -1 0 20496 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2993_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2994_
timestamp 1698431365
transform -1 0 26544 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2995_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2996_
timestamp 1698431365
transform -1 0 24864 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2997_
timestamp 1698431365
transform 1 0 22512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2998_
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2999_
timestamp 1698431365
transform 1 0 30688 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3000_
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3001_
timestamp 1698431365
transform -1 0 57792 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3002_
timestamp 1698431365
transform 1 0 52864 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3003_
timestamp 1698431365
transform -1 0 56224 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3004_
timestamp 1698431365
transform -1 0 57344 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3005_
timestamp 1698431365
transform 1 0 52640 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3006_
timestamp 1698431365
transform 1 0 34384 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3007_
timestamp 1698431365
transform 1 0 31696 0 1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3008_
timestamp 1698431365
transform 1 0 49952 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _3009_
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3010_
timestamp 1698431365
transform -1 0 43680 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3011_
timestamp 1698431365
transform 1 0 46368 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3012_
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3013_
timestamp 1698431365
transform 1 0 44688 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3014_
timestamp 1698431365
transform 1 0 43456 0 -1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3015_
timestamp 1698431365
transform 1 0 49728 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3016_
timestamp 1698431365
transform 1 0 46368 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3017_
timestamp 1698431365
transform -1 0 52416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3018_
timestamp 1698431365
transform 1 0 47824 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _3019_
timestamp 1698431365
transform -1 0 52528 0 -1 23520
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3020_
timestamp 1698431365
transform -1 0 56224 0 1 23520
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3021_
timestamp 1698431365
transform -1 0 56224 0 -1 23520
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3022_
timestamp 1698431365
transform 1 0 44912 0 1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3023_
timestamp 1698431365
transform -1 0 51520 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3024_
timestamp 1698431365
transform 1 0 46032 0 1 21952
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3025_
timestamp 1698431365
transform -1 0 51296 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3026_
timestamp 1698431365
transform -1 0 51072 0 1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3027_
timestamp 1698431365
transform -1 0 33376 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3028_
timestamp 1698431365
transform 1 0 30576 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3029_
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3030_
timestamp 1698431365
transform 1 0 25312 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3031_
timestamp 1698431365
transform -1 0 26208 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3032_
timestamp 1698431365
transform -1 0 32704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3033_
timestamp 1698431365
transform -1 0 32368 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3034_
timestamp 1698431365
transform -1 0 30016 0 -1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3035_
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3036_
timestamp 1698431365
transform 1 0 30800 0 -1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3037_
timestamp 1698431365
transform 1 0 32928 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3038_
timestamp 1698431365
transform -1 0 32144 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3039_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3040_
timestamp 1698431365
transform 1 0 31472 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3041_
timestamp 1698431365
transform 1 0 30240 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3042_
timestamp 1698431365
transform 1 0 31696 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3043_
timestamp 1698431365
transform -1 0 26208 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3044_
timestamp 1698431365
transform -1 0 25088 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3045_
timestamp 1698431365
transform -1 0 24864 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3046_
timestamp 1698431365
transform -1 0 38976 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3047_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3048_
timestamp 1698431365
transform -1 0 24304 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3049_
timestamp 1698431365
transform -1 0 17024 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3050_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3051_
timestamp 1698431365
transform 1 0 52528 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3052_
timestamp 1698431365
transform -1 0 49728 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3053_
timestamp 1698431365
transform 1 0 48944 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3054_
timestamp 1698431365
transform 1 0 51296 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3055_
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3056_
timestamp 1698431365
transform 1 0 21728 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3057_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3058_
timestamp 1698431365
transform 1 0 49840 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3059_
timestamp 1698431365
transform 1 0 46032 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3060_
timestamp 1698431365
transform -1 0 48384 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3061_
timestamp 1698431365
transform -1 0 46368 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3062_
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3063_
timestamp 1698431365
transform 1 0 45584 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3064_
timestamp 1698431365
transform 1 0 46704 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3065_
timestamp 1698431365
transform 1 0 45696 0 -1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3066_
timestamp 1698431365
transform -1 0 44352 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3067_
timestamp 1698431365
transform -1 0 47040 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3068_
timestamp 1698431365
transform 1 0 47824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3069_
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _3070_
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3071_
timestamp 1698431365
transform -1 0 56000 0 -1 10976
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3072_
timestamp 1698431365
transform -1 0 52304 0 -1 10976
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3073_
timestamp 1698431365
transform -1 0 48384 0 1 7840
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3074_
timestamp 1698431365
transform -1 0 48384 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3075_
timestamp 1698431365
transform 1 0 46144 0 1 9408
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3076_
timestamp 1698431365
transform 1 0 47600 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3077_
timestamp 1698431365
transform -1 0 48384 0 -1 12544
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3078_
timestamp 1698431365
transform -1 0 26656 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3079_
timestamp 1698431365
transform -1 0 24528 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3080_
timestamp 1698431365
transform -1 0 21728 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3081_
timestamp 1698431365
transform 1 0 29568 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3082_
timestamp 1698431365
transform 1 0 30016 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3083_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3084_
timestamp 1698431365
transform 1 0 16464 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3085_
timestamp 1698431365
transform 1 0 18928 0 -1 10976
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3086_
timestamp 1698431365
transform -1 0 20608 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3087_
timestamp 1698431365
transform 1 0 19936 0 -1 12544
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3088_
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3089_
timestamp 1698431365
transform 1 0 24192 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3090_
timestamp 1698431365
transform 1 0 22624 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3091_
timestamp 1698431365
transform -1 0 22848 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3092_
timestamp 1698431365
transform 1 0 22848 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3093_
timestamp 1698431365
transform -1 0 23408 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3094_
timestamp 1698431365
transform 1 0 22848 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3095_
timestamp 1698431365
transform 1 0 18256 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3096_
timestamp 1698431365
transform -1 0 20832 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3097_
timestamp 1698431365
transform -1 0 19936 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3098_
timestamp 1698431365
transform -1 0 25536 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3099_
timestamp 1698431365
transform 1 0 21728 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3100_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3101_
timestamp 1698431365
transform -1 0 32704 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3102_
timestamp 1698431365
transform 1 0 36736 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3103_
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3104_
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3105_
timestamp 1698431365
transform -1 0 7504 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3106_
timestamp 1698431365
transform 1 0 10080 0 1 9408
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3107_
timestamp 1698431365
transform 1 0 35840 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3108_
timestamp 1698431365
transform -1 0 36624 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3109_
timestamp 1698431365
transform 1 0 30912 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3110_
timestamp 1698431365
transform -1 0 33824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3111_
timestamp 1698431365
transform -1 0 46032 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3112_
timestamp 1698431365
transform 1 0 43008 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3113_
timestamp 1698431365
transform -1 0 33600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3114_
timestamp 1698431365
transform -1 0 36288 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3115_
timestamp 1698431365
transform 1 0 39088 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3116_
timestamp 1698431365
transform 1 0 34944 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _3117_
timestamp 1698431365
transform -1 0 39088 0 -1 7840
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3118_
timestamp 1698431365
transform 1 0 36176 0 -1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3119_
timestamp 1698431365
transform -1 0 38864 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3120_
timestamp 1698431365
transform -1 0 32816 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3121_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3122_
timestamp 1698431365
transform -1 0 36624 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3123_
timestamp 1698431365
transform 1 0 32816 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3124_
timestamp 1698431365
transform -1 0 32704 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3125_
timestamp 1698431365
transform 1 0 33040 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3126_
timestamp 1698431365
transform -1 0 16912 0 -1 10976
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3127_
timestamp 1698431365
transform 1 0 10976 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3128_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3129_
timestamp 1698431365
transform 1 0 12768 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3130_
timestamp 1698431365
transform -1 0 14336 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3131_
timestamp 1698431365
transform -1 0 23632 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3132_
timestamp 1698431365
transform -1 0 20496 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3133_
timestamp 1698431365
transform -1 0 9744 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3134_
timestamp 1698431365
transform -1 0 11536 0 -1 10976
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3135_
timestamp 1698431365
transform -1 0 13440 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3136_
timestamp 1698431365
transform -1 0 14336 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3137_
timestamp 1698431365
transform -1 0 14784 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3138_
timestamp 1698431365
transform 1 0 11536 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3139_
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3140_
timestamp 1698431365
transform 1 0 12656 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3141_
timestamp 1698431365
transform 1 0 6944 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3142_
timestamp 1698431365
transform -1 0 8736 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3143_
timestamp 1698431365
transform -1 0 6608 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3144_
timestamp 1698431365
transform -1 0 12208 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3145_
timestamp 1698431365
transform 1 0 38752 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3146_
timestamp 1698431365
transform -1 0 40544 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3147_
timestamp 1698431365
transform -1 0 40544 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3148_
timestamp 1698431365
transform 1 0 40320 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3149_
timestamp 1698431365
transform -1 0 40320 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3150_
timestamp 1698431365
transform 1 0 41440 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3151_
timestamp 1698431365
transform 1 0 41216 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3152_
timestamp 1698431365
transform 1 0 41776 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3153_
timestamp 1698431365
transform -1 0 41104 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3154_
timestamp 1698431365
transform 1 0 36512 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3155_
timestamp 1698431365
transform 1 0 38416 0 -1 25088
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3156_
timestamp 1698431365
transform 1 0 37744 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _3157_
timestamp 1698431365
transform 1 0 35728 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3158_
timestamp 1698431365
transform -1 0 46368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3159_
timestamp 1698431365
transform -1 0 26992 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3160_
timestamp 1698431365
transform -1 0 27104 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3161_
timestamp 1698431365
transform -1 0 46256 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3162_
timestamp 1698431365
transform 1 0 51632 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3163_
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3164_
timestamp 1698431365
transform 1 0 61488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3165_
timestamp 1698431365
transform -1 0 62160 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3166_
timestamp 1698431365
transform 1 0 61264 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3167_
timestamp 1698431365
transform 1 0 44912 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3168_
timestamp 1698431365
transform 1 0 43456 0 -1 28224
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3169_
timestamp 1698431365
transform 1 0 60368 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3170_
timestamp 1698431365
transform 1 0 57008 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3171_
timestamp 1698431365
transform -1 0 61264 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3172_
timestamp 1698431365
transform 1 0 60368 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3173_
timestamp 1698431365
transform -1 0 60032 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3174_
timestamp 1698431365
transform -1 0 54432 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3175_
timestamp 1698431365
transform -1 0 57456 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3176_
timestamp 1698431365
transform -1 0 53424 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3177_
timestamp 1698431365
transform -1 0 51632 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3178_
timestamp 1698431365
transform 1 0 54768 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3179_
timestamp 1698431365
transform 1 0 52080 0 -1 29792
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3180_
timestamp 1698431365
transform -1 0 61936 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3181_
timestamp 1698431365
transform -1 0 59136 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3182_
timestamp 1698431365
transform -1 0 62384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3183_
timestamp 1698431365
transform -1 0 58688 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3184_
timestamp 1698431365
transform 1 0 57792 0 -1 28224
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3185_
timestamp 1698431365
transform 1 0 58688 0 -1 32928
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3186_
timestamp 1698431365
transform 1 0 58688 0 -1 29792
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3187_
timestamp 1698431365
transform -1 0 60032 0 1 25088
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3188_
timestamp 1698431365
transform -1 0 61040 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3189_
timestamp 1698431365
transform -1 0 61600 0 -1 26656
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3190_
timestamp 1698431365
transform -1 0 57344 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3191_
timestamp 1698431365
transform -1 0 56112 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3192_
timestamp 1698431365
transform -1 0 50288 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3193_
timestamp 1698431365
transform 1 0 45808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3194_
timestamp 1698431365
transform 1 0 49280 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3195_
timestamp 1698431365
transform 1 0 49728 0 1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3196_
timestamp 1698431365
transform 1 0 45584 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3197_
timestamp 1698431365
transform -1 0 47040 0 -1 23520
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3198_
timestamp 1698431365
transform -1 0 42000 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3199_
timestamp 1698431365
transform 1 0 40880 0 -1 26656
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3200_
timestamp 1698431365
transform 1 0 49504 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3201_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3202_
timestamp 1698431365
transform -1 0 56000 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3203_
timestamp 1698431365
transform 1 0 46368 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3204_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3205_
timestamp 1698431365
transform 1 0 46928 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3206_
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3207_
timestamp 1698431365
transform -1 0 51408 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3208_
timestamp 1698431365
transform -1 0 53648 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3209_
timestamp 1698431365
transform -1 0 48160 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3210_
timestamp 1698431365
transform 1 0 40656 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3211_
timestamp 1698431365
transform -1 0 48608 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3212_
timestamp 1698431365
transform -1 0 34272 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3213_
timestamp 1698431365
transform 1 0 34608 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3214_
timestamp 1698431365
transform -1 0 57344 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3215_
timestamp 1698431365
transform -1 0 57344 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3216_
timestamp 1698431365
transform -1 0 59136 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3217_
timestamp 1698431365
transform -1 0 56224 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3218_
timestamp 1698431365
transform 1 0 54208 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3219_
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3220_
timestamp 1698431365
transform 1 0 37520 0 -1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3221_
timestamp 1698431365
transform 1 0 52528 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3222_
timestamp 1698431365
transform -1 0 54096 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3223_
timestamp 1698431365
transform 1 0 54432 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3224_
timestamp 1698431365
transform -1 0 52080 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3225_
timestamp 1698431365
transform 1 0 52752 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3226_
timestamp 1698431365
transform 1 0 54208 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3227_
timestamp 1698431365
transform -1 0 62384 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3228_
timestamp 1698431365
transform 1 0 57456 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3229_
timestamp 1698431365
transform -1 0 60032 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3230_
timestamp 1698431365
transform -1 0 56224 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3231_
timestamp 1698431365
transform 1 0 61264 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3232_
timestamp 1698431365
transform 1 0 53536 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3233_
timestamp 1698431365
transform 1 0 54096 0 -1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3234_
timestamp 1698431365
transform -1 0 58240 0 1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3235_
timestamp 1698431365
transform 1 0 54208 0 1 18816
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3236_
timestamp 1698431365
transform 1 0 53312 0 1 15680
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3237_
timestamp 1698431365
transform -1 0 58912 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3238_
timestamp 1698431365
transform -1 0 57344 0 1 14112
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3239_
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3240_
timestamp 1698431365
transform -1 0 53536 0 -1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3241_
timestamp 1698431365
transform -1 0 45136 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3242_
timestamp 1698431365
transform 1 0 43568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3243_
timestamp 1698431365
transform -1 0 46704 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3244_
timestamp 1698431365
transform -1 0 50512 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3245_
timestamp 1698431365
transform -1 0 48720 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3246_
timestamp 1698431365
transform -1 0 48944 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3247_
timestamp 1698431365
transform 1 0 46256 0 -1 9408
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3248_
timestamp 1698431365
transform -1 0 46480 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3249_
timestamp 1698431365
transform 1 0 44464 0 -1 12544
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3250_
timestamp 1698431365
transform -1 0 45808 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3251_
timestamp 1698431365
transform 1 0 46704 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3252_
timestamp 1698431365
transform -1 0 43344 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3253_
timestamp 1698431365
transform -1 0 45808 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3254_
timestamp 1698431365
transform -1 0 40880 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3255_
timestamp 1698431365
transform 1 0 39312 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3256_
timestamp 1698431365
transform -1 0 47712 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3257_
timestamp 1698431365
transform 1 0 46368 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3258_
timestamp 1698431365
transform 1 0 47824 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3259_
timestamp 1698431365
transform -1 0 49504 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3260_
timestamp 1698431365
transform 1 0 45584 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3261_
timestamp 1698431365
transform 1 0 37856 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3262_
timestamp 1698431365
transform 1 0 46704 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3263_
timestamp 1698431365
transform -1 0 47712 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3264_
timestamp 1698431365
transform -1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3265_
timestamp 1698431365
transform -1 0 17136 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3266_
timestamp 1698431365
transform 1 0 17136 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3267_
timestamp 1698431365
transform -1 0 42896 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3268_
timestamp 1698431365
transform 1 0 40880 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3269_
timestamp 1698431365
transform 1 0 40992 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3270_
timestamp 1698431365
transform -1 0 44016 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3271_
timestamp 1698431365
transform -1 0 44352 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3272_
timestamp 1698431365
transform 1 0 43456 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3273_
timestamp 1698431365
transform 1 0 41776 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3274_
timestamp 1698431365
transform 1 0 41552 0 1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3275_
timestamp 1698431365
transform -1 0 44464 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3276_
timestamp 1698431365
transform -1 0 43456 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _3277_
timestamp 1698431365
transform 1 0 37968 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3278_
timestamp 1698431365
transform -1 0 37744 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3279_
timestamp 1698431365
transform -1 0 40320 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3280_
timestamp 1698431365
transform -1 0 37744 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3281_
timestamp 1698431365
transform 1 0 38528 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3282_
timestamp 1698431365
transform 1 0 39648 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3283_
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3284_
timestamp 1698431365
transform 1 0 53200 0 -1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3285_
timestamp 1698431365
transform -1 0 46816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3286_
timestamp 1698431365
transform -1 0 40544 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _3287_
timestamp 1698431365
transform 1 0 46928 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3288_
timestamp 1698431365
transform 1 0 40880 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3289_
timestamp 1698431365
transform 1 0 41888 0 1 14112
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3290_
timestamp 1698431365
transform -1 0 45920 0 -1 17248
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3291_
timestamp 1698431365
transform -1 0 45920 0 -1 15680
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3292_
timestamp 1698431365
transform 1 0 39424 0 1 12544
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3293_
timestamp 1698431365
transform -1 0 42336 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _3294_
timestamp 1698431365
transform -1 0 45136 0 -1 14112
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3295_
timestamp 1698431365
transform 1 0 42560 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3296_
timestamp 1698431365
transform 1 0 41664 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3297_
timestamp 1698431365
transform 1 0 40880 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3298_
timestamp 1698431365
transform -1 0 35056 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _3299_
timestamp 1698431365
transform -1 0 39424 0 -1 6272
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3300_
timestamp 1698431365
transform -1 0 35840 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3301_
timestamp 1698431365
transform 1 0 38864 0 1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3302_
timestamp 1698431365
transform -1 0 44464 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3303_
timestamp 1698431365
transform -1 0 45808 0 -1 9408
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3304_
timestamp 1698431365
transform -1 0 41664 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3305_
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3306_
timestamp 1698431365
transform 1 0 41552 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3307_
timestamp 1698431365
transform -1 0 43344 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3308_
timestamp 1698431365
transform -1 0 41664 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3309_
timestamp 1698431365
transform -1 0 40544 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3310_
timestamp 1698431365
transform -1 0 40544 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3311_
timestamp 1698431365
transform -1 0 32704 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3312_
timestamp 1698431365
transform 1 0 34832 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3313_
timestamp 1698431365
transform -1 0 36176 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3314_
timestamp 1698431365
transform 1 0 39088 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3315_
timestamp 1698431365
transform -1 0 38640 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3316_
timestamp 1698431365
transform 1 0 39424 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3317_
timestamp 1698431365
transform -1 0 11088 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3318_
timestamp 1698431365
transform 1 0 23744 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _3319_
timestamp 1698431365
transform -1 0 26096 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3320_
timestamp 1698431365
transform -1 0 27440 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3321_
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3322_
timestamp 1698431365
transform 1 0 37744 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3323_
timestamp 1698431365
transform -1 0 40432 0 1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3324_
timestamp 1698431365
transform -1 0 33376 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3325_
timestamp 1698431365
transform 1 0 30576 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3326_
timestamp 1698431365
transform -1 0 33488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _3327_
timestamp 1698431365
transform 1 0 29568 0 1 32928
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3328_
timestamp 1698431365
transform 1 0 27552 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3329_
timestamp 1698431365
transform 1 0 26992 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3330_
timestamp 1698431365
transform -1 0 24864 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3331_
timestamp 1698431365
transform -1 0 28672 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3332_
timestamp 1698431365
transform -1 0 29456 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3333_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3334_
timestamp 1698431365
transform 1 0 29904 0 -1 14112
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3335_
timestamp 1698431365
transform 1 0 31920 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _3336_
timestamp 1698431365
transform -1 0 31920 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _3337_
timestamp 1698431365
transform -1 0 34832 0 1 12544
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _3338_
timestamp 1698431365
transform 1 0 26656 0 -1 10976
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3339_
timestamp 1698431365
transform -1 0 27888 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _3340_
timestamp 1698431365
transform 1 0 28560 0 -1 12544
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3341_
timestamp 1698431365
transform -1 0 31920 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3342_
timestamp 1698431365
transform -1 0 31024 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3343_
timestamp 1698431365
transform -1 0 31920 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3344_
timestamp 1698431365
transform 1 0 28672 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3345_
timestamp 1698431365
transform -1 0 31472 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3346_
timestamp 1698431365
transform 1 0 33936 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3347_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3348_
timestamp 1698431365
transform 1 0 29344 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3349_
timestamp 1698431365
transform -1 0 28672 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3350_
timestamp 1698431365
transform 1 0 29568 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3351_
timestamp 1698431365
transform -1 0 28448 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3352_
timestamp 1698431365
transform 1 0 28224 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3353_
timestamp 1698431365
transform 1 0 29344 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3354_
timestamp 1698431365
transform 1 0 51968 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3355_
timestamp 1698431365
transform 1 0 48496 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _3356_
timestamp 1698431365
transform -1 0 50624 0 1 40768
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3357_
timestamp 1698431365
transform -1 0 39536 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3358_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3359_
timestamp 1698431365
transform 1 0 50064 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3360_
timestamp 1698431365
transform -1 0 54320 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3361_
timestamp 1698431365
transform -1 0 30800 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3362_
timestamp 1698431365
transform -1 0 33488 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3363_
timestamp 1698431365
transform -1 0 32368 0 1 10976
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3364_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3365_
timestamp 1698431365
transform 1 0 32256 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3366_
timestamp 1698431365
transform -1 0 57344 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3367_
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3368_
timestamp 1698431365
transform 1 0 58016 0 1 26656
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3369_
timestamp 1698431365
transform 1 0 56448 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3370_
timestamp 1698431365
transform -1 0 56224 0 -1 28224
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3371_
timestamp 1698431365
transform 1 0 52304 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3372_
timestamp 1698431365
transform 1 0 50288 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3373_
timestamp 1698431365
transform 1 0 45920 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3374_
timestamp 1698431365
transform -1 0 54096 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3375_
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3376_
timestamp 1698431365
transform -1 0 52304 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3377_
timestamp 1698431365
transform -1 0 52304 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3378_
timestamp 1698431365
transform 1 0 50624 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3379_
timestamp 1698431365
transform 1 0 51296 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3380_
timestamp 1698431365
transform 1 0 38976 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3381_
timestamp 1698431365
transform 1 0 56672 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3382_
timestamp 1698431365
transform 1 0 60368 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3383_
timestamp 1698431365
transform 1 0 55664 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3384_
timestamp 1698431365
transform 1 0 59584 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3385_
timestamp 1698431365
transform 1 0 60368 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3386_
timestamp 1698431365
transform -1 0 61040 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3387_
timestamp 1698431365
transform 1 0 54768 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3388_
timestamp 1698431365
transform -1 0 56224 0 -1 26656
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3389_
timestamp 1698431365
transform 1 0 51072 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3390_
timestamp 1698431365
transform 1 0 51632 0 -1 25088
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3391_
timestamp 1698431365
transform 1 0 57344 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3392_
timestamp 1698431365
transform -1 0 62384 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3393_
timestamp 1698431365
transform -1 0 57568 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3394_
timestamp 1698431365
transform 1 0 57344 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3395_
timestamp 1698431365
transform -1 0 62384 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3396_
timestamp 1698431365
transform -1 0 57344 0 1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3397_
timestamp 1698431365
transform -1 0 58128 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3398_
timestamp 1698431365
transform -1 0 58688 0 -1 21952
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3399_
timestamp 1698431365
transform -1 0 59808 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3400_
timestamp 1698431365
transform -1 0 54544 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3401_
timestamp 1698431365
transform 1 0 53872 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3402_
timestamp 1698431365
transform -1 0 59360 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3403_
timestamp 1698431365
transform 1 0 54320 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3404_
timestamp 1698431365
transform 1 0 60368 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3405_
timestamp 1698431365
transform -1 0 56224 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3406_
timestamp 1698431365
transform 1 0 54096 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3407_
timestamp 1698431365
transform -1 0 57904 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3408_
timestamp 1698431365
transform 1 0 56112 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3409_
timestamp 1698431365
transform 1 0 57344 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3410_
timestamp 1698431365
transform -1 0 56000 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3411_
timestamp 1698431365
transform -1 0 51520 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3412_
timestamp 1698431365
transform 1 0 49280 0 1 17248
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3413_
timestamp 1698431365
transform -1 0 48384 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3414_
timestamp 1698431365
transform 1 0 48496 0 1 10976
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3415_
timestamp 1698431365
transform -1 0 49280 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3416_
timestamp 1698431365
transform 1 0 60368 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3417_
timestamp 1698431365
transform -1 0 59584 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3418_
timestamp 1698431365
transform 1 0 46816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3419_
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3420_
timestamp 1698431365
transform 1 0 42336 0 1 15680
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3421_
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3422_
timestamp 1698431365
transform 1 0 47376 0 1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3423_
timestamp 1698431365
transform -1 0 51408 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3424_
timestamp 1698431365
transform 1 0 49504 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3425_
timestamp 1698431365
transform 1 0 48720 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3426_
timestamp 1698431365
transform -1 0 50288 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3427_
timestamp 1698431365
transform -1 0 50064 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3428_
timestamp 1698431365
transform 1 0 50064 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3429_
timestamp 1698431365
transform 1 0 40768 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3430_
timestamp 1698431365
transform -1 0 42224 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3431_
timestamp 1698431365
transform -1 0 41664 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3432_
timestamp 1698431365
transform 1 0 38752 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3433_
timestamp 1698431365
transform -1 0 39200 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3434_
timestamp 1698431365
transform -1 0 40096 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3435_
timestamp 1698431365
transform -1 0 37744 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3436_
timestamp 1698431365
transform -1 0 34160 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3437_
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3438_
timestamp 1698431365
transform -1 0 36624 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3439_
timestamp 1698431365
transform 1 0 34832 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3440_
timestamp 1698431365
transform 1 0 34608 0 -1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3441_
timestamp 1698431365
transform 1 0 34832 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3442_
timestamp 1698431365
transform -1 0 48048 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3443_
timestamp 1698431365
transform -1 0 47600 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3444_
timestamp 1698431365
transform 1 0 34832 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3445_
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3446_
timestamp 1698431365
transform -1 0 36288 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3447_
timestamp 1698431365
transform 1 0 35504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3448_
timestamp 1698431365
transform 1 0 34608 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3449_
timestamp 1698431365
transform -1 0 37296 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3450_
timestamp 1698431365
transform -1 0 35168 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3451_
timestamp 1698431365
transform 1 0 32816 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3452_
timestamp 1698431365
transform 1 0 33376 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3453_
timestamp 1698431365
transform -1 0 26320 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3454_
timestamp 1698431365
transform -1 0 30576 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3455_
timestamp 1698431365
transform -1 0 28784 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3456_
timestamp 1698431365
transform 1 0 27888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3457_
timestamp 1698431365
transform 1 0 58240 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3458_
timestamp 1698431365
transform -1 0 53648 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3459_
timestamp 1698431365
transform -1 0 50512 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3460_
timestamp 1698431365
transform -1 0 57008 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3461_
timestamp 1698431365
transform -1 0 56000 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3462_
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3463_
timestamp 1698431365
transform -1 0 56112 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3464_
timestamp 1698431365
transform -1 0 48384 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _3465_
timestamp 1698431365
transform 1 0 50176 0 1 43904
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3466_
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _3467_
timestamp 1698431365
transform 1 0 51856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3468_
timestamp 1698431365
transform -1 0 60032 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3469_
timestamp 1698431365
transform -1 0 58128 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3470_
timestamp 1698431365
transform -1 0 57904 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3471_
timestamp 1698431365
transform -1 0 60032 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _3472_
timestamp 1698431365
transform 1 0 57008 0 -1 47040
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3473_
timestamp 1698431365
transform -1 0 56672 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3474_
timestamp 1698431365
transform -1 0 58128 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3475_
timestamp 1698431365
transform 1 0 56224 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _3476_
timestamp 1698431365
transform -1 0 60368 0 -1 39200
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3477_
timestamp 1698431365
transform -1 0 61824 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3478_
timestamp 1698431365
transform -1 0 58352 0 -1 42336
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3479_
timestamp 1698431365
transform -1 0 55216 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3480_
timestamp 1698431365
transform 1 0 53648 0 -1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3481_
timestamp 1698431365
transform 1 0 60368 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3482_
timestamp 1698431365
transform -1 0 54096 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3483_
timestamp 1698431365
transform -1 0 56224 0 -1 45472
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3484_
timestamp 1698431365
transform 1 0 53536 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3485_
timestamp 1698431365
transform 1 0 60368 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3486_
timestamp 1698431365
transform 1 0 60816 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3487_
timestamp 1698431365
transform 1 0 60368 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3488_
timestamp 1698431365
transform -1 0 55328 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3489_
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3490_
timestamp 1698431365
transform 1 0 53200 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3491_
timestamp 1698431365
transform -1 0 54432 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3492_
timestamp 1698431365
transform -1 0 54992 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3493_
timestamp 1698431365
transform 1 0 51520 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3494_
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3495_
timestamp 1698431365
transform 1 0 46928 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3496_
timestamp 1698431365
transform -1 0 54432 0 1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3497_
timestamp 1698431365
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3498_
timestamp 1698431365
transform 1 0 54320 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3499_
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _3500_
timestamp 1698431365
transform 1 0 49280 0 -1 34496
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3501_
timestamp 1698431365
transform 1 0 51520 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3502_
timestamp 1698431365
transform 1 0 53088 0 -1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3503_
timestamp 1698431365
transform -1 0 61824 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3504_
timestamp 1698431365
transform -1 0 57008 0 1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3505_
timestamp 1698431365
transform 1 0 55216 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3506_
timestamp 1698431365
transform -1 0 56112 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3507_
timestamp 1698431365
transform -1 0 53760 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3508_
timestamp 1698431365
transform 1 0 52864 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3509_
timestamp 1698431365
transform 1 0 53200 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3510_
timestamp 1698431365
transform -1 0 45584 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3511_
timestamp 1698431365
transform -1 0 48384 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3512_
timestamp 1698431365
transform -1 0 48608 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3513_
timestamp 1698431365
transform -1 0 48384 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3514_
timestamp 1698431365
transform 1 0 45584 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3515_
timestamp 1698431365
transform -1 0 46928 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3516_
timestamp 1698431365
transform -1 0 45024 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3517_
timestamp 1698431365
transform 1 0 41104 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3518_
timestamp 1698431365
transform 1 0 41888 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3519_
timestamp 1698431365
transform -1 0 40768 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3520_
timestamp 1698431365
transform 1 0 40656 0 1 39200
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3521_
timestamp 1698431365
transform -1 0 47488 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3522_
timestamp 1698431365
transform -1 0 43456 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3523_
timestamp 1698431365
transform 1 0 34944 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _3524_
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3525_
timestamp 1698431365
transform -1 0 40544 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3526_
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3527_
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3528_
timestamp 1698431365
transform 1 0 45920 0 1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3529_
timestamp 1698431365
transform -1 0 45584 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3530_
timestamp 1698431365
transform -1 0 44352 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3531_
timestamp 1698431365
transform 1 0 43008 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3532_
timestamp 1698431365
transform 1 0 41776 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3533_
timestamp 1698431365
transform -1 0 42000 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3534_
timestamp 1698431365
transform 1 0 37296 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3535_
timestamp 1698431365
transform -1 0 40544 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3536_
timestamp 1698431365
transform -1 0 36512 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3537_
timestamp 1698431365
transform 1 0 39984 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3538_
timestamp 1698431365
transform 1 0 39984 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3539_
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3540_
timestamp 1698431365
transform 1 0 30240 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3541_
timestamp 1698431365
transform -1 0 26992 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3542_
timestamp 1698431365
transform 1 0 30688 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3543_
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3544_
timestamp 1698431365
transform -1 0 34832 0 -1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3545_
timestamp 1698431365
transform 1 0 33600 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3546_
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3547_
timestamp 1698431365
transform 1 0 42672 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3548_
timestamp 1698431365
transform -1 0 39200 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3549_
timestamp 1698431365
transform -1 0 38192 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3550_
timestamp 1698431365
transform -1 0 36176 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3551_
timestamp 1698431365
transform 1 0 35728 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3552_
timestamp 1698431365
transform 1 0 32592 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3553_
timestamp 1698431365
transform 1 0 34048 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3554_
timestamp 1698431365
transform -1 0 35056 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3555_
timestamp 1698431365
transform -1 0 35728 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3556_
timestamp 1698431365
transform 1 0 34048 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3557_
timestamp 1698431365
transform 1 0 35056 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3558_
timestamp 1698431365
transform -1 0 37520 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3559_
timestamp 1698431365
transform 1 0 35504 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3560_
timestamp 1698431365
transform -1 0 36960 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3561_
timestamp 1698431365
transform 1 0 38640 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3562_
timestamp 1698431365
transform 1 0 35392 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3563_
timestamp 1698431365
transform -1 0 36288 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3564_
timestamp 1698431365
transform -1 0 35056 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3565_
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3566_
timestamp 1698431365
transform -1 0 33824 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3567_
timestamp 1698431365
transform -1 0 34384 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3568_
timestamp 1698431365
transform -1 0 32704 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3569_
timestamp 1698431365
transform -1 0 41104 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3570_
timestamp 1698431365
transform 1 0 52528 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3571_
timestamp 1698431365
transform 1 0 44464 0 -1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3572_
timestamp 1698431365
transform -1 0 48384 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3573_
timestamp 1698431365
transform 1 0 42448 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3574_
timestamp 1698431365
transform 1 0 51296 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3575_
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3576_
timestamp 1698431365
transform -1 0 52080 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3577_
timestamp 1698431365
transform -1 0 54208 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3578_
timestamp 1698431365
transform -1 0 51632 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3579_
timestamp 1698431365
transform 1 0 43680 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3580_
timestamp 1698431365
transform 1 0 42224 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3581_
timestamp 1698431365
transform 1 0 42224 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3582_
timestamp 1698431365
transform -1 0 48160 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3583_
timestamp 1698431365
transform -1 0 43232 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3584_
timestamp 1698431365
transform 1 0 32704 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3585_
timestamp 1698431365
transform 1 0 29904 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3586_
timestamp 1698431365
transform -1 0 32480 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3587_
timestamp 1698431365
transform 1 0 26768 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3588_
timestamp 1698431365
transform -1 0 33152 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3589_
timestamp 1698431365
transform -1 0 29904 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3590_
timestamp 1698431365
transform 1 0 29232 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3591_
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3592_
timestamp 1698431365
transform 1 0 30800 0 1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3593_
timestamp 1698431365
transform 1 0 30912 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3594_
timestamp 1698431365
transform -1 0 31584 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3595_
timestamp 1698431365
transform 1 0 37408 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3596_
timestamp 1698431365
transform -1 0 35616 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3597_
timestamp 1698431365
transform -1 0 40544 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3598_
timestamp 1698431365
transform 1 0 36288 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3599_
timestamp 1698431365
transform -1 0 9184 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3600_
timestamp 1698431365
transform -1 0 14560 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3601_
timestamp 1698431365
transform -1 0 13440 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3602_
timestamp 1698431365
transform 1 0 10976 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3603_
timestamp 1698431365
transform -1 0 12320 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3604_
timestamp 1698431365
transform -1 0 2800 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3605_
timestamp 1698431365
transform -1 0 3248 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3606_
timestamp 1698431365
transform -1 0 9184 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3607_
timestamp 1698431365
transform 1 0 4928 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3608_
timestamp 1698431365
transform 1 0 2240 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3609_
timestamp 1698431365
transform -1 0 5264 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3610_
timestamp 1698431365
transform 1 0 2128 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3611_
timestamp 1698431365
transform -1 0 14672 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3612_
timestamp 1698431365
transform 1 0 18032 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3613_
timestamp 1698431365
transform 1 0 14784 0 -1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3614_
timestamp 1698431365
transform -1 0 19824 0 -1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3615_
timestamp 1698431365
transform 1 0 14224 0 -1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3616_
timestamp 1698431365
transform 1 0 27888 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3617_
timestamp 1698431365
transform -1 0 22400 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3618_
timestamp 1698431365
transform -1 0 26768 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3619_
timestamp 1698431365
transform -1 0 28784 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3620_
timestamp 1698431365
transform -1 0 28336 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3621_
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3622_
timestamp 1698431365
transform 1 0 13664 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3623_
timestamp 1698431365
transform -1 0 17472 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3624_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3625_
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3626_
timestamp 1698431365
transform -1 0 2800 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3627_
timestamp 1698431365
transform 1 0 5600 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3628_
timestamp 1698431365
transform 1 0 7504 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3629_
timestamp 1698431365
transform -1 0 10080 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3630_
timestamp 1698431365
transform -1 0 8176 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3631_
timestamp 1698431365
transform -1 0 9184 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3632_
timestamp 1698431365
transform 1 0 20608 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3633_
timestamp 1698431365
transform 1 0 15680 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3634_
timestamp 1698431365
transform 1 0 16576 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3635_
timestamp 1698431365
transform 1 0 23184 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3636_
timestamp 1698431365
transform -1 0 18928 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3637_
timestamp 1698431365
transform 1 0 23968 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3638_
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3639_
timestamp 1698431365
transform -1 0 15344 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3640_
timestamp 1698431365
transform 1 0 21728 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _3641_
timestamp 1698431365
transform -1 0 24080 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3642_
timestamp 1698431365
transform -1 0 7056 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3643_
timestamp 1698431365
transform 1 0 13440 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3644_
timestamp 1698431365
transform 1 0 14336 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3645_
timestamp 1698431365
transform 1 0 13664 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3646_
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3647_
timestamp 1698431365
transform -1 0 5936 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3648_
timestamp 1698431365
transform 1 0 4144 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3649_
timestamp 1698431365
transform -1 0 9968 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3650_
timestamp 1698431365
transform 1 0 7392 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3651_
timestamp 1698431365
transform 1 0 7616 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3652_
timestamp 1698431365
transform 1 0 8176 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3653_
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3654_
timestamp 1698431365
transform -1 0 38864 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3655_
timestamp 1698431365
transform 1 0 22960 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3656_
timestamp 1698431365
transform 1 0 17808 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3657_
timestamp 1698431365
transform -1 0 15008 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3658_
timestamp 1698431365
transform -1 0 18368 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3659_
timestamp 1698431365
transform -1 0 49952 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3660_
timestamp 1698431365
transform 1 0 29680 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3661_
timestamp 1698431365
transform 1 0 30800 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3662_
timestamp 1698431365
transform 1 0 31024 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3663_
timestamp 1698431365
transform -1 0 32368 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3664_
timestamp 1698431365
transform -1 0 47824 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3665_
timestamp 1698431365
transform -1 0 19264 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3666_
timestamp 1698431365
transform 1 0 19264 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3667_
timestamp 1698431365
transform 1 0 18592 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3668_
timestamp 1698431365
transform -1 0 22288 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3669_
timestamp 1698431365
transform 1 0 9408 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3670_
timestamp 1698431365
transform 1 0 8400 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3671_
timestamp 1698431365
transform 1 0 14560 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3672_
timestamp 1698431365
transform -1 0 7504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3673_
timestamp 1698431365
transform 1 0 7504 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3674_
timestamp 1698431365
transform 1 0 8064 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3675_
timestamp 1698431365
transform -1 0 47936 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3676_
timestamp 1698431365
transform 1 0 40880 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3677_
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3678_
timestamp 1698431365
transform 1 0 46144 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3679_
timestamp 1698431365
transform -1 0 44128 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3680_
timestamp 1698431365
transform 1 0 51408 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3681_
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3682_
timestamp 1698431365
transform 1 0 43792 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3683_
timestamp 1698431365
transform 1 0 35392 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3684_
timestamp 1698431365
transform -1 0 43232 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3685_
timestamp 1698431365
transform -1 0 39312 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3686_
timestamp 1698431365
transform -1 0 45584 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3687_
timestamp 1698431365
transform -1 0 44800 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3688_
timestamp 1698431365
transform -1 0 42224 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3689_
timestamp 1698431365
transform -1 0 43904 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3690_
timestamp 1698431365
transform 1 0 28448 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3691_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3692_
timestamp 1698431365
transform 1 0 32144 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3693_
timestamp 1698431365
transform -1 0 33936 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3694_
timestamp 1698431365
transform -1 0 28784 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3695_
timestamp 1698431365
transform -1 0 31584 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3696_
timestamp 1698431365
transform -1 0 26768 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3697_
timestamp 1698431365
transform -1 0 40432 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3698_
timestamp 1698431365
transform 1 0 47488 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3699_
timestamp 1698431365
transform -1 0 48384 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3700_
timestamp 1698431365
transform -1 0 55888 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3701_
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3702_
timestamp 1698431365
transform 1 0 47264 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3703_
timestamp 1698431365
transform -1 0 54544 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3704_
timestamp 1698431365
transform -1 0 55328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3705_
timestamp 1698431365
transform -1 0 54992 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3706_
timestamp 1698431365
transform 1 0 61264 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3707_
timestamp 1698431365
transform 1 0 60368 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3708_
timestamp 1698431365
transform 1 0 56224 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3709_
timestamp 1698431365
transform -1 0 49504 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3710_
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3711_
timestamp 1698431365
transform 1 0 49840 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3712_
timestamp 1698431365
transform 1 0 47712 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3713_
timestamp 1698431365
transform 1 0 51184 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3714_
timestamp 1698431365
transform 1 0 50176 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3715_
timestamp 1698431365
transform 1 0 35056 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3716_
timestamp 1698431365
transform -1 0 37072 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3717_
timestamp 1698431365
transform -1 0 33824 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3718_
timestamp 1698431365
transform 1 0 33712 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3719_
timestamp 1698431365
transform 1 0 33712 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3720_
timestamp 1698431365
transform -1 0 33712 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3721_
timestamp 1698431365
transform 1 0 58240 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3722_
timestamp 1698431365
transform 1 0 59248 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3723_
timestamp 1698431365
transform 1 0 61488 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3724_
timestamp 1698431365
transform -1 0 58240 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3725_
timestamp 1698431365
transform -1 0 62384 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3726_
timestamp 1698431365
transform 1 0 60368 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3727_
timestamp 1698431365
transform -1 0 53200 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3728_
timestamp 1698431365
transform 1 0 61264 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3729_
timestamp 1698431365
transform -1 0 53424 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3730_
timestamp 1698431365
transform 1 0 53424 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3731_
timestamp 1698431365
transform 1 0 53760 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3732_
timestamp 1698431365
transform 1 0 54096 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3733_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3734_
timestamp 1698431365
transform 1 0 46144 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3735_
timestamp 1698431365
transform 1 0 42448 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3736_
timestamp 1698431365
transform 1 0 41664 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3737_
timestamp 1698431365
transform -1 0 44352 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3738_
timestamp 1698431365
transform 1 0 41328 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3739_
timestamp 1698431365
transform -1 0 40096 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3740_
timestamp 1698431365
transform -1 0 41328 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3741_
timestamp 1698431365
transform -1 0 38080 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3742_
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3743_
timestamp 1698431365
transform 1 0 30688 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3744_
timestamp 1698431365
transform -1 0 32704 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3745_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 49280 0 1 56448
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3746_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41216 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3747_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43904 0 -1 58016
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3748_
timestamp 1698431365
transform 1 0 46816 0 1 56448
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3749_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45920 0 1 53312
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3750_
timestamp 1698431365
transform 1 0 42448 0 -1 56448
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3751_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3752_
timestamp 1698431365
transform 1 0 56896 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3753_
timestamp 1698431365
transform 1 0 53088 0 1 56448
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3754_
timestamp 1698431365
transform -1 0 60256 0 -1 54880
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3755_
timestamp 1698431365
transform 1 0 52080 0 -1 50176
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3756_
timestamp 1698431365
transform 1 0 49056 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3757_
timestamp 1698431365
transform -1 0 57680 0 1 50176
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3758_
timestamp 1698431365
transform -1 0 57680 0 1 48608
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3759_
timestamp 1698431365
transform 1 0 50960 0 -1 47040
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3760_
timestamp 1698431365
transform 1 0 51968 0 -1 48608
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3761_
timestamp 1698431365
transform 1 0 45024 0 -1 51744
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3762_
timestamp 1698431365
transform 1 0 40096 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3763_
timestamp 1698431365
transform 1 0 41888 0 -1 53312
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3764_
timestamp 1698431365
transform 1 0 41216 0 -1 51744
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3765_
timestamp 1698431365
transform 1 0 44912 0 -1 45472
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3766_
timestamp 1698431365
transform 1 0 41216 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3767_
timestamp 1698431365
transform 1 0 43456 0 -1 40768
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3768_
timestamp 1698431365
transform -1 0 47152 0 1 39200
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3769_
timestamp 1698431365
transform 1 0 44800 0 -1 43904
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3770_
timestamp 1698431365
transform 1 0 42000 0 1 40768
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3771_
timestamp 1698431365
transform 1 0 38304 0 1 47040
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3772_
timestamp 1698431365
transform 1 0 34048 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3773_
timestamp 1698431365
transform -1 0 39088 0 1 45472
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3774_
timestamp 1698431365
transform 1 0 37408 0 -1 47040
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3775_
timestamp 1698431365
transform 1 0 31584 0 1 45472
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3776_
timestamp 1698431365
transform 1 0 29120 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3777_
timestamp 1698431365
transform -1 0 37632 0 -1 42336
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3778_
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3779_
timestamp 1698431365
transform 1 0 30464 0 1 43904
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3780_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3781_
timestamp 1698431365
transform 1 0 26320 0 1 40768
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3782_
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3783_
timestamp 1698431365
transform -1 0 28112 0 -1 39200
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3784_
timestamp 1698431365
transform 1 0 28336 0 -1 36064
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3785_
timestamp 1698431365
transform -1 0 27216 0 1 59584
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3786_
timestamp 1698431365
transform -1 0 28336 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3787_
timestamp 1698431365
transform 1 0 21280 0 1 59584
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3788_
timestamp 1698431365
transform -1 0 22960 0 -1 59584
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3789_
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3790_
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3791_
timestamp 1698431365
transform -1 0 36064 0 1 58016
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3792_
timestamp 1698431365
transform 1 0 34272 0 1 56448
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3793_
timestamp 1698431365
transform 1 0 32928 0 1 54880
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3794_
timestamp 1698431365
transform 1 0 30240 0 -1 59584
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3795_
timestamp 1698431365
transform 1 0 27328 0 -1 53312
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3796_
timestamp 1698431365
transform 1 0 25200 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3797_
timestamp 1698431365
transform 1 0 26992 0 -1 51744
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3798_
timestamp 1698431365
transform 1 0 26320 0 -1 50176
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3799_
timestamp 1698431365
transform 1 0 33488 0 1 53312
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3800_
timestamp 1698431365
transform 1 0 34944 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3801_
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3802_
timestamp 1698431365
transform 1 0 37632 0 1 51744
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3803_
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3804_
timestamp 1698431365
transform 1 0 36176 0 -1 50176
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3805_
timestamp 1698431365
transform 1 0 19264 0 -1 51744
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3806_
timestamp 1698431365
transform 1 0 13776 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3807_
timestamp 1698431365
transform 1 0 17584 0 -1 50176
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3808_
timestamp 1698431365
transform -1 0 19600 0 1 50176
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3809_
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3810_
timestamp 1698431365
transform 1 0 7056 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3811_
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3812_
timestamp 1698431365
transform -1 0 12432 0 1 51744
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3813_
timestamp 1698431365
transform 1 0 10080 0 -1 48608
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3814_
timestamp 1698431365
transform 1 0 10640 0 1 50176
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3815_
timestamp 1698431365
transform 1 0 5824 0 1 47040
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3816_
timestamp 1698431365
transform 1 0 2016 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3817_
timestamp 1698431365
transform 1 0 4368 0 -1 42336
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3818_
timestamp 1698431365
transform 1 0 4368 0 -1 40768
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3819_
timestamp 1698431365
transform 1 0 2240 0 -1 48608
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3820_
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3821_
timestamp 1698431365
transform -1 0 3808 0 1 45472
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3822_
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3823_
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3824_
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3825_
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3826_
timestamp 1698431365
transform -1 0 14672 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3827_
timestamp 1698431365
transform 1 0 14224 0 -1 59584
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3828_
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3829_
timestamp 1698431365
transform 1 0 16016 0 1 54880
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3830_
timestamp 1698431365
transform 1 0 14224 0 1 58016
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3831_
timestamp 1698431365
transform 1 0 18480 0 1 54880
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3832_
timestamp 1698431365
transform -1 0 20720 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3833_
timestamp 1698431365
transform 1 0 18032 0 -1 53312
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3834_
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3835_
timestamp 1698431365
transform 1 0 21392 0 -1 48608
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3836_
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3837_
timestamp 1698431365
transform -1 0 27440 0 1 48608
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3838_
timestamp 1698431365
transform -1 0 28112 0 -1 48608
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3839_
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3840_
timestamp 1698431365
transform -1 0 28784 0 -1 45472
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3841_
timestamp 1698431365
transform 1 0 20944 0 -1 43904
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3842_
timestamp 1698431365
transform 1 0 17696 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3843_
timestamp 1698431365
transform -1 0 22400 0 -1 39200
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3844_
timestamp 1698431365
transform 1 0 20944 0 -1 37632
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3845_
timestamp 1698431365
transform -1 0 19264 0 1 37632
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3846_
timestamp 1698431365
transform 1 0 13664 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3847_
timestamp 1698431365
transform 1 0 18368 0 1 42336
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3848_
timestamp 1698431365
transform 1 0 16016 0 1 45472
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3849_
timestamp 1698431365
transform 1 0 15680 0 1 42336
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3850_
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3851_
timestamp 1698431365
transform 1 0 10080 0 1 40768
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3852_
timestamp 1698431365
transform -1 0 17024 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3853_
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3854_
timestamp 1698431365
transform 1 0 10080 0 -1 42336
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3855_
timestamp 1698431365
transform -1 0 11648 0 -1 34496
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3856_
timestamp 1698431365
transform 1 0 6048 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3857_
timestamp 1698431365
transform -1 0 8736 0 1 36064
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3858_
timestamp 1698431365
transform -1 0 8512 0 -1 28224
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3859_
timestamp 1698431365
transform -1 0 10080 0 1 32928
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3860_
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3861_
timestamp 1698431365
transform 1 0 4816 0 -1 29792
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3862_
timestamp 1698431365
transform -1 0 4816 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3863_
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3864_
timestamp 1698431365
transform -1 0 5152 0 1 28224
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3865_
timestamp 1698431365
transform 1 0 10416 0 -1 32928
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3866_
timestamp 1698431365
transform 1 0 7616 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3867_
timestamp 1698431365
transform 1 0 9744 0 -1 31360
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3868_
timestamp 1698431365
transform 1 0 10080 0 -1 29792
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3869_
timestamp 1698431365
transform 1 0 18032 0 -1 31360
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3870_
timestamp 1698431365
transform 1 0 24976 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3871_
timestamp 1698431365
transform 1 0 19152 0 -1 34496
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3872_
timestamp 1698431365
transform 1 0 26320 0 1 32928
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3873_
timestamp 1698431365
transform 1 0 22624 0 1 32928
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3874_
timestamp 1698431365
transform 1 0 17696 0 1 34496
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3875_
timestamp 1698431365
transform -1 0 26992 0 1 28224
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3876_
timestamp 1698431365
transform 1 0 21504 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3877_
timestamp 1698431365
transform 1 0 26544 0 1 29792
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3878_
timestamp 1698431365
transform 1 0 27888 0 -1 28224
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3879_
timestamp 1698431365
transform 1 0 10640 0 1 28224
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3880_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3881_
timestamp 1698431365
transform 1 0 9744 0 -1 28224
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3882_
timestamp 1698431365
transform 1 0 20272 0 -1 36064
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3883_
timestamp 1698431365
transform 1 0 14112 0 1 25088
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3884_
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3885_
timestamp 1698431365
transform 1 0 10752 0 -1 23520
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3886_
timestamp 1698431365
transform 1 0 21168 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3887_
timestamp 1698431365
transform -1 0 17808 0 1 17248
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3888_
timestamp 1698431365
transform 1 0 16576 0 1 15680
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3889_
timestamp 1698431365
transform 1 0 9856 0 1 20384
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3890_
timestamp 1698431365
transform 1 0 11424 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3891_
timestamp 1698431365
transform 1 0 10192 0 -1 17248
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3892_
timestamp 1698431365
transform -1 0 17024 0 -1 14112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3893_
timestamp 1698431365
transform 1 0 14224 0 -1 15680
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3894_
timestamp 1698431365
transform 1 0 10752 0 -1 18816
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3895_
timestamp 1698431365
transform 1 0 2128 0 1 18816
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3896_
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3897_
timestamp 1698431365
transform 1 0 3024 0 1 17248
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3898_
timestamp 1698431365
transform 1 0 4144 0 -1 18816
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3899_
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3900_
timestamp 1698431365
transform 1 0 6608 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3901_
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3902_
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3903_
timestamp 1698431365
transform -1 0 4032 0 1 21952
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3904_
timestamp 1698431365
transform 1 0 2352 0 -1 26656
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3905_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3906_
timestamp 1698431365
transform 1 0 17472 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3907_
timestamp 1698431365
transform -1 0 22064 0 -1 26656
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3908_
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3909_
timestamp 1698431365
transform -1 0 17808 0 1 23520
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3910_
timestamp 1698431365
transform 1 0 17360 0 -1 26656
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3911_
timestamp 1698431365
transform 1 0 22624 0 1 21952
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3912_
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3913_
timestamp 1698431365
transform -1 0 27328 0 -1 21952
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3914_
timestamp 1698431365
transform 1 0 22624 0 -1 26656
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3915_
timestamp 1698431365
transform 1 0 27328 0 -1 21952
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3916_
timestamp 1698431365
transform 1 0 32144 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3917_
timestamp 1698431365
transform 1 0 33488 0 -1 23520
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3918_
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3919_
timestamp 1698431365
transform -1 0 32368 0 -1 23520
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3920_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3921_
timestamp 1698431365
transform 1 0 30352 0 1 18816
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3922_
timestamp 1698431365
transform 1 0 21840 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3923_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3924_
timestamp 1698431365
transform 1 0 31696 0 1 17248
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3925_
timestamp 1698431365
transform -1 0 26096 0 1 15680
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3926_
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3927_
timestamp 1698431365
transform 1 0 18704 0 1 14112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3928_
timestamp 1698431365
transform -1 0 20944 0 -1 15680
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3929_
timestamp 1698431365
transform -1 0 25088 0 1 14112
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3930_
timestamp 1698431365
transform 1 0 19152 0 -1 14112
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3931_
timestamp 1698431365
transform -1 0 19712 0 -1 6272
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3932_
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3933_
timestamp 1698431365
transform 1 0 17696 0 1 6272
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3934_
timestamp 1698431365
transform -1 0 19488 0 -1 7840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3935_
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3936_
timestamp 1698431365
transform 1 0 12544 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3937_
timestamp 1698431365
transform 1 0 10080 0 -1 7840
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3938_
timestamp 1698431365
transform -1 0 12656 0 -1 9408
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3939_
timestamp 1698431365
transform -1 0 15792 0 1 10976
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3940_
timestamp 1698431365
transform 1 0 8624 0 1 7840
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3941_
timestamp 1698431365
transform 1 0 2800 0 1 10976
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3942_
timestamp 1698431365
transform -1 0 12992 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3943_
timestamp 1698431365
transform 1 0 3024 0 1 12544
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3944_
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3945_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3946_
timestamp 1698431365
transform 1 0 34832 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3947_
timestamp 1698431365
transform 1 0 35504 0 -1 26656
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3948_
timestamp 1698431365
transform 1 0 35616 0 -1 25088
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3949_
timestamp 1698431365
transform 1 0 42000 0 1 21952
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3950_
timestamp 1698431365
transform -1 0 49728 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3951_
timestamp 1698431365
transform -1 0 49616 0 1 26656
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3952_
timestamp 1698431365
transform 1 0 41216 0 -1 25088
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3953_
timestamp 1698431365
transform -1 0 45248 0 -1 26656
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3954_
timestamp 1698431365
transform 1 0 42000 0 1 23520
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3955_
timestamp 1698431365
transform -1 0 51744 0 1 20384
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3956_
timestamp 1698431365
transform 1 0 47488 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3957_
timestamp 1698431365
transform 1 0 49728 0 -1 20384
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3958_
timestamp 1698431365
transform 1 0 50624 0 -1 21952
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3959_
timestamp 1698431365
transform 1 0 43344 0 -1 20384
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3960_
timestamp 1698431365
transform 1 0 37296 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3961_
timestamp 1698431365
transform 1 0 41104 0 -1 20384
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3962_
timestamp 1698431365
transform -1 0 39312 0 1 18816
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3963_
timestamp 1698431365
transform -1 0 47712 0 1 17248
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3964_
timestamp 1698431365
transform 1 0 39648 0 1 18816
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3965_
timestamp 1698431365
transform 1 0 42896 0 -1 10976
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3966_
timestamp 1698431365
transform 1 0 46592 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3967_
timestamp 1698431365
transform -1 0 50848 0 -1 7840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3968_
timestamp 1698431365
transform 1 0 49504 0 1 7840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3969_
timestamp 1698431365
transform -1 0 42784 0 1 4704
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3970_
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3971_
timestamp 1698431365
transform -1 0 46480 0 -1 4704
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3972_
timestamp 1698431365
transform -1 0 43008 0 -1 4704
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3973_
timestamp 1698431365
transform -1 0 42448 0 1 6272
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3974_
timestamp 1698431365
transform 1 0 42672 0 -1 6272
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3975_
timestamp 1698431365
transform -1 0 39984 0 1 6272
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3976_
timestamp 1698431365
transform -1 0 40096 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3977_
timestamp 1698431365
transform -1 0 38080 0 1 3136
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _3978_
timestamp 1698431365
transform -1 0 36736 0 -1 4704
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3979_
timestamp 1698431365
transform 1 0 29456 0 -1 4704
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3980_
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3981_
timestamp 1698431365
transform 1 0 25536 0 -1 6272
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3982_
timestamp 1698431365
transform -1 0 26992 0 1 7840
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3983_
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3984_
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3985_
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3986_
timestamp 1698431365
transform 1 0 50736 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3987_
timestamp 1698431365
transform -1 0 51072 0 -1 28224
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3988_
timestamp 1698431365
transform 1 0 45248 0 1 29792
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3989_
timestamp 1698431365
transform 1 0 49616 0 -1 29792
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3990_
timestamp 1698431365
transform 1 0 47488 0 1 28224
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3991_
timestamp 1698431365
transform -1 0 62384 0 -1 28224
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3992_
timestamp 1698431365
transform 1 0 59136 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3993_
timestamp 1698431365
transform 1 0 57904 0 1 29792
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3994_
timestamp 1698431365
transform -1 0 60144 0 1 28224
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3995_
timestamp 1698431365
transform 1 0 60144 0 -1 23520
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3996_
timestamp 1698431365
transform 1 0 58016 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _3997_
timestamp 1698431365
transform -1 0 62384 0 -1 21952
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _3998_
timestamp 1698431365
transform -1 0 60144 0 1 21952
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _3999_
timestamp 1698431365
transform 1 0 54656 0 1 21952
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4000_
timestamp 1698431365
transform 1 0 57680 0 1 23520
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4001_
timestamp 1698431365
transform -1 0 60144 0 1 17248
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4002_
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4003_
timestamp 1698431365
transform -1 0 60144 0 -1 17248
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4004_
timestamp 1698431365
transform -1 0 60704 0 -1 18816
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4005_
timestamp 1698431365
transform -1 0 54320 0 -1 15680
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4006_
timestamp 1698431365
transform 1 0 49952 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4007_
timestamp 1698431365
transform 1 0 53424 0 1 10976
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4008_
timestamp 1698431365
transform -1 0 54768 0 1 9408
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4009_
timestamp 1698431365
transform 1 0 49280 0 1 14112
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4010_
timestamp 1698431365
transform 1 0 52864 0 -1 12544
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4011_
timestamp 1698431365
transform 1 0 45920 0 -1 15680
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4012_
timestamp 1698431365
transform 1 0 38416 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4013_
timestamp 1698431365
transform -1 0 46928 0 1 14112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4014_
timestamp 1698431365
transform -1 0 47600 0 -1 14112
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4015_
timestamp 1698431365
transform -1 0 39648 0 -1 15680
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4016_
timestamp 1698431365
transform 1 0 33376 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4017_
timestamp 1698431365
transform -1 0 40320 0 1 10976
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4018_
timestamp 1698431365
transform -1 0 38752 0 -1 10976
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4019_
timestamp 1698431365
transform 1 0 34944 0 -1 15680
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4020_
timestamp 1698431365
transform 1 0 33488 0 -1 12544
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4021_
timestamp 1698431365
transform 1 0 29904 0 -1 15680
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4022_
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4023_
timestamp 1698431365
transform 1 0 26320 0 -1 12544
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4024_
timestamp 1698431365
transform -1 0 28560 0 1 12544
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4025_
timestamp 1698431365
transform 1 0 51296 0 -1 42336
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4026_
timestamp 1698431365
transform -1 0 53424 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4027_
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _4028_
timestamp 1698431365
transform -1 0 50288 0 1 42336
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4029_
timestamp 1698431365
transform 1 0 57904 0 1 43904
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4030_
timestamp 1698431365
transform 1 0 58576 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4031_
timestamp 1698431365
transform 1 0 57904 0 1 45472
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4032_
timestamp 1698431365
transform 1 0 57008 0 -1 43904
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4033_
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4034_
timestamp 1698431365
transform 1 0 59136 0 -1 48608
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _4035_
timestamp 1698431365
transform 1 0 57008 0 1 40768
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4036_
timestamp 1698431365
transform 1 0 58688 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4037_
timestamp 1698431365
transform 1 0 53984 0 -1 39200
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _4038_
timestamp 1698431365
transform -1 0 60144 0 1 36064
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4039_
timestamp 1698431365
transform -1 0 61600 0 -1 34496
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4040_
timestamp 1698431365
transform 1 0 51072 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4041_
timestamp 1698431365
transform -1 0 60144 0 1 32928
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4042_
timestamp 1698431365
transform -1 0 59696 0 1 31360
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4043_
timestamp 1698431365
transform 1 0 54768 0 1 31360
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4044_
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _4045_
timestamp 1698431365
transform 1 0 48608 0 1 31360
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4046_
timestamp 1698431365
transform 1 0 45136 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4047_
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _4048_
timestamp 1698431365
transform 1 0 48048 0 1 32928
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4049_
timestamp 1698431365
transform -1 0 46144 0 -1 34496
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4050_
timestamp 1698431365
transform 1 0 42000 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4051_
timestamp 1698431365
transform 1 0 42896 0 -1 31360
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  _4052_
timestamp 1698431365
transform 1 0 41440 0 1 31360
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4053_
timestamp 1698431365
transform -1 0 44464 0 1 36064
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4054_
timestamp 1698431365
transform 1 0 41776 0 1 32928
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _4055_
timestamp 1698431365
transform 1 0 39200 0 1 37632
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4056_
timestamp 1698431365
transform 1 0 36960 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4057_
timestamp 1698431365
transform 1 0 37856 0 -1 39200
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  _4058_
timestamp 1698431365
transform -1 0 39984 0 -1 40768
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4059_
timestamp 1698431365
transform -1 0 39536 0 -1 31360
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _4060_
timestamp 1698431365
transform 1 0 34048 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4061_
timestamp 1698431365
transform 1 0 30352 0 1 31360
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _4062_
timestamp 1698431365
transform -1 0 31360 0 -1 32928
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4063_
timestamp 1698431365
transform -1 0 36848 0 -1 32928
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _4064_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__I test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40992 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A1
timestamp 1698431365
transform 1 0 42896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A2
timestamp 1698431365
transform 1 0 36848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__I1
timestamp 1698431365
transform -1 0 49504 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A1
timestamp 1698431365
transform 1 0 61264 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__B
timestamp 1698431365
transform -1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__I1
timestamp 1698431365
transform 1 0 60368 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__A1
timestamp 1698431365
transform 1 0 49168 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A2
timestamp 1698431365
transform -1 0 47712 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__B
timestamp 1698431365
transform 1 0 60704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__A2
timestamp 1698431365
transform -1 0 60144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__I1
timestamp 1698431365
transform -1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1863__I1
timestamp 1698431365
transform -1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__A2
timestamp 1698431365
transform 1 0 14000 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__A2
timestamp 1698431365
transform 1 0 37072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__A2
timestamp 1698431365
transform 1 0 14000 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A1
timestamp 1698431365
transform -1 0 36176 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__A1
timestamp 1698431365
transform 1 0 41104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__A2
timestamp 1698431365
transform -1 0 40880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__I
timestamp 1698431365
transform 1 0 29680 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__I0
timestamp 1698431365
transform -1 0 22736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__A1
timestamp 1698431365
transform 1 0 29232 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__A2
timestamp 1698431365
transform -1 0 27888 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__I
timestamp 1698431365
transform 1 0 61824 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A1
timestamp 1698431365
transform -1 0 60816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A2
timestamp 1698431365
transform -1 0 61152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1698431365
transform 1 0 61936 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__I1
timestamp 1698431365
transform 1 0 57792 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__C
timestamp 1698431365
transform -1 0 42336 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1936__A1
timestamp 1698431365
transform 1 0 59248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__A2
timestamp 1698431365
transform -1 0 46144 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__A2
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__I
timestamp 1698431365
transform 1 0 38304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__A2
timestamp 1698431365
transform -1 0 45696 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A1
timestamp 1698431365
transform -1 0 45248 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A2
timestamp 1698431365
transform 1 0 43680 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__A1
timestamp 1698431365
transform -1 0 46592 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__A1
timestamp 1698431365
transform -1 0 56896 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__A2
timestamp 1698431365
transform 1 0 48048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1961__S
timestamp 1698431365
transform -1 0 54544 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__A1
timestamp 1698431365
transform 1 0 61264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A1
timestamp 1698431365
transform 1 0 61488 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A2
timestamp 1698431365
transform -1 0 61376 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__I1
timestamp 1698431365
transform 1 0 36288 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A2
timestamp 1698431365
transform 1 0 38864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__A1
timestamp 1698431365
transform 1 0 44240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__A1
timestamp 1698431365
transform -1 0 48160 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__A2
timestamp 1698431365
transform -1 0 49056 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__B
timestamp 1698431365
transform 1 0 47488 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__I0
timestamp 1698431365
transform 1 0 44912 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A2
timestamp 1698431365
transform -1 0 47152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2067__I
timestamp 1698431365
transform 1 0 30128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2070__A2
timestamp 1698431365
transform -1 0 51408 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A1
timestamp 1698431365
transform 1 0 50176 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__A2
timestamp 1698431365
transform 1 0 44016 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__S
timestamp 1698431365
transform -1 0 42000 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__I1
timestamp 1698431365
transform -1 0 61264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2107__A2
timestamp 1698431365
transform 1 0 60256 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2112__A1
timestamp 1698431365
transform 1 0 62160 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2112__A2
timestamp 1698431365
transform -1 0 51296 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__I1
timestamp 1698431365
transform 1 0 6720 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__I
timestamp 1698431365
transform -1 0 6496 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__I1
timestamp 1698431365
transform -1 0 13552 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A2
timestamp 1698431365
transform -1 0 8512 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__A2
timestamp 1698431365
transform 1 0 9856 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2141__A1
timestamp 1698431365
transform 1 0 11200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__A1
timestamp 1698431365
transform 1 0 42336 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__A2
timestamp 1698431365
transform 1 0 44240 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__B
timestamp 1698431365
transform 1 0 46368 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__A1
timestamp 1698431365
transform 1 0 54992 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__A2
timestamp 1698431365
transform 1 0 54992 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2160__I1
timestamp 1698431365
transform -1 0 41216 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__C
timestamp 1698431365
transform -1 0 7616 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2171__A1
timestamp 1698431365
transform -1 0 40768 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2171__B
timestamp 1698431365
transform 1 0 35616 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__A2
timestamp 1698431365
transform 1 0 46704 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__A1
timestamp 1698431365
transform 1 0 42224 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__A1
timestamp 1698431365
transform 1 0 37184 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__B
timestamp 1698431365
transform -1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__S
timestamp 1698431365
transform 1 0 36288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__I1
timestamp 1698431365
transform -1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2212__A2
timestamp 1698431365
transform 1 0 40432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2217__A2
timestamp 1698431365
transform -1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2228__I1
timestamp 1698431365
transform 1 0 7616 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2239__A2
timestamp 1698431365
transform -1 0 7952 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2245__A1
timestamp 1698431365
transform -1 0 6272 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__A1
timestamp 1698431365
transform 1 0 24640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__A2
timestamp 1698431365
transform 1 0 12880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__B
timestamp 1698431365
transform -1 0 20048 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__A2
timestamp 1698431365
transform 1 0 8064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__A1
timestamp 1698431365
transform 1 0 30352 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__I
timestamp 1698431365
transform 1 0 25312 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A2
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2267__A1
timestamp 1698431365
transform -1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2268__A1
timestamp 1698431365
transform 1 0 18592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2268__A2
timestamp 1698431365
transform -1 0 27664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__I
timestamp 1698431365
transform -1 0 11536 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__A2
timestamp 1698431365
transform 1 0 13104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2272__A1
timestamp 1698431365
transform -1 0 12656 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2272__A2
timestamp 1698431365
transform 1 0 13552 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2276__A2
timestamp 1698431365
transform 1 0 37744 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2279__A2
timestamp 1698431365
transform -1 0 13664 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__A2
timestamp 1698431365
transform -1 0 34720 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A1
timestamp 1698431365
transform -1 0 7840 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A2
timestamp 1698431365
transform -1 0 7392 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2313__A2
timestamp 1698431365
transform 1 0 38864 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A1
timestamp 1698431365
transform 1 0 37296 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A2
timestamp 1698431365
transform -1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2332__I
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2334__A2
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2336__B
timestamp 1698431365
transform -1 0 36512 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2337__A2
timestamp 1698431365
transform 1 0 35504 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__A1
timestamp 1698431365
transform 1 0 36400 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__A2
timestamp 1698431365
transform -1 0 36176 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2341__A1
timestamp 1698431365
transform -1 0 11536 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2341__A2
timestamp 1698431365
transform -1 0 17248 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__A1
timestamp 1698431365
transform 1 0 42224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__A2
timestamp 1698431365
transform -1 0 43568 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2356__A1
timestamp 1698431365
transform -1 0 2128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2356__A2
timestamp 1698431365
transform -1 0 2016 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2359__I1
timestamp 1698431365
transform 1 0 25312 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2372__A2
timestamp 1698431365
transform 1 0 13664 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2373__A2
timestamp 1698431365
transform 1 0 25312 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__A2
timestamp 1698431365
transform -1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2386__B
timestamp 1698431365
transform -1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2387__A1
timestamp 1698431365
transform 1 0 41664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2387__A2
timestamp 1698431365
transform 1 0 40320 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2387__B
timestamp 1698431365
transform 1 0 40208 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__A2
timestamp 1698431365
transform -1 0 6496 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2393__A1
timestamp 1698431365
transform 1 0 39984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2393__B
timestamp 1698431365
transform 1 0 41664 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A2
timestamp 1698431365
transform -1 0 8288 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__A1
timestamp 1698431365
transform -1 0 10640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__A2
timestamp 1698431365
transform -1 0 6720 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2399__A2
timestamp 1698431365
transform 1 0 9632 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2407__A2
timestamp 1698431365
transform 1 0 10976 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2415__A1
timestamp 1698431365
transform 1 0 7504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2415__A2
timestamp 1698431365
transform -1 0 10192 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2415__B
timestamp 1698431365
transform -1 0 10192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2431__A1
timestamp 1698431365
transform -1 0 2688 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2431__A2
timestamp 1698431365
transform -1 0 4592 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2431__B
timestamp 1698431365
transform 1 0 10304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__A2
timestamp 1698431365
transform 1 0 13776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2448__A2
timestamp 1698431365
transform -1 0 12432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2449__B
timestamp 1698431365
transform 1 0 8512 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2450__A2
timestamp 1698431365
transform 1 0 8064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2454__I
timestamp 1698431365
transform -1 0 13776 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2455__A1
timestamp 1698431365
transform 1 0 7168 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2455__A2
timestamp 1698431365
transform -1 0 8400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2456__A1
timestamp 1698431365
transform -1 0 6944 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2457__A2
timestamp 1698431365
transform 1 0 4368 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__A1
timestamp 1698431365
transform 1 0 4480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__A2
timestamp 1698431365
transform 1 0 4928 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__B
timestamp 1698431365
transform -1 0 5600 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__I
timestamp 1698431365
transform -1 0 4928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__A2
timestamp 1698431365
transform 1 0 9968 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2502__A1
timestamp 1698431365
transform 1 0 4144 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A2
timestamp 1698431365
transform -1 0 12208 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2515__I1
timestamp 1698431365
transform -1 0 2352 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__I1
timestamp 1698431365
transform 1 0 3024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__A1
timestamp 1698431365
transform 1 0 3920 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A2
timestamp 1698431365
transform 1 0 5824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__A2
timestamp 1698431365
transform -1 0 2128 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__A1
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A1
timestamp 1698431365
transform -1 0 10304 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A2
timestamp 1698431365
transform -1 0 12656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__B
timestamp 1698431365
transform -1 0 11984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__A2
timestamp 1698431365
transform -1 0 10192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__A2
timestamp 1698431365
transform -1 0 11088 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__A2
timestamp 1698431365
transform 1 0 8624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2556__A2
timestamp 1698431365
transform -1 0 11760 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2557__A1
timestamp 1698431365
transform -1 0 10752 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2563__A2
timestamp 1698431365
transform 1 0 10864 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2566__A2
timestamp 1698431365
transform 1 0 39312 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__I1
timestamp 1698431365
transform 1 0 52080 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__I1
timestamp 1698431365
transform -1 0 13888 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__A1
timestamp 1698431365
transform 1 0 26768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2591__A2
timestamp 1698431365
transform 1 0 31920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__A2
timestamp 1698431365
transform -1 0 29904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__A2
timestamp 1698431365
transform -1 0 10528 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2613__A1
timestamp 1698431365
transform 1 0 8064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__I
timestamp 1698431365
transform -1 0 21056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__A2
timestamp 1698431365
transform -1 0 12208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__A2
timestamp 1698431365
transform -1 0 2128 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2620__A1
timestamp 1698431365
transform -1 0 2240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2622__A2
timestamp 1698431365
transform -1 0 8736 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__I1
timestamp 1698431365
transform -1 0 21616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__A1
timestamp 1698431365
transform 1 0 23408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__A2
timestamp 1698431365
transform 1 0 21952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__A1
timestamp 1698431365
transform -1 0 18928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__A1
timestamp 1698431365
transform -1 0 2352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__A2
timestamp 1698431365
transform -1 0 2016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2667__A2
timestamp 1698431365
transform -1 0 10976 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__A1
timestamp 1698431365
transform 1 0 7840 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__A2
timestamp 1698431365
transform -1 0 9856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__A1
timestamp 1698431365
transform 1 0 5040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__I1
timestamp 1698431365
transform 1 0 3696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__A2
timestamp 1698431365
transform -1 0 3024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__B
timestamp 1698431365
transform -1 0 7504 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__A1
timestamp 1698431365
transform -1 0 8848 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__A2
timestamp 1698431365
transform -1 0 2016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2715__B
timestamp 1698431365
transform -1 0 3696 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2716__A2
timestamp 1698431365
transform -1 0 4368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2719__A1
timestamp 1698431365
transform -1 0 2128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2720__A2
timestamp 1698431365
transform -1 0 2688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2722__A2
timestamp 1698431365
transform -1 0 11424 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2723__A1
timestamp 1698431365
transform -1 0 2800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2723__A2
timestamp 1698431365
transform -1 0 3696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__A2
timestamp 1698431365
transform -1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__A1
timestamp 1698431365
transform -1 0 4928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__A1
timestamp 1698431365
transform 1 0 29232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__A2
timestamp 1698431365
transform 1 0 28784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__A1
timestamp 1698431365
transform -1 0 31472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__A2
timestamp 1698431365
transform 1 0 43568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__B
timestamp 1698431365
transform -1 0 32816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__A2
timestamp 1698431365
transform 1 0 33376 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2749__I0
timestamp 1698431365
transform 1 0 39760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2761__A1
timestamp 1698431365
transform 1 0 48160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2761__A2
timestamp 1698431365
transform -1 0 23968 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2761__B
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2779__A2
timestamp 1698431365
transform 1 0 14000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2781__B
timestamp 1698431365
transform -1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2782__A2
timestamp 1698431365
transform 1 0 10192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2784__A2
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2786__A2
timestamp 1698431365
transform 1 0 9296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2787__A1
timestamp 1698431365
transform 1 0 8736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2789__A2
timestamp 1698431365
transform -1 0 21728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2798__A1
timestamp 1698431365
transform 1 0 57568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2800__A2
timestamp 1698431365
transform 1 0 13552 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2801__I1
timestamp 1698431365
transform -1 0 9856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2815__A2
timestamp 1698431365
transform 1 0 23744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2820__C
timestamp 1698431365
transform -1 0 24416 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2822__A1
timestamp 1698431365
transform -1 0 2800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2822__A2
timestamp 1698431365
transform -1 0 2240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2832__I
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2833__A1
timestamp 1698431365
transform -1 0 3920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2833__A2
timestamp 1698431365
transform -1 0 3248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2835__A2
timestamp 1698431365
transform -1 0 3920 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2836__A1
timestamp 1698431365
transform -1 0 2352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2837__I
timestamp 1698431365
transform -1 0 21504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2840__A1
timestamp 1698431365
transform 1 0 16240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2840__A2
timestamp 1698431365
transform -1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2842__A2
timestamp 1698431365
transform 1 0 17472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2847__A1
timestamp 1698431365
transform -1 0 15008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2847__A2
timestamp 1698431365
transform -1 0 14560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2854__A1
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2854__A2
timestamp 1698431365
transform 1 0 22400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2854__B
timestamp 1698431365
transform -1 0 24752 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__A2
timestamp 1698431365
transform -1 0 15456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2870__A1
timestamp 1698431365
transform -1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2870__A2
timestamp 1698431365
transform -1 0 25984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2870__B
timestamp 1698431365
transform -1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2886__I
timestamp 1698431365
transform 1 0 56224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2888__A2
timestamp 1698431365
transform 1 0 15792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2889__B
timestamp 1698431365
transform 1 0 9968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2890__A2
timestamp 1698431365
transform -1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2894__A2
timestamp 1698431365
transform -1 0 6944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2895__A1
timestamp 1698431365
transform -1 0 3024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2896__A2
timestamp 1698431365
transform -1 0 2576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2900__I
timestamp 1698431365
transform -1 0 2128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2915__I0
timestamp 1698431365
transform -1 0 4928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2924__A2
timestamp 1698431365
transform -1 0 10080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2926__A2
timestamp 1698431365
transform -1 0 2576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2936__A2
timestamp 1698431365
transform -1 0 3472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2937__A1
timestamp 1698431365
transform 1 0 3248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2939__A2
timestamp 1698431365
transform -1 0 4480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2948__I1
timestamp 1698431365
transform -1 0 50624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2960__I1
timestamp 1698431365
transform 1 0 51408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2962__A2
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2965__A2
timestamp 1698431365
transform 1 0 57792 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2968__A2
timestamp 1698431365
transform 1 0 49728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2970__C
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2972__A2
timestamp 1698431365
transform -1 0 3584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2984__A2
timestamp 1698431365
transform 1 0 2800 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2986__A2
timestamp 1698431365
transform -1 0 16016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2987__A2
timestamp 1698431365
transform -1 0 2576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2989__A2
timestamp 1698431365
transform 1 0 24640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2990__A1
timestamp 1698431365
transform -1 0 19488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2996__A1
timestamp 1698431365
transform -1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2996__A2
timestamp 1698431365
transform -1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2999__A2
timestamp 1698431365
transform -1 0 23296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3008__I1
timestamp 1698431365
transform 1 0 58240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3021__A2
timestamp 1698431365
transform -1 0 58016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3026__C
timestamp 1698431365
transform 1 0 51968 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3028__A2
timestamp 1698431365
transform -1 0 31024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3039__A2
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3041__A2
timestamp 1698431365
transform 1 0 28448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3042__A1
timestamp 1698431365
transform 1 0 13552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3044__A2
timestamp 1698431365
transform -1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3047__A2
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3050__A2
timestamp 1698431365
transform 1 0 22400 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3058__I1
timestamp 1698431365
transform 1 0 52864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3072__A2
timestamp 1698431365
transform 1 0 51632 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3077__C
timestamp 1698431365
transform 1 0 51184 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3079__A2
timestamp 1698431365
transform -1 0 24752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3091__A2
timestamp 1698431365
transform -1 0 23072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3093__A2
timestamp 1698431365
transform -1 0 23632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3094__A1
timestamp 1698431365
transform 1 0 24080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3098__A2
timestamp 1698431365
transform -1 0 25312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3108__I1
timestamp 1698431365
transform 1 0 26992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3119__A2
timestamp 1698431365
transform 1 0 45472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3126__A1
timestamp 1698431365
transform 1 0 16912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3126__A2
timestamp 1698431365
transform 1 0 16352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3126__B
timestamp 1698431365
transform 1 0 16800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3139__B
timestamp 1698431365
transform -1 0 13328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3140__A2
timestamp 1698431365
transform 1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3141__A2
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3143__A1
timestamp 1698431365
transform -1 0 6048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3144__A1
timestamp 1698431365
transform -1 0 8400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3144__A2
timestamp 1698431365
transform 1 0 12432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3145__I
timestamp 1698431365
transform 1 0 43568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3147__A2
timestamp 1698431365
transform 1 0 47824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3149__A2
timestamp 1698431365
transform -1 0 57792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3151__A2
timestamp 1698431365
transform 1 0 60816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3152__A1
timestamp 1698431365
transform -1 0 43904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3154__A2
timestamp 1698431365
transform 1 0 44912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3161__A1
timestamp 1698431365
transform 1 0 61488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3161__A2
timestamp 1698431365
transform 1 0 59248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3165__A1
timestamp 1698431365
transform 1 0 61712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3165__A2
timestamp 1698431365
transform -1 0 61488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3166__A1
timestamp 1698431365
transform 1 0 62160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3168__A2
timestamp 1698431365
transform 1 0 49728 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3185__A1
timestamp 1698431365
transform 1 0 62160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3203__A2
timestamp 1698431365
transform 1 0 59920 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3204__B
timestamp 1698431365
transform 1 0 60592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3205__A2
timestamp 1698431365
transform 1 0 59920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3208__A2
timestamp 1698431365
transform 1 0 59808 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3210__A2
timestamp 1698431365
transform 1 0 60368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3211__A1
timestamp 1698431365
transform 1 0 49392 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3221__I1
timestamp 1698431365
transform -1 0 53424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3235__A2
timestamp 1698431365
transform 1 0 54544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3240__C
timestamp 1698431365
transform -1 0 52192 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3254__A2
timestamp 1698431365
transform 1 0 46704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3255__A1
timestamp 1698431365
transform 1 0 56896 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3259__A2
timestamp 1698431365
transform -1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3262__A2
timestamp 1698431365
transform 1 0 49280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3263__A1
timestamp 1698431365
transform 1 0 52080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3267__A1
timestamp 1698431365
transform 1 0 50736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3267__A2
timestamp 1698431365
transform 1 0 54992 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3272__A1
timestamp 1698431365
transform -1 0 45248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3272__A2
timestamp 1698431365
transform -1 0 58912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3274__A2
timestamp 1698431365
transform 1 0 50736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3290__A1
timestamp 1698431365
transform 1 0 53648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3290__A2
timestamp 1698431365
transform 1 0 60592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3307__A2
timestamp 1698431365
transform -1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3309__B
timestamp 1698431365
transform -1 0 51744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3310__A2
timestamp 1698431365
transform -1 0 47376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3313__A2
timestamp 1698431365
transform 1 0 26544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3315__A2
timestamp 1698431365
transform 1 0 47488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3316__A1
timestamp 1698431365
transform 1 0 50288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3317__B
timestamp 1698431365
transform 1 0 3248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3318__A1
timestamp 1698431365
transform -1 0 22848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3318__A2
timestamp 1698431365
transform -1 0 23744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3318__B
timestamp 1698431365
transform -1 0 23296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3331__I0
timestamp 1698431365
transform -1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3340__A2
timestamp 1698431365
transform 1 0 29232 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3352__A1
timestamp 1698431365
transform -1 0 10976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3352__A2
timestamp 1698431365
transform 1 0 9184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3353__A1
timestamp 1698431365
transform -1 0 27552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3371__A2
timestamp 1698431365
transform -1 0 56336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3375__A2
timestamp 1698431365
transform -1 0 56784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3376__B
timestamp 1698431365
transform 1 0 58464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3377__A2
timestamp 1698431365
transform 1 0 61936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3380__I
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3384__A2
timestamp 1698431365
transform 1 0 59584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3385__A1
timestamp 1698431365
transform 1 0 61040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3388__A1
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3388__A2
timestamp 1698431365
transform 1 0 59136 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3403__B
timestamp 1698431365
transform 1 0 59584 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3404__A2
timestamp 1698431365
transform 1 0 61152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3406__A2
timestamp 1698431365
transform 1 0 55888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3408__A2
timestamp 1698431365
transform 1 0 56336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3409__A1
timestamp 1698431365
transform 1 0 57120 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3412__A1
timestamp 1698431365
transform 1 0 52416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3412__A2
timestamp 1698431365
transform -1 0 53872 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3412__B
timestamp 1698431365
transform -1 0 55664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3427__B
timestamp 1698431365
transform 1 0 54096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3428__A2
timestamp 1698431365
transform -1 0 58912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3433__A2
timestamp 1698431365
transform -1 0 59360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3434__A1
timestamp 1698431365
transform -1 0 47712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3437__A1
timestamp 1698431365
transform -1 0 29680 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3437__A2
timestamp 1698431365
transform -1 0 27664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3439__A1
timestamp 1698431365
transform 1 0 37072 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3440__A1
timestamp 1698431365
transform 1 0 51968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3440__A2
timestamp 1698431365
transform -1 0 45248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3440__B
timestamp 1698431365
transform -1 0 39088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3451__A2
timestamp 1698431365
transform -1 0 30016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3452__A1
timestamp 1698431365
transform -1 0 31136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3453__A2
timestamp 1698431365
transform 1 0 25648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3455__A1
timestamp 1698431365
transform -1 0 29008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3456__A1
timestamp 1698431365
transform -1 0 29008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3456__A2
timestamp 1698431365
transform -1 0 27216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3458__A2
timestamp 1698431365
transform 1 0 61936 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3459__A2
timestamp 1698431365
transform -1 0 49952 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3461__A2
timestamp 1698431365
transform 1 0 60816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3462__A1
timestamp 1698431365
transform -1 0 52976 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3464__A1
timestamp 1698431365
transform -1 0 48608 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3468__I
timestamp 1698431365
transform -1 0 61600 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3474__A2
timestamp 1698431365
transform -1 0 60816 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3483__A2
timestamp 1698431365
transform 1 0 61040 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3484__B
timestamp 1698431365
transform 1 0 54208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3485__A2
timestamp 1698431365
transform 1 0 62160 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3490__A2
timestamp 1698431365
transform -1 0 58464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3491__A1
timestamp 1698431365
transform 1 0 60592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3496__A1
timestamp 1698431365
transform 1 0 59920 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3496__A2
timestamp 1698431365
transform 1 0 56672 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3508__B
timestamp 1698431365
transform 1 0 62160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3509__A2
timestamp 1698431365
transform 1 0 61264 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3512__A2
timestamp 1698431365
transform 1 0 62048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3514__A2
timestamp 1698431365
transform 1 0 56672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3515__A1
timestamp 1698431365
transform 1 0 48832 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3522__A2
timestamp 1698431365
transform 1 0 51072 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3531__A2
timestamp 1698431365
transform 1 0 49504 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3532__B
timestamp 1698431365
transform -1 0 41216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3533__A2
timestamp 1698431365
transform 1 0 43008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3536__A1
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3536__A2
timestamp 1698431365
transform 1 0 43568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3538__A2
timestamp 1698431365
transform 1 0 45808 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3539__A1
timestamp 1698431365
transform 1 0 41888 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3544__A1
timestamp 1698431365
transform 1 0 38752 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3544__A2
timestamp 1698431365
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3546__A2
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3549__A2
timestamp 1698431365
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3552__A2
timestamp 1698431365
transform -1 0 30352 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3553__B
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3554__I
timestamp 1698431365
transform 1 0 34160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3555__A2
timestamp 1698431365
transform -1 0 42560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3555__A3
timestamp 1698431365
transform -1 0 34944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3557__I
timestamp 1698431365
transform -1 0 45136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3558__A2
timestamp 1698431365
transform -1 0 48272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3559__A2
timestamp 1698431365
transform 1 0 46144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3560__A2
timestamp 1698431365
transform 1 0 45808 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3562__A1
timestamp 1698431365
transform 1 0 38864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3562__A2
timestamp 1698431365
transform -1 0 36848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3563__A1
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3563__A2
timestamp 1698431365
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3565__I
timestamp 1698431365
transform -1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3566__A2
timestamp 1698431365
transform 1 0 33600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3567__A2
timestamp 1698431365
transform -1 0 31472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3569__A1
timestamp 1698431365
transform 1 0 39984 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3569__A2
timestamp 1698431365
transform 1 0 39536 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3571__I0
timestamp 1698431365
transform -1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3574__A1
timestamp 1698431365
transform 1 0 52080 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3574__A2
timestamp 1698431365
transform 1 0 51632 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3574__B
timestamp 1698431365
transform -1 0 50848 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3577__A1
timestamp 1698431365
transform -1 0 60816 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3577__A2
timestamp 1698431365
transform 1 0 61712 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3579__A1
timestamp 1698431365
transform 1 0 44912 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3579__A2
timestamp 1698431365
transform 1 0 44240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3579__B
timestamp 1698431365
transform -1 0 44016 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3582__A1
timestamp 1698431365
transform -1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3582__A2
timestamp 1698431365
transform 1 0 62048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3584__A2
timestamp 1698431365
transform -1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3587__A1
timestamp 1698431365
transform 1 0 40992 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3587__A2
timestamp 1698431365
transform 1 0 2912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3587__B
timestamp 1698431365
transform -1 0 6160 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3592__I1
timestamp 1698431365
transform 1 0 38976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3594__A2
timestamp 1698431365
transform 1 0 39200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3595__A1
timestamp 1698431365
transform 1 0 39760 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3595__A2
timestamp 1698431365
transform -1 0 37744 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3595__B
timestamp 1698431365
transform 1 0 40208 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3597__A1
timestamp 1698431365
transform 1 0 40992 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3597__A2
timestamp 1698431365
transform 1 0 41440 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3600__A2
timestamp 1698431365
transform -1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3602__I1
timestamp 1698431365
transform 1 0 11760 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3605__A1
timestamp 1698431365
transform -1 0 4144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3605__A2
timestamp 1698431365
transform -1 0 3696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3605__B
timestamp 1698431365
transform -1 0 4032 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3611__A1
timestamp 1698431365
transform 1 0 9072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3611__A2
timestamp 1698431365
transform -1 0 12208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3611__B
timestamp 1698431365
transform -1 0 9744 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3613__I0
timestamp 1698431365
transform -1 0 10640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3614__A2
timestamp 1698431365
transform 1 0 12656 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3616__A2
timestamp 1698431365
transform 1 0 27664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3619__A2
timestamp 1698431365
transform 1 0 37072 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3621__A1
timestamp 1698431365
transform 1 0 10304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3621__A2
timestamp 1698431365
transform -1 0 2016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3624__A2
timestamp 1698431365
transform 1 0 11760 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3629__A1
timestamp 1698431365
transform -1 0 6048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3629__A2
timestamp 1698431365
transform -1 0 7168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3635__I1
timestamp 1698431365
transform -1 0 10640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3635__S
timestamp 1698431365
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3640__A2
timestamp 1698431365
transform 1 0 22960 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3640__C
timestamp 1698431365
transform -1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3641__A1
timestamp 1698431365
transform 1 0 9856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3645__I1
timestamp 1698431365
transform -1 0 3696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3645__S
timestamp 1698431365
transform 1 0 15344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3647__A2
timestamp 1698431365
transform 1 0 2800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3656__I0
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3657__A2
timestamp 1698431365
transform -1 0 4032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3657__C
timestamp 1698431365
transform -1 0 11872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3658__A1
timestamp 1698431365
transform -1 0 2128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3658__A2
timestamp 1698431365
transform -1 0 16352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3662__A2
timestamp 1698431365
transform -1 0 30800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3662__C
timestamp 1698431365
transform -1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3663__A1
timestamp 1698431365
transform 1 0 48832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3667__A2
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3667__C
timestamp 1698431365
transform 1 0 20272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3668__A1
timestamp 1698431365
transform -1 0 21168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3668__A2
timestamp 1698431365
transform -1 0 23072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3671__A1
timestamp 1698431365
transform 1 0 15456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3671__A2
timestamp 1698431365
transform 1 0 16352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3671__B
timestamp 1698431365
transform -1 0 16128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3678__I1
timestamp 1698431365
transform -1 0 46928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3678__S
timestamp 1698431365
transform 1 0 49952 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3683__C
timestamp 1698431365
transform 1 0 45360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3684__A1
timestamp 1698431365
transform 1 0 57344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3688__I1
timestamp 1698431365
transform -1 0 46144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3688__S
timestamp 1698431365
transform 1 0 47600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3691__A1
timestamp 1698431365
transform 1 0 23632 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3691__A2
timestamp 1698431365
transform 1 0 24976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3691__B
timestamp 1698431365
transform 1 0 24080 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3701__I1
timestamp 1698431365
transform 1 0 57792 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3704__A1
timestamp 1698431365
transform -1 0 57232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3704__A2
timestamp 1698431365
transform -1 0 57680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3710__A1
timestamp 1698431365
transform -1 0 50064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3710__A2
timestamp 1698431365
transform 1 0 60704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3711__A1
timestamp 1698431365
transform 1 0 60256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3717__A1
timestamp 1698431365
transform 1 0 27888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3717__A2
timestamp 1698431365
transform -1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3718__A1
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3718__A2
timestamp 1698431365
transform 1 0 46032 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3718__B
timestamp 1698431365
transform 1 0 50624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3725__A2
timestamp 1698431365
transform 1 0 62160 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3726__A1
timestamp 1698431365
transform -1 0 61936 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3727__A1
timestamp 1698431365
transform -1 0 52304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3727__A2
timestamp 1698431365
transform 1 0 61824 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3737__A2
timestamp 1698431365
transform 1 0 51072 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3738__A1
timestamp 1698431365
transform -1 0 47264 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3740__A2
timestamp 1698431365
transform -1 0 43680 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3742__A1
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3742__A2
timestamp 1698431365
transform 1 0 32480 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3744__A2
timestamp 1698431365
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3752__CLK
timestamp 1698431365
transform 1 0 60480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3754__D
timestamp 1698431365
transform 1 0 61040 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3756__CLK
timestamp 1698431365
transform 1 0 61936 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3776__CLK
timestamp 1698431365
transform 1 0 44016 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3782__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3786__CLK
timestamp 1698431365
transform -1 0 14448 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3796__CLK
timestamp 1698431365
transform 1 0 9520 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3802__D
timestamp 1698431365
transform 1 0 40096 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3806__CLK
timestamp 1698431365
transform 1 0 6832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3810__CLK
timestamp 1698431365
transform 1 0 5824 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3816__CLK
timestamp 1698431365
transform -1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3820__CLK
timestamp 1698431365
transform 1 0 4816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3826__CLK
timestamp 1698431365
transform -1 0 7840 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3832__CLK
timestamp 1698431365
transform -1 0 13104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3836__CLK
timestamp 1698431365
transform -1 0 12432 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3842__CLK
timestamp 1698431365
transform -1 0 4368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3846__CLK
timestamp 1698431365
transform 1 0 9072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3852__CLK
timestamp 1698431365
transform 1 0 6832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3866__CLK
timestamp 1698431365
transform -1 0 4368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3870__CLK
timestamp 1698431365
transform -1 0 9968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3880__CLK
timestamp 1698431365
transform 1 0 2800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3890__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3915__D
timestamp 1698431365
transform -1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3926__CLK
timestamp 1698431365
transform -1 0 22064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3932__CLK
timestamp 1698431365
transform -1 0 21616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3936__CLK
timestamp 1698431365
transform -1 0 12544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3942__CLK
timestamp 1698431365
transform 1 0 6272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3950__CLK
timestamp 1698431365
transform 1 0 57344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3956__CLK
timestamp 1698431365
transform -1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3966__CLK
timestamp 1698431365
transform -1 0 50288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3970__CLK
timestamp 1698431365
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3976__CLK
timestamp 1698431365
transform -1 0 46592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3980__CLK
timestamp 1698431365
transform -1 0 26768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3986__CLK
timestamp 1698431365
transform 1 0 58912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3987__D
timestamp 1698431365
transform -1 0 59808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3992__CLK
timestamp 1698431365
transform 1 0 59136 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3996__CLK
timestamp 1698431365
transform -1 0 58128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4002__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4006__CLK
timestamp 1698431365
transform 1 0 54096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4012__CLK
timestamp 1698431365
transform 1 0 58016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4016__CLK
timestamp 1698431365
transform 1 0 61040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4022__CLK
timestamp 1698431365
transform 1 0 26096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4026__CLK
timestamp 1698431365
transform -1 0 47264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4030__CLK
timestamp 1698431365
transform 1 0 60256 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4036__CLK
timestamp 1698431365
transform 1 0 61488 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4040__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4046__CLK
timestamp 1698431365
transform 1 0 59136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4050__CLK
timestamp 1698431365
transform 1 0 44800 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4056__CLK
timestamp 1698431365
transform 1 0 41776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__4060__CLK
timestamp 1698431365
transform 1 0 47040 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout42_I
timestamp 1698431365
transform 1 0 61488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout90_I
timestamp 1698431365
transform -1 0 40208 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout106_I
timestamp 1698431365
transform 1 0 58240 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout110_I
timestamp 1698431365
transform -1 0 2128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout111_I
timestamp 1698431365
transform 1 0 1904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout113_I
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout114_I
timestamp 1698431365
transform -1 0 15904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout115_I
timestamp 1698431365
transform -1 0 2576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout116_I
timestamp 1698431365
transform -1 0 2912 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout117_I
timestamp 1698431365
transform -1 0 2016 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout118_I
timestamp 1698431365
transform -1 0 11760 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout119_I
timestamp 1698431365
transform -1 0 11312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout120_I
timestamp 1698431365
transform -1 0 2464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout121_I
timestamp 1698431365
transform 1 0 2912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout122_I
timestamp 1698431365
transform -1 0 18704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout123_I
timestamp 1698431365
transform 1 0 51968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout124_I
timestamp 1698431365
transform 1 0 51072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout125_I
timestamp 1698431365
transform 1 0 59360 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout126_I
timestamp 1698431365
transform 1 0 46144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout127_I
timestamp 1698431365
transform 1 0 37968 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout128_I
timestamp 1698431365
transform -1 0 41888 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout129_I
timestamp 1698431365
transform 1 0 41216 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout130_I
timestamp 1698431365
transform -1 0 50736 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout131_I
timestamp 1698431365
transform -1 0 47712 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout132_I
timestamp 1698431365
transform -1 0 38640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout133_I
timestamp 1698431365
transform 1 0 36848 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 2464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 62384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 59696 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 26656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 27104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 62272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 61824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 61936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 47936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 61712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 26208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 25760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 3024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 2128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 1792 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 34944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output20_I
timestamp 1698431365
transform 1 0 48048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output21_I
timestamp 1698431365
transform -1 0 2800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout27
timestamp 1698431365
transform -1 0 37184 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout28
timestamp 1698431365
transform 1 0 37968 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout29
timestamp 1698431365
transform -1 0 49280 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout30
timestamp 1698431365
transform -1 0 46032 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout31
timestamp 1698431365
transform -1 0 53872 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout32
timestamp 1698431365
transform -1 0 62272 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout33
timestamp 1698431365
transform -1 0 62384 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout34
timestamp 1698431365
transform 1 0 61600 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout35
timestamp 1698431365
transform 1 0 31136 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout36
timestamp 1698431365
transform 1 0 38640 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout37
timestamp 1698431365
transform 1 0 37296 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout38
timestamp 1698431365
transform -1 0 57120 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout39
timestamp 1698431365
transform -1 0 53312 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout40
timestamp 1698431365
transform 1 0 61040 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout41
timestamp 1698431365
transform -1 0 61376 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout42
timestamp 1698431365
transform -1 0 54768 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout43
timestamp 1698431365
transform -1 0 54096 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout44
timestamp 1698431365
transform -1 0 26208 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout45
timestamp 1698431365
transform -1 0 28560 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout46
timestamp 1698431365
transform 1 0 41104 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout47
timestamp 1698431365
transform 1 0 44128 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout48
timestamp 1698431365
transform -1 0 50512 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout49
timestamp 1698431365
transform 1 0 39872 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout50
timestamp 1698431365
transform 1 0 41216 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout51
timestamp 1698431365
transform -1 0 45136 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout52
timestamp 1698431365
transform -1 0 54880 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout53
timestamp 1698431365
transform -1 0 14000 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout54
timestamp 1698431365
transform -1 0 14896 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout55
timestamp 1698431365
transform -1 0 21840 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout56
timestamp 1698431365
transform -1 0 25200 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout57
timestamp 1698431365
transform -1 0 25984 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout58
timestamp 1698431365
transform 1 0 21952 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout59
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout60
timestamp 1698431365
transform -1 0 36288 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout61
timestamp 1698431365
transform 1 0 21168 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout62
timestamp 1698431365
transform -1 0 22064 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout63
timestamp 1698431365
transform -1 0 21840 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout64
timestamp 1698431365
transform -1 0 5936 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout65
timestamp 1698431365
transform -1 0 5264 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout66
timestamp 1698431365
transform -1 0 11648 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout67
timestamp 1698431365
transform 1 0 14784 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout68
timestamp 1698431365
transform 1 0 16800 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout69
timestamp 1698431365
transform -1 0 12208 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout70
timestamp 1698431365
transform 1 0 21504 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout71
timestamp 1698431365
transform 1 0 17360 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout72
timestamp 1698431365
transform -1 0 20944 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout73
timestamp 1698431365
transform -1 0 27888 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout74
timestamp 1698431365
transform -1 0 9968 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout75
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout76
timestamp 1698431365
transform -1 0 12320 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout77
timestamp 1698431365
transform 1 0 16352 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout78
timestamp 1698431365
transform 1 0 15680 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout79
timestamp 1698431365
transform -1 0 20048 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout80
timestamp 1698431365
transform -1 0 27216 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout81
timestamp 1698431365
transform -1 0 29008 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout82
timestamp 1698431365
transform -1 0 18368 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout83
timestamp 1698431365
transform -1 0 13104 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout84
timestamp 1698431365
transform 1 0 13664 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout85
timestamp 1698431365
transform -1 0 5152 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout86
timestamp 1698431365
transform -1 0 3696 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout87
timestamp 1698431365
transform 1 0 9072 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout88
timestamp 1698431365
transform 1 0 12432 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout89
timestamp 1698431365
transform -1 0 17472 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout90
timestamp 1698431365
transform -1 0 41440 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout91
timestamp 1698431365
transform 1 0 37968 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout92
timestamp 1698431365
transform -1 0 35280 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout93
timestamp 1698431365
transform -1 0 35728 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout94
timestamp 1698431365
transform -1 0 29680 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout95
timestamp 1698431365
transform -1 0 29680 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout96
timestamp 1698431365
transform 1 0 32928 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout97
timestamp 1698431365
transform 1 0 33824 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout98
timestamp 1698431365
transform -1 0 38416 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout99
timestamp 1698431365
transform 1 0 38416 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout100
timestamp 1698431365
transform -1 0 47040 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout101
timestamp 1698431365
transform -1 0 45472 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout102
timestamp 1698431365
transform -1 0 43568 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout103
timestamp 1698431365
transform -1 0 48608 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout104
timestamp 1698431365
transform -1 0 58016 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout105
timestamp 1698431365
transform -1 0 59024 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout106
timestamp 1698431365
transform -1 0 57568 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout107
timestamp 1698431365
transform -1 0 59808 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout108
timestamp 1698431365
transform -1 0 46032 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout109
timestamp 1698431365
transform 1 0 46032 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout110
timestamp 1698431365
transform -1 0 4032 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout111
timestamp 1698431365
transform 1 0 1680 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout112
timestamp 1698431365
transform 1 0 16352 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout113
timestamp 1698431365
transform -1 0 23968 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout114
timestamp 1698431365
transform 1 0 15456 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout115
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout116
timestamp 1698431365
transform -1 0 2240 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout117
timestamp 1698431365
transform 1 0 2240 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout118
timestamp 1698431365
transform 1 0 14000 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout119
timestamp 1698431365
transform 1 0 14112 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout120
timestamp 1698431365
transform -1 0 2240 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout121
timestamp 1698431365
transform -1 0 2912 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout122
timestamp 1698431365
transform 1 0 33040 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout123
timestamp 1698431365
transform -1 0 35392 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout124
timestamp 1698431365
transform 1 0 48608 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout125
timestamp 1698431365
transform -1 0 51968 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout126
timestamp 1698431365
transform 1 0 34048 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout127
timestamp 1698431365
transform 1 0 32032 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout128
timestamp 1698431365
transform -1 0 41440 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout129
timestamp 1698431365
transform -1 0 42112 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout130
timestamp 1698431365
transform 1 0 49504 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout131
timestamp 1698431365
transform 1 0 49616 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout132
timestamp 1698431365
transform 1 0 35392 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout133
timestamp 1698431365
transform 1 0 32704 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout134
timestamp 1698431365
transform 1 0 2912 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_36 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_52 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_54 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7392 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_59 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7952 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_188
timestamp 1698431365
transform 1 0 22400 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_196
timestamp 1698431365
transform 1 0 23296 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_199
timestamp 1698431365
transform 1 0 23632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_210
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_214
timestamp 1698431365
transform 1 0 25312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_218
timestamp 1698431365
transform 1 0 25760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_222
timestamp 1698431365
transform 1 0 26208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_226
timestamp 1698431365
transform 1 0 26656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_230
timestamp 1698431365
transform 1 0 27104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_234
timestamp 1698431365
transform 1 0 27552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_240 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_244
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_247
timestamp 1698431365
transform 1 0 29008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_259
timestamp 1698431365
transform 1 0 30352 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_263
timestamp 1698431365
transform 1 0 30800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_302
timestamp 1698431365
transform 1 0 35168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_333
timestamp 1698431365
transform 1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_337
timestamp 1698431365
transform 1 0 39088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_371
timestamp 1698431365
transform 1 0 42896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_373
timestamp 1698431365
transform 1 0 43120 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_380
timestamp 1698431365
transform 1 0 43904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_388
timestamp 1698431365
transform 1 0 44800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_392
timestamp 1698431365
transform 1 0 45248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_396
timestamp 1698431365
transform 1 0 45696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_400
timestamp 1698431365
transform 1 0 46144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_404
timestamp 1698431365
transform 1 0 46592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_414
timestamp 1698431365
transform 1 0 47712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_418
timestamp 1698431365
transform 1 0 48160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_422
timestamp 1698431365
transform 1 0 48608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_438
timestamp 1698431365
transform 1 0 50400 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_512
timestamp 1698431365
transform 1 0 58688 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_544
timestamp 1698431365
transform 1 0 62272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_174
timestamp 1698431365
transform 1 0 20832 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_177
timestamp 1698431365
transform 1 0 21168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_181
timestamp 1698431365
transform 1 0 21616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_185
timestamp 1698431365
transform 1 0 22064 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_189
timestamp 1698431365
transform 1 0 22512 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_192
timestamp 1698431365
transform 1 0 22848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_196
timestamp 1698431365
transform 1 0 23296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_200
timestamp 1698431365
transform 1 0 23744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_202
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_205
timestamp 1698431365
transform 1 0 24304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_216
timestamp 1698431365
transform 1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_224
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_227
timestamp 1698431365
transform 1 0 26768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_231
timestamp 1698431365
transform 1 0 27216 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_235
timestamp 1698431365
transform 1 0 27664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_239
timestamp 1698431365
transform 1 0 28112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_243
timestamp 1698431365
transform 1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_247
timestamp 1698431365
transform 1 0 29008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_271
timestamp 1698431365
transform 1 0 31696 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_372
timestamp 1698431365
transform 1 0 43008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_374
timestamp 1698431365
transform 1 0 43232 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_403
timestamp 1698431365
transform 1 0 46480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_407
timestamp 1698431365
transform 1 0 46928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_411
timestamp 1698431365
transform 1 0 47376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_415
timestamp 1698431365
transform 1 0 47824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_419
timestamp 1698431365
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_426
timestamp 1698431365
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_430
timestamp 1698431365
transform 1 0 49504 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_462
timestamp 1698431365
transform 1 0 53088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_478
timestamp 1698431365
transform 1 0 54880 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_524
timestamp 1698431365
transform 1 0 60032 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_540
timestamp 1698431365
transform 1 0 61824 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_544
timestamp 1698431365
transform 1 0 62272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_113
timestamp 1698431365
transform 1 0 14000 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_121
timestamp 1698431365
transform 1 0 14896 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_125
timestamp 1698431365
transform 1 0 15344 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_128
timestamp 1698431365
transform 1 0 15680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_132
timestamp 1698431365
transform 1 0 16128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_136
timestamp 1698431365
transform 1 0 16576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_138
timestamp 1698431365
transform 1 0 16800 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_141
timestamp 1698431365
transform 1 0 17136 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_149
timestamp 1698431365
transform 1 0 18032 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_153
timestamp 1698431365
transform 1 0 18480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_157
timestamp 1698431365
transform 1 0 18928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_159
timestamp 1698431365
transform 1 0 19152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_162
timestamp 1698431365
transform 1 0 19488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_164
timestamp 1698431365
transform 1 0 19712 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_167
timestamp 1698431365
transform 1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_181
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_185
timestamp 1698431365
transform 1 0 22064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_187
timestamp 1698431365
transform 1 0 22288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_190
timestamp 1698431365
transform 1 0 22624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_194
timestamp 1698431365
transform 1 0 23072 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_198
timestamp 1698431365
transform 1 0 23520 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_201
timestamp 1698431365
transform 1 0 23856 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_205
timestamp 1698431365
transform 1 0 24304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_209
timestamp 1698431365
transform 1 0 24752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_213
timestamp 1698431365
transform 1 0 25200 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_219
timestamp 1698431365
transform 1 0 25872 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_223
timestamp 1698431365
transform 1 0 26320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_227
timestamp 1698431365
transform 1 0 26768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698431365
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_312
timestamp 1698431365
transform 1 0 36288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698431365
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_346
timestamp 1698431365
transform 1 0 40096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_402
timestamp 1698431365
transform 1 0 46368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_433
timestamp 1698431365
transform 1 0 49840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_437
timestamp 1698431365
transform 1 0 50288 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_453
timestamp 1698431365
transform 1 0 52080 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_521
timestamp 1698431365
transform 1 0 59696 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_527
timestamp 1698431365
transform 1 0 60368 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_543
timestamp 1698431365
transform 1 0 62160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_88
timestamp 1698431365
transform 1 0 11200 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_96
timestamp 1698431365
transform 1 0 12096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_100
timestamp 1698431365
transform 1 0 12544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_104
timestamp 1698431365
transform 1 0 12992 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_113
timestamp 1698431365
transform 1 0 14000 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_115
timestamp 1698431365
transform 1 0 14224 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_118
timestamp 1698431365
transform 1 0 14560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_122
timestamp 1698431365
transform 1 0 15008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_126
timestamp 1698431365
transform 1 0 15456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_130
timestamp 1698431365
transform 1 0 15904 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_172
timestamp 1698431365
transform 1 0 20608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_176
timestamp 1698431365
transform 1 0 21056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_180
timestamp 1698431365
transform 1 0 21504 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_186
timestamp 1698431365
transform 1 0 22176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_190
timestamp 1698431365
transform 1 0 22624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_194
timestamp 1698431365
transform 1 0 23072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_196
timestamp 1698431365
transform 1 0 23296 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_199
timestamp 1698431365
transform 1 0 23632 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_203
timestamp 1698431365
transform 1 0 24080 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_251
timestamp 1698431365
transform 1 0 29456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_253
timestamp 1698431365
transform 1 0 29680 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_348
timestamp 1698431365
transform 1 0 40320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_354
timestamp 1698431365
transform 1 0 40992 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_410
timestamp 1698431365
transform 1 0 47264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_414
timestamp 1698431365
transform 1 0 47712 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_419
timestamp 1698431365
transform 1 0 48272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_427
timestamp 1698431365
transform 1 0 49168 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_431
timestamp 1698431365
transform 1 0 49616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_435
timestamp 1698431365
transform 1 0 50064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_439
timestamp 1698431365
transform 1 0 50512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_443
timestamp 1698431365
transform 1 0 50960 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_475
timestamp 1698431365
transform 1 0 54544 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_483
timestamp 1698431365
transform 1 0 55440 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_487
timestamp 1698431365
transform 1 0 55888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_489
timestamp 1698431365
transform 1 0 56112 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_524
timestamp 1698431365
transform 1 0 60032 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_540
timestamp 1698431365
transform 1 0 61824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_544
timestamp 1698431365
transform 1 0 62272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_69
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_71
timestamp 1698431365
transform 1 0 9296 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_95
timestamp 1698431365
transform 1 0 11984 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_113
timestamp 1698431365
transform 1 0 14000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_121
timestamp 1698431365
transform 1 0 14896 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_127
timestamp 1698431365
transform 1 0 15568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_131
timestamp 1698431365
transform 1 0 16016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_140
timestamp 1698431365
transform 1 0 17024 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_189
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_191
timestamp 1698431365
transform 1 0 22736 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_197
timestamp 1698431365
transform 1 0 23408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_199
timestamp 1698431365
transform 1 0 23632 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_202
timestamp 1698431365
transform 1 0 23968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_206
timestamp 1698431365
transform 1 0 24416 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_210
timestamp 1698431365
transform 1 0 24864 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_237
timestamp 1698431365
transform 1 0 27888 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_249
timestamp 1698431365
transform 1 0 29232 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_260
timestamp 1698431365
transform 1 0 30464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_262
timestamp 1698431365
transform 1 0 30688 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_371
timestamp 1698431365
transform 1 0 42896 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_403
timestamp 1698431365
transform 1 0 46480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_405
timestamp 1698431365
transform 1 0 46704 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_439
timestamp 1698431365
transform 1 0 50512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_443
timestamp 1698431365
transform 1 0 50960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_447
timestamp 1698431365
transform 1 0 51408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_521
timestamp 1698431365
transform 1 0 59696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_527
timestamp 1698431365
transform 1 0 60368 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_543
timestamp 1698431365
transform 1 0 62160 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_50
timestamp 1698431365
transform 1 0 6944 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_58
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_65
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_162
timestamp 1698431365
transform 1 0 19488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_207
timestamp 1698431365
transform 1 0 24528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_240
timestamp 1698431365
transform 1 0 28224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_270
timestamp 1698431365
transform 1 0 31584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_299
timestamp 1698431365
transform 1 0 34832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_301
timestamp 1698431365
transform 1 0 35056 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_368
timestamp 1698431365
transform 1 0 42560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_388
timestamp 1698431365
transform 1 0 44800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_392
timestamp 1698431365
transform 1 0 45248 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_442
timestamp 1698431365
transform 1 0 50848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_446
timestamp 1698431365
transform 1 0 51296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_450
timestamp 1698431365
transform 1 0 51744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_454
timestamp 1698431365
transform 1 0 52192 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_458
timestamp 1698431365
transform 1 0 52640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_462
timestamp 1698431365
transform 1 0 53088 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_478
timestamp 1698431365
transform 1 0 54880 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_524
timestamp 1698431365
transform 1 0 60032 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_540
timestamp 1698431365
transform 1 0 61824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_544
timestamp 1698431365
transform 1 0 62272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_53
timestamp 1698431365
transform 1 0 7280 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_87
timestamp 1698431365
transform 1 0 11088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_89
timestamp 1698431365
transform 1 0 11312 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_127
timestamp 1698431365
transform 1 0 15568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_206
timestamp 1698431365
transform 1 0 24416 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_237
timestamp 1698431365
transform 1 0 27888 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_299
timestamp 1698431365
transform 1 0 34832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_352
timestamp 1698431365
transform 1 0 40768 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_383
timestamp 1698431365
transform 1 0 44240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_450
timestamp 1698431365
transform 1 0 51744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_454
timestamp 1698431365
transform 1 0 52192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_461
timestamp 1698431365
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_465
timestamp 1698431365
transform 1 0 53424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_469
timestamp 1698431365
transform 1 0 53872 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_473
timestamp 1698431365
transform 1 0 54320 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_505
timestamp 1698431365
transform 1 0 57904 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_521
timestamp 1698431365
transform 1 0 59696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_527
timestamp 1698431365
transform 1 0 60368 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_543
timestamp 1698431365
transform 1 0 62160 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_42
timestamp 1698431365
transform 1 0 6048 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_46
timestamp 1698431365
transform 1 0 6496 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_76
timestamp 1698431365
transform 1 0 9856 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_101
timestamp 1698431365
transform 1 0 12656 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_233
timestamp 1698431365
transform 1 0 27440 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_261
timestamp 1698431365
transform 1 0 30576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_273
timestamp 1698431365
transform 1 0 31920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_329
timestamp 1698431365
transform 1 0 38192 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_363
timestamp 1698431365
transform 1 0 42000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_375
timestamp 1698431365
transform 1 0 43344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_379
timestamp 1698431365
transform 1 0 43792 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_397
timestamp 1698431365
transform 1 0 45808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_465
timestamp 1698431365
transform 1 0 53424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_469
timestamp 1698431365
transform 1 0 53872 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_473
timestamp 1698431365
transform 1 0 54320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_477
timestamp 1698431365
transform 1 0 54768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_485
timestamp 1698431365
transform 1 0 55664 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_489
timestamp 1698431365
transform 1 0 56112 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_524
timestamp 1698431365
transform 1 0 60032 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_540
timestamp 1698431365
transform 1 0 61824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_544
timestamp 1698431365
transform 1 0 62272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_39
timestamp 1698431365
transform 1 0 5712 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_42
timestamp 1698431365
transform 1 0 6048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_46
timestamp 1698431365
transform 1 0 6496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_58
timestamp 1698431365
transform 1 0 7840 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_60
timestamp 1698431365
transform 1 0 8064 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_102
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_109
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_199
timestamp 1698431365
transform 1 0 23632 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_265
timestamp 1698431365
transform 1 0 31024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_269
timestamp 1698431365
transform 1 0 31472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_271
timestamp 1698431365
transform 1 0 31696 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_293
timestamp 1698431365
transform 1 0 34160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_339
timestamp 1698431365
transform 1 0 39312 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_371
timestamp 1698431365
transform 1 0 42896 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_454
timestamp 1698431365
transform 1 0 52192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_477
timestamp 1698431365
transform 1 0 54768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_481
timestamp 1698431365
transform 1 0 55216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_485
timestamp 1698431365
transform 1 0 55664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_489
timestamp 1698431365
transform 1 0 56112 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_493
timestamp 1698431365
transform 1 0 56560 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_527
timestamp 1698431365
transform 1 0 60368 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_543
timestamp 1698431365
transform 1 0 62160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_18
timestamp 1698431365
transform 1 0 3360 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_26
timestamp 1698431365
transform 1 0 4256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_32
timestamp 1698431365
transform 1 0 4928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_36
timestamp 1698431365
transform 1 0 5376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_45
timestamp 1698431365
transform 1 0 6384 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_119
timestamp 1698431365
transform 1 0 14672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_121
timestamp 1698431365
transform 1 0 14896 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_190
timestamp 1698431365
transform 1 0 22624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_203
timestamp 1698431365
transform 1 0 24080 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_277
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_334
timestamp 1698431365
transform 1 0 38752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_336
timestamp 1698431365
transform 1 0 38976 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_341
timestamp 1698431365
transform 1 0 39536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_345
timestamp 1698431365
transform 1 0 39984 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_369
timestamp 1698431365
transform 1 0 42672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_399
timestamp 1698431365
transform 1 0 46032 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_401
timestamp 1698431365
transform 1 0 46256 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_488
timestamp 1698431365
transform 1 0 56000 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_496
timestamp 1698431365
transform 1 0 56896 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_500
timestamp 1698431365
transform 1 0 57344 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_532
timestamp 1698431365
transform 1 0 60928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_540
timestamp 1698431365
transform 1 0 61824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_544
timestamp 1698431365
transform 1 0 62272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_12
timestamp 1698431365
transform 1 0 2688 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_88
timestamp 1698431365
transform 1 0 11200 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_129
timestamp 1698431365
transform 1 0 15792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_131
timestamp 1698431365
transform 1 0 16016 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_214
timestamp 1698431365
transform 1 0 25312 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_255
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_257
timestamp 1698431365
transform 1 0 30128 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_277
timestamp 1698431365
transform 1 0 32368 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_304
timestamp 1698431365
transform 1 0 35392 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_306
timestamp 1698431365
transform 1 0 35616 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_353
timestamp 1698431365
transform 1 0 40880 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_403
timestamp 1698431365
transform 1 0 46480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_454
timestamp 1698431365
transform 1 0 52192 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_487
timestamp 1698431365
transform 1 0 55888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_491
timestamp 1698431365
transform 1 0 56336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_495
timestamp 1698431365
transform 1 0 56784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_499
timestamp 1698431365
transform 1 0 57232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_503
timestamp 1698431365
transform 1 0 57680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_507
timestamp 1698431365
transform 1 0 58128 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_523
timestamp 1698431365
transform 1 0 59920 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_527
timestamp 1698431365
transform 1 0 60368 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_543
timestamp 1698431365
transform 1 0 62160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_8
timestamp 1698431365
transform 1 0 2240 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_12
timestamp 1698431365
transform 1 0 2688 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_15
timestamp 1698431365
transform 1 0 3024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_19
timestamp 1698431365
transform 1 0 3472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_95
timestamp 1698431365
transform 1 0 11984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_97
timestamp 1698431365
transform 1 0 12208 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_183
timestamp 1698431365
transform 1 0 21840 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_354
timestamp 1698431365
transform 1 0 40992 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_430
timestamp 1698431365
transform 1 0 49504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_434
timestamp 1698431365
transform 1 0 49952 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_488
timestamp 1698431365
transform 1 0 56000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_498
timestamp 1698431365
transform 1 0 57120 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_502
timestamp 1698431365
transform 1 0 57568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_506
timestamp 1698431365
transform 1 0 58016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_510
timestamp 1698431365
transform 1 0 58464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_514
timestamp 1698431365
transform 1 0 58912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_518
timestamp 1698431365
transform 1 0 59360 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_522
timestamp 1698431365
transform 1 0 59808 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_538
timestamp 1698431365
transform 1 0 61600 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_542
timestamp 1698431365
transform 1 0 62048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_544
timestamp 1698431365
transform 1 0 62272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_4
timestamp 1698431365
transform 1 0 1792 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_7
timestamp 1698431365
transform 1 0 2128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_11
timestamp 1698431365
transform 1 0 2576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_145
timestamp 1698431365
transform 1 0 17584 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_313
timestamp 1698431365
transform 1 0 36400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_391
timestamp 1698431365
transform 1 0 45136 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_395
timestamp 1698431365
transform 1 0 45584 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_397
timestamp 1698431365
transform 1 0 45808 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_432
timestamp 1698431365
transform 1 0 49728 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_454
timestamp 1698431365
transform 1 0 52192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_494
timestamp 1698431365
transform 1 0 56672 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_498
timestamp 1698431365
transform 1 0 57120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_502
timestamp 1698431365
transform 1 0 57568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_506
timestamp 1698431365
transform 1 0 58016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_510
timestamp 1698431365
transform 1 0 58464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_514
timestamp 1698431365
transform 1 0 58912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_518
timestamp 1698431365
transform 1 0 59360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_522
timestamp 1698431365
transform 1 0 59808 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_524
timestamp 1698431365
transform 1 0 60032 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_527
timestamp 1698431365
transform 1 0 60368 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_535
timestamp 1698431365
transform 1 0 61264 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_541
timestamp 1698431365
transform 1 0 61936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_6
timestamp 1698431365
transform 1 0 2016 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_9
timestamp 1698431365
transform 1 0 2352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_13
timestamp 1698431365
transform 1 0 2800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_17
timestamp 1698431365
transform 1 0 3248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_60
timestamp 1698431365
transform 1 0 8064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_87
timestamp 1698431365
transform 1 0 11088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_89
timestamp 1698431365
transform 1 0 11312 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_119
timestamp 1698431365
transform 1 0 14672 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_152
timestamp 1698431365
transform 1 0 18368 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_189
timestamp 1698431365
transform 1 0 22512 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_274
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_333
timestamp 1698431365
transform 1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_413
timestamp 1698431365
transform 1 0 47600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_417
timestamp 1698431365
transform 1 0 48048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_419
timestamp 1698431365
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_438
timestamp 1698431365
transform 1 0 50400 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_442
timestamp 1698431365
transform 1 0 50848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_444
timestamp 1698431365
transform 1 0 51072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_460
timestamp 1698431365
transform 1 0 52864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_462
timestamp 1698431365
transform 1 0 53088 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_487
timestamp 1698431365
transform 1 0 55888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_489
timestamp 1698431365
transform 1 0 56112 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_500
timestamp 1698431365
transform 1 0 57344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_504
timestamp 1698431365
transform 1 0 57792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_512
timestamp 1698431365
transform 1 0 58688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_516
timestamp 1698431365
transform 1 0 59136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_520
timestamp 1698431365
transform 1 0 59584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_524
timestamp 1698431365
transform 1 0 60032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_528
timestamp 1698431365
transform 1 0 60480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_532
timestamp 1698431365
transform 1 0 60928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_536
timestamp 1698431365
transform 1 0 61376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_540
timestamp 1698431365
transform 1 0 61824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_544
timestamp 1698431365
transform 1 0 62272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_4
timestamp 1698431365
transform 1 0 1792 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_7
timestamp 1698431365
transform 1 0 2128 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_11
timestamp 1698431365
transform 1 0 2576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_15
timestamp 1698431365
transform 1 0 3024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_19
timestamp 1698431365
transform 1 0 3472 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_23
timestamp 1698431365
transform 1 0 3920 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698431365
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_150
timestamp 1698431365
transform 1 0 18144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_152
timestamp 1698431365
transform 1 0 18368 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_236
timestamp 1698431365
transform 1 0 27776 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_291
timestamp 1698431365
transform 1 0 33936 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_312
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_349
timestamp 1698431365
transform 1 0 40432 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_351
timestamp 1698431365
transform 1 0 40656 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_450
timestamp 1698431365
transform 1 0 51744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_454
timestamp 1698431365
transform 1 0 52192 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_514
timestamp 1698431365
transform 1 0 58912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_518
timestamp 1698431365
transform 1 0 59360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_522
timestamp 1698431365
transform 1 0 59808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_524
timestamp 1698431365
transform 1 0 60032 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_527
timestamp 1698431365
transform 1 0 60368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_531
timestamp 1698431365
transform 1 0 60816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_535
timestamp 1698431365
transform 1 0 61264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_539
timestamp 1698431365
transform 1 0 61712 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_4
timestamp 1698431365
transform 1 0 1792 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_7
timestamp 1698431365
transform 1 0 2128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_11
timestamp 1698431365
transform 1 0 2576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_15
timestamp 1698431365
transform 1 0 3024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_19
timestamp 1698431365
transform 1 0 3472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_23
timestamp 1698431365
transform 1 0 3920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_59
timestamp 1698431365
transform 1 0 7952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_61
timestamp 1698431365
transform 1 0 8176 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_97
timestamp 1698431365
transform 1 0 12208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_152
timestamp 1698431365
transform 1 0 18368 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_175
timestamp 1698431365
transform 1 0 20944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_192
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_218
timestamp 1698431365
transform 1 0 25760 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_220
timestamp 1698431365
transform 1 0 25984 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_254
timestamp 1698431365
transform 1 0 29792 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698431365
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_297
timestamp 1698431365
transform 1 0 34608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_299
timestamp 1698431365
transform 1 0 34832 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_354
timestamp 1698431365
transform 1 0 40992 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_418
timestamp 1698431365
transform 1 0 48160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_473
timestamp 1698431365
transform 1 0 54320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_521
timestamp 1698431365
transform 1 0 59696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_525
timestamp 1698431365
transform 1 0 60144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_529
timestamp 1698431365
transform 1 0 60592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_533
timestamp 1698431365
transform 1 0 61040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_537
timestamp 1698431365
transform 1 0 61488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_541
timestamp 1698431365
transform 1 0 61936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_6
timestamp 1698431365
transform 1 0 2016 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_9
timestamp 1698431365
transform 1 0 2352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_13
timestamp 1698431365
transform 1 0 2800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_17
timestamp 1698431365
transform 1 0 3248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_91
timestamp 1698431365
transform 1 0 11536 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_93
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_164
timestamp 1698431365
transform 1 0 19712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_166
timestamp 1698431365
transform 1 0 19936 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_229
timestamp 1698431365
transform 1 0 26992 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_259
timestamp 1698431365
transform 1 0 30352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_397
timestamp 1698431365
transform 1 0 45808 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_422
timestamp 1698431365
transform 1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_445
timestamp 1698431365
transform 1 0 51184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_449
timestamp 1698431365
transform 1 0 51632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_453
timestamp 1698431365
transform 1 0 52080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_497
timestamp 1698431365
transform 1 0 57008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_499
timestamp 1698431365
transform 1 0 57232 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_524
timestamp 1698431365
transform 1 0 60032 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_527
timestamp 1698431365
transform 1 0 60368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_531
timestamp 1698431365
transform 1 0 60816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_535
timestamp 1698431365
transform 1 0 61264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_539
timestamp 1698431365
transform 1 0 61712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_543
timestamp 1698431365
transform 1 0 62160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_8
timestamp 1698431365
transform 1 0 2240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_12
timestamp 1698431365
transform 1 0 2688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_16
timestamp 1698431365
transform 1 0 3136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_20
timestamp 1698431365
transform 1 0 3584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_24
timestamp 1698431365
transform 1 0 4032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_28
timestamp 1698431365
transform 1 0 4480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_76
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_107
timestamp 1698431365
transform 1 0 13328 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_109
timestamp 1698431365
transform 1 0 13552 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_256
timestamp 1698431365
transform 1 0 30016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_313
timestamp 1698431365
transform 1 0 36400 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_317
timestamp 1698431365
transform 1 0 36848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_354
timestamp 1698431365
transform 1 0 40992 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_398
timestamp 1698431365
transform 1 0 45920 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_417
timestamp 1698431365
transform 1 0 48048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_430
timestamp 1698431365
transform 1 0 49504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_471
timestamp 1698431365
transform 1 0 54096 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_525
timestamp 1698431365
transform 1 0 60144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_4
timestamp 1698431365
transform 1 0 1792 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_7
timestamp 1698431365
transform 1 0 2128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_11
timestamp 1698431365
transform 1 0 2576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_86
timestamp 1698431365
transform 1 0 10976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_147
timestamp 1698431365
transform 1 0 17808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_255
timestamp 1698431365
transform 1 0 29904 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_304
timestamp 1698431365
transform 1 0 35392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_333
timestamp 1698431365
transform 1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_337
timestamp 1698431365
transform 1 0 39088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_350
timestamp 1698431365
transform 1 0 40544 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_384
timestamp 1698431365
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_391
timestamp 1698431365
transform 1 0 45136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_445
timestamp 1698431365
transform 1 0 51184 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_447
timestamp 1698431365
transform 1 0 51408 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_470
timestamp 1698431365
transform 1 0 53984 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_500
timestamp 1698431365
transform 1 0 57344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_502
timestamp 1698431365
transform 1 0 57568 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_6
timestamp 1698431365
transform 1 0 2016 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_9
timestamp 1698431365
transform 1 0 2352 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_13
timestamp 1698431365
transform 1 0 2800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_17
timestamp 1698431365
transform 1 0 3248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_21
timestamp 1698431365
transform 1 0 3696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_53
timestamp 1698431365
transform 1 0 7280 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_67
timestamp 1698431365
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_116
timestamp 1698431365
transform 1 0 14336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_118
timestamp 1698431365
transform 1 0 14560 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_198
timestamp 1698431365
transform 1 0 23520 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_232
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_234
timestamp 1698431365
transform 1 0 27552 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_270
timestamp 1698431365
transform 1 0 31584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_295
timestamp 1698431365
transform 1 0 34384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_315
timestamp 1698431365
transform 1 0 36624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_319
timestamp 1698431365
transform 1 0 37072 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_375
timestamp 1698431365
transform 1 0 43344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_394
timestamp 1698431365
transform 1 0 45472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_441
timestamp 1698431365
transform 1 0 50736 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_507
timestamp 1698431365
transform 1 0 58128 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_536
timestamp 1698431365
transform 1 0 61376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_538
timestamp 1698431365
transform 1 0 61600 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_4
timestamp 1698431365
transform 1 0 1792 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_192
timestamp 1698431365
transform 1 0 22848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_294
timestamp 1698431365
transform 1 0 34272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_296
timestamp 1698431365
transform 1 0 34496 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_339
timestamp 1698431365
transform 1 0 39312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_341
timestamp 1698431365
transform 1 0 39536 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_374
timestamp 1698431365
transform 1 0 43232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_376
timestamp 1698431365
transform 1 0 43456 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_411
timestamp 1698431365
transform 1 0 47376 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_31
timestamp 1698431365
transform 1 0 4816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_33
timestamp 1698431365
transform 1 0 5040 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_59
timestamp 1698431365
transform 1 0 7952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_61
timestamp 1698431365
transform 1 0 8176 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_257
timestamp 1698431365
transform 1 0 30128 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_354
timestamp 1698431365
transform 1 0 40992 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_418
timestamp 1698431365
transform 1 0 48160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_430
timestamp 1698431365
transform 1 0 49504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_456
timestamp 1698431365
transform 1 0 52416 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_480
timestamp 1698431365
transform 1 0 55104 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_489
timestamp 1698431365
transform 1 0 56112 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_543
timestamp 1698431365
transform 1 0 62160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_66
timestamp 1698431365
transform 1 0 8736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_163
timestamp 1698431365
transform 1 0 19600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_165
timestamp 1698431365
transform 1 0 19824 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_323
timestamp 1698431365
transform 1 0 37520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_342
timestamp 1698431365
transform 1 0 39648 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_355
timestamp 1698431365
transform 1 0 41104 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_362
timestamp 1698431365
transform 1 0 41888 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_450
timestamp 1698431365
transform 1 0 51744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_454
timestamp 1698431365
transform 1 0 52192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_465
timestamp 1698431365
transform 1 0 53424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_524
timestamp 1698431365
transform 1 0 60032 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_22
timestamp 1698431365
transform 1 0 3808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_24
timestamp 1698431365
transform 1 0 4032 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_51
timestamp 1698431365
transform 1 0 7056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_53
timestamp 1698431365
transform 1 0 7280 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_107
timestamp 1698431365
transform 1 0 13328 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_260
timestamp 1698431365
transform 1 0 30464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_262
timestamp 1698431365
transform 1 0 30688 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698431365
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_298
timestamp 1698431365
transform 1 0 34720 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_369
timestamp 1698431365
transform 1 0 42672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_401
timestamp 1698431365
transform 1 0 46256 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_417
timestamp 1698431365
transform 1 0 48048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_419
timestamp 1698431365
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_468
timestamp 1698431365
transform 1 0 53760 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_494
timestamp 1698431365
transform 1 0 56672 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_522
timestamp 1698431365
transform 1 0 59808 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_24
timestamp 1698431365
transform 1 0 4032 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_26
timestamp 1698431365
transform 1 0 4256 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_135
timestamp 1698431365
transform 1 0 16464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_137
timestamp 1698431365
transform 1 0 16688 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_304
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_306
timestamp 1698431365
transform 1 0 35616 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_347
timestamp 1698431365
transform 1 0 40208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_349
timestamp 1698431365
transform 1 0 40432 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_395
timestamp 1698431365
transform 1 0 45584 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_451
timestamp 1698431365
transform 1 0 51856 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_475
timestamp 1698431365
transform 1 0 54544 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_504
timestamp 1698431365
transform 1 0 57792 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_542
timestamp 1698431365
transform 1 0 62048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_544
timestamp 1698431365
transform 1 0 62272 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_45
timestamp 1698431365
transform 1 0 6384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_47
timestamp 1698431365
transform 1 0 6608 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_190
timestamp 1698431365
transform 1 0 22624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_192
timestamp 1698431365
transform 1 0 22848 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_201
timestamp 1698431365
transform 1 0 23856 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_286
timestamp 1698431365
transform 1 0 33376 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_313
timestamp 1698431365
transform 1 0 36400 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_500
timestamp 1698431365
transform 1 0 57344 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_22
timestamp 1698431365
transform 1 0 3808 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_39
timestamp 1698431365
transform 1 0 5712 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_62
timestamp 1698431365
transform 1 0 8288 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_68
timestamp 1698431365
transform 1 0 8960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_77
timestamp 1698431365
transform 1 0 9968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_79
timestamp 1698431365
transform 1 0 10192 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_82
timestamp 1698431365
transform 1 0 10528 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_102
timestamp 1698431365
transform 1 0 12768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_117
timestamp 1698431365
transform 1 0 14448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_265
timestamp 1698431365
transform 1 0 31024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_279
timestamp 1698431365
transform 1 0 32592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_281
timestamp 1698431365
transform 1 0 32816 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_323
timestamp 1698431365
transform 1 0 37520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_423
timestamp 1698431365
transform 1 0 48720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_425
timestamp 1698431365
transform 1 0 48944 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_452
timestamp 1698431365
transform 1 0 51968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_454
timestamp 1698431365
transform 1 0 52192 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_500
timestamp 1698431365
transform 1 0 57344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_502
timestamp 1698431365
transform 1 0 57568 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_542
timestamp 1698431365
transform 1 0 62048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_544
timestamp 1698431365
transform 1 0 62272 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_43
timestamp 1698431365
transform 1 0 6160 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_65
timestamp 1698431365
transform 1 0 8624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_67
timestamp 1698431365
transform 1 0 8848 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_101
timestamp 1698431365
transform 1 0 12656 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_125
timestamp 1698431365
transform 1 0 15344 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_161
timestamp 1698431365
transform 1 0 19376 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_183
timestamp 1698431365
transform 1 0 21840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_201
timestamp 1698431365
transform 1 0 23856 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_266
timestamp 1698431365
transform 1 0 31136 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_304
timestamp 1698431365
transform 1 0 35392 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_76
timestamp 1698431365
transform 1 0 9856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_113
timestamp 1698431365
transform 1 0 14000 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_136
timestamp 1698431365
transform 1 0 16576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_138
timestamp 1698431365
transform 1 0 16800 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_158
timestamp 1698431365
transform 1 0 19040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_295
timestamp 1698431365
transform 1 0 34384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_297
timestamp 1698431365
transform 1 0 34608 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698431365
transform 1 0 36288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_402
timestamp 1698431365
transform 1 0 46368 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_452
timestamp 1698431365
transform 1 0 51968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_490
timestamp 1698431365
transform 1 0 56224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_524
timestamp 1698431365
transform 1 0 60032 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_542
timestamp 1698431365
transform 1 0 62048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_544
timestamp 1698431365
transform 1 0 62272 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_46
timestamp 1698431365
transform 1 0 6496 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_94
timestamp 1698431365
transform 1 0 11872 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_114
timestamp 1698431365
transform 1 0 14112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_214
timestamp 1698431365
transform 1 0 25312 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_225
timestamp 1698431365
transform 1 0 26544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_262
timestamp 1698431365
transform 1 0 30688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_264
timestamp 1698431365
transform 1 0 30912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_286
timestamp 1698431365
transform 1 0 33376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_290
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_292
timestamp 1698431365
transform 1 0 34048 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_303
timestamp 1698431365
transform 1 0 35280 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_325
timestamp 1698431365
transform 1 0 37744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_335
timestamp 1698431365
transform 1 0 38864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_337
timestamp 1698431365
transform 1 0 39088 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_417
timestamp 1698431365
transform 1 0 48048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1698431365
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_438
timestamp 1698431365
transform 1 0 50400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_440
timestamp 1698431365
transform 1 0 50624 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_470
timestamp 1698431365
transform 1 0 53984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_472
timestamp 1698431365
transform 1 0 54208 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_500
timestamp 1698431365
transform 1 0 57344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_504
timestamp 1698431365
transform 1 0 57792 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_69
timestamp 1698431365
transform 1 0 9072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_73
timestamp 1698431365
transform 1 0 9520 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_77
timestamp 1698431365
transform 1 0 9968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_102
timestamp 1698431365
transform 1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_168
timestamp 1698431365
transform 1 0 20160 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_179
timestamp 1698431365
transform 1 0 21392 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_186
timestamp 1698431365
transform 1 0 22176 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_252
timestamp 1698431365
transform 1 0 29568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_288
timestamp 1698431365
transform 1 0 33600 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_310
timestamp 1698431365
transform 1 0 36064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_382
timestamp 1698431365
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_398
timestamp 1698431365
transform 1 0 45920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_402
timestamp 1698431365
transform 1 0 46368 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_502
timestamp 1698431365
transform 1 0 57568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_24
timestamp 1698431365
transform 1 0 4032 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_41
timestamp 1698431365
transform 1 0 5936 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_64
timestamp 1698431365
transform 1 0 8512 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_74
timestamp 1698431365
transform 1 0 9632 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_167
timestamp 1698431365
transform 1 0 20048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_169
timestamp 1698431365
transform 1 0 20272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_229
timestamp 1698431365
transform 1 0 26992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_275
timestamp 1698431365
transform 1 0 32144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_295
timestamp 1698431365
transform 1 0 34384 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_301
timestamp 1698431365
transform 1 0 35056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_303
timestamp 1698431365
transform 1 0 35280 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_318
timestamp 1698431365
transform 1 0 36960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_375
timestamp 1698431365
transform 1 0 43344 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_415
timestamp 1698431365
transform 1 0 47824 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_419
timestamp 1698431365
transform 1 0 48272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_77
timestamp 1698431365
transform 1 0 9968 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_109
timestamp 1698431365
transform 1 0 13552 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_179
timestamp 1698431365
transform 1 0 21392 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_229
timestamp 1698431365
transform 1 0 26992 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_231
timestamp 1698431365
transform 1 0 27216 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_323
timestamp 1698431365
transform 1 0 37520 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_327
timestamp 1698431365
transform 1 0 37968 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_382
timestamp 1698431365
transform 1 0 44128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_401
timestamp 1698431365
transform 1 0 46256 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_488
timestamp 1698431365
transform 1 0 56000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_152
timestamp 1698431365
transform 1 0 18368 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_219
timestamp 1698431365
transform 1 0 25872 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_270
timestamp 1698431365
transform 1 0 31584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_272
timestamp 1698431365
transform 1 0 31808 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_325
timestamp 1698431365
transform 1 0 37744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_339
timestamp 1698431365
transform 1 0 39312 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_341
timestamp 1698431365
transform 1 0 39536 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_360
timestamp 1698431365
transform 1 0 41664 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_430
timestamp 1698431365
transform 1 0 49504 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_22
timestamp 1698431365
transform 1 0 3808 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_24
timestamp 1698431365
transform 1 0 4032 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_85
timestamp 1698431365
transform 1 0 10864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_109
timestamp 1698431365
transform 1 0 13552 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_151
timestamp 1698431365
transform 1 0 18256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_224
timestamp 1698431365
transform 1 0 26432 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_280
timestamp 1698431365
transform 1 0 32704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_290
timestamp 1698431365
transform 1 0 33824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_312
timestamp 1698431365
transform 1 0 36288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_354
timestamp 1698431365
transform 1 0 40992 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_364
timestamp 1698431365
transform 1 0 42112 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_391
timestamp 1698431365
transform 1 0 45136 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_436
timestamp 1698431365
transform 1 0 50176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_477
timestamp 1698431365
transform 1 0 54768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_489
timestamp 1698431365
transform 1 0 56112 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_535
timestamp 1698431365
transform 1 0 61264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_4
timestamp 1698431365
transform 1 0 1792 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_74
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_95
timestamp 1698431365
transform 1 0 11984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_97
timestamp 1698431365
transform 1 0 12208 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_171
timestamp 1698431365
transform 1 0 20496 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_214
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_238
timestamp 1698431365
transform 1 0 28000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_279
timestamp 1698431365
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_288
timestamp 1698431365
transform 1 0 33600 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_368
timestamp 1698431365
transform 1 0 42560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_370
timestamp 1698431365
transform 1 0 42784 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_406
timestamp 1698431365
transform 1 0 46816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_442
timestamp 1698431365
transform 1 0 50848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_458
timestamp 1698431365
transform 1 0 52640 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_477
timestamp 1698431365
transform 1 0 54768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_481
timestamp 1698431365
transform 1 0 55216 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_515
timestamp 1698431365
transform 1 0 59024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_47
timestamp 1698431365
transform 1 0 6608 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_81
timestamp 1698431365
transform 1 0 10416 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_103
timestamp 1698431365
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_142
timestamp 1698431365
transform 1 0 17248 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_183
timestamp 1698431365
transform 1 0 21840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_255
timestamp 1698431365
transform 1 0 29904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_289
timestamp 1698431365
transform 1 0 33712 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_291
timestamp 1698431365
transform 1 0 33936 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_319
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_380
timestamp 1698431365
transform 1 0 43904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698431365
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_389
timestamp 1698431365
transform 1 0 44912 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_406
timestamp 1698431365
transform 1 0 46816 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_415
timestamp 1698431365
transform 1 0 47824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_419
timestamp 1698431365
transform 1 0 48272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_421
timestamp 1698431365
transform 1 0 48496 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_450
timestamp 1698431365
transform 1 0 51744 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_521
timestamp 1698431365
transform 1 0 59696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_543
timestamp 1698431365
transform 1 0 62160 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_17
timestamp 1698431365
transform 1 0 3248 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_80
timestamp 1698431365
transform 1 0 10304 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_111
timestamp 1698431365
transform 1 0 13776 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_194
timestamp 1698431365
transform 1 0 23072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_292
timestamp 1698431365
transform 1 0 34048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_294
timestamp 1698431365
transform 1 0 34272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_317
timestamp 1698431365
transform 1 0 36848 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_390
timestamp 1698431365
transform 1 0 45024 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_428
timestamp 1698431365
transform 1 0 49280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_432
timestamp 1698431365
transform 1 0 49728 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_434
timestamp 1698431365
transform 1 0 49952 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_441
timestamp 1698431365
transform 1 0 50736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_443
timestamp 1698431365
transform 1 0 50960 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_479
timestamp 1698431365
transform 1 0 54992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_481
timestamp 1698431365
transform 1 0 55216 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_28
timestamp 1698431365
transform 1 0 4480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_54
timestamp 1698431365
transform 1 0 7392 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_179
timestamp 1698431365
transform 1 0 21392 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_222
timestamp 1698431365
transform 1 0 26208 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_243
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_287
timestamp 1698431365
transform 1 0 33488 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_383
timestamp 1698431365
transform 1 0 44240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_408
timestamp 1698431365
transform 1 0 47040 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_453
timestamp 1698431365
transform 1 0 52080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_476
timestamp 1698431365
transform 1 0 54656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_502
timestamp 1698431365
transform 1 0 57568 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_504
timestamp 1698431365
transform 1 0 57792 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_533
timestamp 1698431365
transform 1 0 61040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_543
timestamp 1698431365
transform 1 0 62160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_4
timestamp 1698431365
transform 1 0 1792 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_64
timestamp 1698431365
transform 1 0 8512 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_98
timestamp 1698431365
transform 1 0 12320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_100
timestamp 1698431365
transform 1 0 12544 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_116
timestamp 1698431365
transform 1 0 14336 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_131
timestamp 1698431365
transform 1 0 16016 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_157
timestamp 1698431365
transform 1 0 18928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_187
timestamp 1698431365
transform 1 0 22288 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_214
timestamp 1698431365
transform 1 0 25312 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_243
timestamp 1698431365
transform 1 0 28560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_320
timestamp 1698431365
transform 1 0 37184 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_375
timestamp 1698431365
transform 1 0 43344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_379
timestamp 1698431365
transform 1 0 43792 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_489
timestamp 1698431365
transform 1 0 56112 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_514
timestamp 1698431365
transform 1 0 58912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_544
timestamp 1698431365
transform 1 0 62272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_53
timestamp 1698431365
transform 1 0 7280 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_122
timestamp 1698431365
transform 1 0 15008 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_144
timestamp 1698431365
transform 1 0 17472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_168
timestamp 1698431365
transform 1 0 20160 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_192
timestamp 1698431365
transform 1 0 22848 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_225
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_227
timestamp 1698431365
transform 1 0 26768 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_236
timestamp 1698431365
transform 1 0 27776 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_253
timestamp 1698431365
transform 1 0 29680 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_298
timestamp 1698431365
transform 1 0 34720 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_395
timestamp 1698431365
transform 1 0 45584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_399
timestamp 1698431365
transform 1 0 46032 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_454
timestamp 1698431365
transform 1 0 52192 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_459
timestamp 1698431365
transform 1 0 52752 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_543
timestamp 1698431365
transform 1 0 62160 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_48
timestamp 1698431365
transform 1 0 6720 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_96
timestamp 1698431365
transform 1 0 12096 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_158
timestamp 1698431365
transform 1 0 19040 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_160
timestamp 1698431365
transform 1 0 19264 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_191
timestamp 1698431365
transform 1 0 22736 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_269
timestamp 1698431365
transform 1 0 31472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_271
timestamp 1698431365
transform 1 0 31696 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_299
timestamp 1698431365
transform 1 0 34832 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_479
timestamp 1698431365
transform 1 0 54992 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_481
timestamp 1698431365
transform 1 0 55216 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_496
timestamp 1698431365
transform 1 0 56896 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_541
timestamp 1698431365
transform 1 0 61936 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_4
timestamp 1698431365
transform 1 0 1792 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_31
timestamp 1698431365
transform 1 0 4816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_43
timestamp 1698431365
transform 1 0 6160 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_140
timestamp 1698431365
transform 1 0 17024 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_232
timestamp 1698431365
transform 1 0 27328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_234
timestamp 1698431365
transform 1 0 27552 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_289
timestamp 1698431365
transform 1 0 33712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_291
timestamp 1698431365
transform 1 0 33936 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_360
timestamp 1698431365
transform 1 0 41664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_362
timestamp 1698431365
transform 1 0 41888 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_395
timestamp 1698431365
transform 1 0 45584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_397
timestamp 1698431365
transform 1 0 45808 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_453
timestamp 1698431365
transform 1 0 52080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_543
timestamp 1698431365
transform 1 0 62160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_4
timestamp 1698431365
transform 1 0 1792 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698431365
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_207
timestamp 1698431365
transform 1 0 24528 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_275
timestamp 1698431365
transform 1 0 32144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_277
timestamp 1698431365
transform 1 0 32368 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_296
timestamp 1698431365
transform 1 0 34496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_298
timestamp 1698431365
transform 1 0 34720 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_332
timestamp 1698431365
transform 1 0 38528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_336
timestamp 1698431365
transform 1 0 38976 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_360
timestamp 1698431365
transform 1 0 41664 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_390
timestamp 1698431365
transform 1 0 45024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_392
timestamp 1698431365
transform 1 0 45248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_406
timestamp 1698431365
transform 1 0 46816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_464
timestamp 1698431365
transform 1 0 53312 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_474
timestamp 1698431365
transform 1 0 54432 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_476
timestamp 1698431365
transform 1 0 54656 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_497
timestamp 1698431365
transform 1 0 57008 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_4
timestamp 1698431365
transform 1 0 1792 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_160
timestamp 1698431365
transform 1 0 19264 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_233
timestamp 1698431365
transform 1 0 27440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_337
timestamp 1698431365
transform 1 0 39088 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_376
timestamp 1698431365
transform 1 0 43456 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_474
timestamp 1698431365
transform 1 0 54432 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_523
timestamp 1698431365
transform 1 0 59920 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_81
timestamp 1698431365
transform 1 0 10416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_131
timestamp 1698431365
transform 1 0 16016 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_192
timestamp 1698431365
transform 1 0 22848 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_194
timestamp 1698431365
transform 1 0 23072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_239
timestamp 1698431365
transform 1 0 28112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_241
timestamp 1698431365
transform 1 0 28336 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_290
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_292
timestamp 1698431365
transform 1 0 34048 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_392
timestamp 1698431365
transform 1 0 45248 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_407
timestamp 1698431365
transform 1 0 46928 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_418
timestamp 1698431365
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_468
timestamp 1698431365
transform 1 0 53760 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_543
timestamp 1698431365
transform 1 0 62160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_32
timestamp 1698431365
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_109
timestamp 1698431365
transform 1 0 13552 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_150
timestamp 1698431365
transform 1 0 18144 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_276
timestamp 1698431365
transform 1 0 32256 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_312
timestamp 1698431365
transform 1 0 36288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698431365
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_347
timestamp 1698431365
transform 1 0 40208 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_374
timestamp 1698431365
transform 1 0 43232 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_378
timestamp 1698431365
transform 1 0 43680 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_417
timestamp 1698431365
transform 1 0 48048 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_471
timestamp 1698431365
transform 1 0 54096 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_540
timestamp 1698431365
transform 1 0 61824 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_6
timestamp 1698431365
transform 1 0 2016 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_24
timestamp 1698431365
transform 1 0 4032 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_26
timestamp 1698431365
transform 1 0 4256 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_124
timestamp 1698431365
transform 1 0 15232 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_130
timestamp 1698431365
transform 1 0 15904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_164
timestamp 1698431365
transform 1 0 19712 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_166
timestamp 1698431365
transform 1 0 19936 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_224
timestamp 1698431365
transform 1 0 26432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_275
timestamp 1698431365
transform 1 0 32144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_277
timestamp 1698431365
transform 1 0 32368 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_302
timestamp 1698431365
transform 1 0 35168 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_360
timestamp 1698431365
transform 1 0 41664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_374
timestamp 1698431365
transform 1 0 43232 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_465
timestamp 1698431365
transform 1 0 53424 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_467
timestamp 1698431365
transform 1 0 53648 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_488
timestamp 1698431365
transform 1 0 56000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_540
timestamp 1698431365
transform 1 0 61824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_544
timestamp 1698431365
transform 1 0 62272 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_68
timestamp 1698431365
transform 1 0 8960 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_109
timestamp 1698431365
transform 1 0 13552 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_118
timestamp 1698431365
transform 1 0 14560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_143
timestamp 1698431365
transform 1 0 17360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_145
timestamp 1698431365
transform 1 0 17584 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_220
timestamp 1698431365
transform 1 0 25984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_222
timestamp 1698431365
transform 1 0 26208 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_284
timestamp 1698431365
transform 1 0 33152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_341
timestamp 1698431365
transform 1 0 39536 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_343
timestamp 1698431365
transform 1 0 39760 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_359
timestamp 1698431365
transform 1 0 41552 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_402
timestamp 1698431365
transform 1 0 46368 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_454
timestamp 1698431365
transform 1 0 52192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_465
timestamp 1698431365
transform 1 0 53424 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_495
timestamp 1698431365
transform 1 0 56784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_8
timestamp 1698431365
transform 1 0 2240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_12
timestamp 1698431365
transform 1 0 2688 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_26
timestamp 1698431365
transform 1 0 4256 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_77
timestamp 1698431365
transform 1 0 9968 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_245
timestamp 1698431365
transform 1 0 28784 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_254
timestamp 1698431365
transform 1 0 29792 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_278
timestamp 1698431365
transform 1 0 32480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_332
timestamp 1698431365
transform 1 0 38528 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_334
timestamp 1698431365
transform 1 0 38752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_387
timestamp 1698431365
transform 1 0 44688 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_389
timestamp 1698431365
transform 1 0 44912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_442
timestamp 1698431365
transform 1 0 50848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_489
timestamp 1698431365
transform 1 0 56112 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_509
timestamp 1698431365
transform 1 0 58352 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_540
timestamp 1698431365
transform 1 0 61824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_544
timestamp 1698431365
transform 1 0 62272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_90
timestamp 1698431365
transform 1 0 11424 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_94
timestamp 1698431365
transform 1 0 11872 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_150
timestamp 1698431365
transform 1 0 18144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_172
timestamp 1698431365
transform 1 0 20608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_186
timestamp 1698431365
transform 1 0 22176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_224
timestamp 1698431365
transform 1 0 26432 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_226
timestamp 1698431365
transform 1 0 26656 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_281
timestamp 1698431365
transform 1 0 32816 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_380
timestamp 1698431365
transform 1 0 43904 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_408
timestamp 1698431365
transform 1 0 47040 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_437
timestamp 1698431365
transform 1 0 50288 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_439
timestamp 1698431365
transform 1 0 50512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_524
timestamp 1698431365
transform 1 0 60032 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_542
timestamp 1698431365
transform 1 0 62048 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_544
timestamp 1698431365
transform 1 0 62272 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_105
timestamp 1698431365
transform 1 0 13104 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_122
timestamp 1698431365
transform 1 0 15008 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_150
timestamp 1698431365
transform 1 0 18144 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_273
timestamp 1698431365
transform 1 0 31920 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_288
timestamp 1698431365
transform 1 0 33600 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_330
timestamp 1698431365
transform 1 0 38304 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_376
timestamp 1698431365
transform 1 0 43456 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_410
timestamp 1698431365
transform 1 0 47264 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_430
timestamp 1698431365
transform 1 0 49504 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_466
timestamp 1698431365
transform 1 0 53536 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_489
timestamp 1698431365
transform 1 0 56112 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_89
timestamp 1698431365
transform 1 0 11312 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_91
timestamp 1698431365
transform 1 0 11536 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_100
timestamp 1698431365
transform 1 0 12544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_102
timestamp 1698431365
transform 1 0 12768 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_109
timestamp 1698431365
transform 1 0 13552 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_179
timestamp 1698431365
transform 1 0 21392 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_196
timestamp 1698431365
transform 1 0 23296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_228
timestamp 1698431365
transform 1 0 26880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_230
timestamp 1698431365
transform 1 0 27104 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_251
timestamp 1698431365
transform 1 0 29456 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_255
timestamp 1698431365
transform 1 0 29904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_259
timestamp 1698431365
transform 1 0 30352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_328
timestamp 1698431365
transform 1 0 38080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_332
timestamp 1698431365
transform 1 0 38528 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1698431365
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_395
timestamp 1698431365
transform 1 0 45584 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_434
timestamp 1698431365
transform 1 0 49952 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_467
timestamp 1698431365
transform 1 0 53648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_502
timestamp 1698431365
transform 1 0 57568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_504
timestamp 1698431365
transform 1 0 57792 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_542
timestamp 1698431365
transform 1 0 62048 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_544
timestamp 1698431365
transform 1 0 62272 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_4
timestamp 1698431365
transform 1 0 1792 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_28
timestamp 1698431365
transform 1 0 4480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_152
timestamp 1698431365
transform 1 0 18368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_214
timestamp 1698431365
transform 1 0 25312 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_245
timestamp 1698431365
transform 1 0 28784 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_247
timestamp 1698431365
transform 1 0 29008 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_277
timestamp 1698431365
transform 1 0 32368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_279
timestamp 1698431365
transform 1 0 32592 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_304
timestamp 1698431365
transform 1 0 35392 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698431365
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_358
timestamp 1698431365
transform 1 0 41440 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_387
timestamp 1698431365
transform 1 0 44688 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_417
timestamp 1698431365
transform 1 0 48048 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698431365
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_460
timestamp 1698431365
transform 1 0 52864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_472
timestamp 1698431365
transform 1 0 54208 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_514
timestamp 1698431365
transform 1 0 58912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_516
timestamp 1698431365
transform 1 0 59136 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_541
timestamp 1698431365
transform 1 0 61936 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_22
timestamp 1698431365
transform 1 0 3808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_24
timestamp 1698431365
transform 1 0 4032 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_84
timestamp 1698431365
transform 1 0 10752 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_86
timestamp 1698431365
transform 1 0 10976 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_255
timestamp 1698431365
transform 1 0 29904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_261
timestamp 1698431365
transform 1 0 30576 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_311
timestamp 1698431365
transform 1 0 36176 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_352
timestamp 1698431365
transform 1 0 40768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_395
timestamp 1698431365
transform 1 0 45584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_453
timestamp 1698431365
transform 1 0 52080 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_25
timestamp 1698431365
transform 1 0 4144 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_37
timestamp 1698431365
transform 1 0 5488 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_57
timestamp 1698431365
transform 1 0 7728 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_59
timestamp 1698431365
transform 1 0 7952 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_91
timestamp 1698431365
transform 1 0 11536 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_279
timestamp 1698431365
transform 1 0 32592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_321
timestamp 1698431365
transform 1 0 37296 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_360
timestamp 1698431365
transform 1 0 41664 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_362
timestamp 1698431365
transform 1 0 41888 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_386
timestamp 1698431365
transform 1 0 44576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_422
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_442
timestamp 1698431365
transform 1 0 50848 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_489
timestamp 1698431365
transform 1 0 56112 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_533
timestamp 1698431365
transform 1 0 61040 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_39
timestamp 1698431365
transform 1 0 5712 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_90
timestamp 1698431365
transform 1 0 11424 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_128
timestamp 1698431365
transform 1 0 15680 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_190
timestamp 1698431365
transform 1 0 22624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_192
timestamp 1698431365
transform 1 0 22848 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_231
timestamp 1698431365
transform 1 0 27216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_310
timestamp 1698431365
transform 1 0 36064 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_314
timestamp 1698431365
transform 1 0 36512 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_319
timestamp 1698431365
transform 1 0 37072 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_381
timestamp 1698431365
transform 1 0 44016 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_393
timestamp 1698431365
transform 1 0 45360 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_427
timestamp 1698431365
transform 1 0 49168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_524
timestamp 1698431365
transform 1 0 60032 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_535
timestamp 1698431365
transform 1 0 61264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_58
timestamp 1698431365
transform 1 0 7840 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_100
timestamp 1698431365
transform 1 0 12544 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_207
timestamp 1698431365
transform 1 0 24528 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_209
timestamp 1698431365
transform 1 0 24752 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_216
timestamp 1698431365
transform 1 0 25536 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_239
timestamp 1698431365
transform 1 0 28112 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_273
timestamp 1698431365
transform 1 0 31920 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_277
timestamp 1698431365
transform 1 0 32368 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_336
timestamp 1698431365
transform 1 0 38976 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_370
timestamp 1698431365
transform 1 0 42784 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_496
timestamp 1698431365
transform 1 0 56896 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_515
timestamp 1698431365
transform 1 0 59024 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_544
timestamp 1698431365
transform 1 0 62272 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_14
timestamp 1698431365
transform 1 0 2912 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_21
timestamp 1698431365
transform 1 0 3696 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_45
timestamp 1698431365
transform 1 0 6384 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_98
timestamp 1698431365
transform 1 0 12320 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_109
timestamp 1698431365
transform 1 0 13552 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_174
timestamp 1698431365
transform 1 0 20832 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_233
timestamp 1698431365
transform 1 0 27440 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_249
timestamp 1698431365
transform 1 0 29232 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_314
timestamp 1698431365
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_361
timestamp 1698431365
transform 1 0 41776 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_363
timestamp 1698431365
transform 1 0 42000 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_379
timestamp 1698431365
transform 1 0 43792 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_383
timestamp 1698431365
transform 1 0 44240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_420
timestamp 1698431365
transform 1 0 48384 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_453
timestamp 1698431365
transform 1 0 52080 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_465
timestamp 1698431365
transform 1 0 53424 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_535
timestamp 1698431365
transform 1 0 61264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_6
timestamp 1698431365
transform 1 0 2016 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_20
timestamp 1698431365
transform 1 0 3584 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_24
timestamp 1698431365
transform 1 0 4032 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_30
timestamp 1698431365
transform 1 0 4704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_34
timestamp 1698431365
transform 1 0 5152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_38
timestamp 1698431365
transform 1 0 5600 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_42
timestamp 1698431365
transform 1 0 6048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_46
timestamp 1698431365
transform 1 0 6496 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_50
timestamp 1698431365
transform 1 0 6944 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_54
timestamp 1698431365
transform 1 0 7392 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_58
timestamp 1698431365
transform 1 0 7840 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_94
timestamp 1698431365
transform 1 0 11872 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_96
timestamp 1698431365
transform 1 0 12096 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_120
timestamp 1698431365
transform 1 0 14784 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_144
timestamp 1698431365
transform 1 0 17472 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_220
timestamp 1698431365
transform 1 0 25984 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_222
timestamp 1698431365
transform 1 0 26208 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_251
timestamp 1698431365
transform 1 0 29456 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_337
timestamp 1698431365
transform 1 0 39088 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_346
timestamp 1698431365
transform 1 0 40096 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_435
timestamp 1698431365
transform 1 0 50064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_452
timestamp 1698431365
transform 1 0 51968 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_524
timestamp 1698431365
transform 1 0 60032 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_528
timestamp 1698431365
transform 1 0 60480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_538
timestamp 1698431365
transform 1 0 61600 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_542
timestamp 1698431365
transform 1 0 62048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_544
timestamp 1698431365
transform 1 0 62272 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_6
timestamp 1698431365
transform 1 0 2016 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_10
timestamp 1698431365
transform 1 0 2464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_14
timestamp 1698431365
transform 1 0 2912 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_18
timestamp 1698431365
transform 1 0 3360 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_21
timestamp 1698431365
transform 1 0 3696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_25
timestamp 1698431365
transform 1 0 4144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_29
timestamp 1698431365
transform 1 0 4592 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_41
timestamp 1698431365
transform 1 0 5936 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_44
timestamp 1698431365
transform 1 0 6272 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_48
timestamp 1698431365
transform 1 0 6720 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_52
timestamp 1698431365
transform 1 0 7168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_56
timestamp 1698431365
transform 1 0 7616 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_60
timestamp 1698431365
transform 1 0 8064 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_163
timestamp 1698431365
transform 1 0 19600 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_179
timestamp 1698431365
transform 1 0 21392 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_201
timestamp 1698431365
transform 1 0 23856 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_235
timestamp 1698431365
transform 1 0 27664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_292
timestamp 1698431365
transform 1 0 34048 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_294
timestamp 1698431365
transform 1 0 34272 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_314
timestamp 1698431365
transform 1 0 36512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_339
timestamp 1698431365
transform 1 0 39312 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_341
timestamp 1698431365
transform 1 0 39536 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_358
timestamp 1698431365
transform 1 0 41440 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_362
timestamp 1698431365
transform 1 0 41888 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_400
timestamp 1698431365
transform 1 0 46144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_454
timestamp 1698431365
transform 1 0 52192 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_521
timestamp 1698431365
transform 1 0 59696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_527
timestamp 1698431365
transform 1 0 60368 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_531
timestamp 1698431365
transform 1 0 60816 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_535
timestamp 1698431365
transform 1 0 61264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_539
timestamp 1698431365
transform 1 0 61712 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_543
timestamp 1698431365
transform 1 0 62160 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_10
timestamp 1698431365
transform 1 0 2464 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_16
timestamp 1698431365
transform 1 0 3136 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_24
timestamp 1698431365
transform 1 0 4032 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_27
timestamp 1698431365
transform 1 0 4368 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_33
timestamp 1698431365
transform 1 0 5040 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_37
timestamp 1698431365
transform 1 0 5488 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_39
timestamp 1698431365
transform 1 0 5712 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_42
timestamp 1698431365
transform 1 0 6048 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_46
timestamp 1698431365
transform 1 0 6496 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_50
timestamp 1698431365
transform 1 0 6944 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_54
timestamp 1698431365
transform 1 0 7392 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_58
timestamp 1698431365
transform 1 0 7840 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_62
timestamp 1698431365
transform 1 0 8288 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_66
timestamp 1698431365
transform 1 0 8736 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_188
timestamp 1698431365
transform 1 0 22400 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_220
timestamp 1698431365
transform 1 0 25984 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_321
timestamp 1698431365
transform 1 0 37296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_323
timestamp 1698431365
transform 1 0 37520 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_345
timestamp 1698431365
transform 1 0 39984 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_349
timestamp 1698431365
transform 1 0 40432 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_376
timestamp 1698431365
transform 1 0 43456 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_418
timestamp 1698431365
transform 1 0 48160 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_422
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_455
timestamp 1698431365
transform 1 0 52304 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_525
timestamp 1698431365
transform 1 0 60144 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_529
timestamp 1698431365
transform 1 0 60592 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_533
timestamp 1698431365
transform 1 0 61040 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_537
timestamp 1698431365
transform 1 0 61488 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_541
timestamp 1698431365
transform 1 0 61936 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_45
timestamp 1698431365
transform 1 0 6384 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_51
timestamp 1698431365
transform 1 0 7056 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_55
timestamp 1698431365
transform 1 0 7504 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_59
timestamp 1698431365
transform 1 0 7952 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_63
timestamp 1698431365
transform 1 0 8400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_67
timestamp 1698431365
transform 1 0 8848 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_71
timestamp 1698431365
transform 1 0 9296 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_75
timestamp 1698431365
transform 1 0 9744 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_137
timestamp 1698431365
transform 1 0 16688 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_173
timestamp 1698431365
transform 1 0 20720 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_211
timestamp 1698431365
transform 1 0 24976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_242
timestamp 1698431365
transform 1 0 28448 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_244
timestamp 1698431365
transform 1 0 28672 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_314
timestamp 1698431365
transform 1 0 36512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_323
timestamp 1698431365
transform 1 0 37520 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_381
timestamp 1698431365
transform 1 0 44016 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_403
timestamp 1698431365
transform 1 0 46480 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_407
timestamp 1698431365
transform 1 0 46928 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_473
timestamp 1698431365
transform 1 0 54320 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_475
timestamp 1698431365
transform 1 0 54544 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_517
timestamp 1698431365
transform 1 0 59248 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_521
timestamp 1698431365
transform 1 0 59696 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_527
timestamp 1698431365
transform 1 0 60368 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_531
timestamp 1698431365
transform 1 0 60816 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_535
timestamp 1698431365
transform 1 0 61264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_539
timestamp 1698431365
transform 1 0 61712 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_543
timestamp 1698431365
transform 1 0 62160 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_34
timestamp 1698431365
transform 1 0 5152 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_50
timestamp 1698431365
transform 1 0 6944 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_54
timestamp 1698431365
transform 1 0 7392 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_58
timestamp 1698431365
transform 1 0 7840 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_62
timestamp 1698431365
transform 1 0 8288 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_78
timestamp 1698431365
transform 1 0 10080 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_82
timestamp 1698431365
transform 1 0 10528 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_86
timestamp 1698431365
transform 1 0 10976 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_119
timestamp 1698431365
transform 1 0 14672 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_138
timestamp 1698431365
transform 1 0 16800 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_231
timestamp 1698431365
transform 1 0 27216 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_358
timestamp 1698431365
transform 1 0 41440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_388
timestamp 1698431365
transform 1 0 44800 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_407
timestamp 1698431365
transform 1 0 46928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_409
timestamp 1698431365
transform 1 0 47152 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_440
timestamp 1698431365
transform 1 0 50624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_506
timestamp 1698431365
transform 1 0 58016 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_510
timestamp 1698431365
transform 1 0 58464 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_524
timestamp 1698431365
transform 1 0 60032 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_528
timestamp 1698431365
transform 1 0 60480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_532
timestamp 1698431365
transform 1 0 60928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_536
timestamp 1698431365
transform 1 0 61376 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_540
timestamp 1698431365
transform 1 0 61824 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_543
timestamp 1698431365
transform 1 0 62160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_53
timestamp 1698431365
transform 1 0 7280 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_61
timestamp 1698431365
transform 1 0 8176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_67
timestamp 1698431365
transform 1 0 8848 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_71
timestamp 1698431365
transform 1 0 9296 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_75
timestamp 1698431365
transform 1 0 9744 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_79
timestamp 1698431365
transform 1 0 10192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_83
timestamp 1698431365
transform 1 0 10640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_87
timestamp 1698431365
transform 1 0 11088 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_91
timestamp 1698431365
transform 1 0 11536 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_95
timestamp 1698431365
transform 1 0 11984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_145
timestamp 1698431365
transform 1 0 17584 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_179
timestamp 1698431365
transform 1 0 21392 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_195
timestamp 1698431365
transform 1 0 23184 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_286
timestamp 1698431365
transform 1 0 33376 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_307
timestamp 1698431365
transform 1 0 35728 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_313
timestamp 1698431365
transform 1 0 36400 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_343
timestamp 1698431365
transform 1 0 39760 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_347
timestamp 1698431365
transform 1 0 40208 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_349
timestamp 1698431365
transform 1 0 40432 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_364
timestamp 1698431365
transform 1 0 42112 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_368
timestamp 1698431365
transform 1 0 42560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_370
timestamp 1698431365
transform 1 0 42784 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_420
timestamp 1698431365
transform 1 0 48384 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_422
timestamp 1698431365
transform 1 0 48608 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_454
timestamp 1698431365
transform 1 0 52192 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_465
timestamp 1698431365
transform 1 0 53424 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_522
timestamp 1698431365
transform 1 0 59808 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_524
timestamp 1698431365
transform 1 0 60032 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_527
timestamp 1698431365
transform 1 0 60368 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_531
timestamp 1698431365
transform 1 0 60816 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_537
timestamp 1698431365
transform 1 0 61488 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_541
timestamp 1698431365
transform 1 0 61936 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_76
timestamp 1698431365
transform 1 0 9856 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_80
timestamp 1698431365
transform 1 0 10304 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_84
timestamp 1698431365
transform 1 0 10752 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_88
timestamp 1698431365
transform 1 0 11200 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_92
timestamp 1698431365
transform 1 0 11648 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_255
timestamp 1698431365
transform 1 0 29904 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_273
timestamp 1698431365
transform 1 0 31920 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_333
timestamp 1698431365
transform 1 0 38640 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_337
timestamp 1698431365
transform 1 0 39088 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_341
timestamp 1698431365
transform 1 0 39536 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_345
timestamp 1698431365
transform 1 0 39984 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_349
timestamp 1698431365
transform 1 0 40432 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_430
timestamp 1698431365
transform 1 0 49504 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_526
timestamp 1698431365
transform 1 0 60256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_530
timestamp 1698431365
transform 1 0 60704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_534
timestamp 1698431365
transform 1 0 61152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_538
timestamp 1698431365
transform 1 0 61600 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_542
timestamp 1698431365
transform 1 0 62048 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_544
timestamp 1698431365
transform 1 0 62272 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_8
timestamp 1698431365
transform 1 0 2240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_12
timestamp 1698431365
transform 1 0 2688 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_28
timestamp 1698431365
transform 1 0 4480 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_32
timestamp 1698431365
transform 1 0 4928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_69
timestamp 1698431365
transform 1 0 9072 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_79
timestamp 1698431365
transform 1 0 10192 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_83
timestamp 1698431365
transform 1 0 10640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_87
timestamp 1698431365
transform 1 0 11088 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_91
timestamp 1698431365
transform 1 0 11536 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_95
timestamp 1698431365
transform 1 0 11984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_99
timestamp 1698431365
transform 1 0 12432 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_129
timestamp 1698431365
transform 1 0 15792 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_220
timestamp 1698431365
transform 1 0 25984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_222
timestamp 1698431365
transform 1 0 26208 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_244
timestamp 1698431365
transform 1 0 28672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_310
timestamp 1698431365
transform 1 0 36064 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_314
timestamp 1698431365
transform 1 0 36512 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_323
timestamp 1698431365
transform 1 0 37520 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_357
timestamp 1698431365
transform 1 0 41328 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_363
timestamp 1698431365
transform 1 0 42000 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_377
timestamp 1698431365
transform 1 0 43568 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_381
timestamp 1698431365
transform 1 0 44016 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_406
timestamp 1698431365
transform 1 0 46816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_442
timestamp 1698431365
transform 1 0 50848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_446
timestamp 1698431365
transform 1 0 51296 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_473
timestamp 1698431365
transform 1 0 54320 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_475
timestamp 1698431365
transform 1 0 54544 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_522
timestamp 1698431365
transform 1 0 59808 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_524
timestamp 1698431365
transform 1 0 60032 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_527
timestamp 1698431365
transform 1 0 60368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_531
timestamp 1698431365
transform 1 0 60816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_535
timestamp 1698431365
transform 1 0 61264 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_543
timestamp 1698431365
transform 1 0 62160 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_66
timestamp 1698431365
transform 1 0 8736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_80
timestamp 1698431365
transform 1 0 10304 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_84
timestamp 1698431365
transform 1 0 10752 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_86
timestamp 1698431365
transform 1 0 10976 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_89
timestamp 1698431365
transform 1 0 11312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_93
timestamp 1698431365
transform 1 0 11760 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_97
timestamp 1698431365
transform 1 0 12208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_101
timestamp 1698431365
transform 1 0 12656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_105
timestamp 1698431365
transform 1 0 13104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_109
timestamp 1698431365
transform 1 0 13552 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_113
timestamp 1698431365
transform 1 0 14000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_166
timestamp 1698431365
transform 1 0 19936 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_208
timestamp 1698431365
transform 1 0 24640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_293
timestamp 1698431365
transform 1 0 34160 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_334
timestamp 1698431365
transform 1 0 38752 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_338
timestamp 1698431365
transform 1 0 39200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_342
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_348
timestamp 1698431365
transform 1 0 40320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_356
timestamp 1698431365
transform 1 0 41216 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_360
timestamp 1698431365
transform 1 0 41664 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_364
timestamp 1698431365
transform 1 0 42112 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_410
timestamp 1698431365
transform 1 0 47264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_441
timestamp 1698431365
transform 1 0 50736 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_470
timestamp 1698431365
transform 1 0 53984 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_474
timestamp 1698431365
transform 1 0 54432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_486
timestamp 1698431365
transform 1 0 55776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_515
timestamp 1698431365
transform 1 0 59024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_519
timestamp 1698431365
transform 1 0 59472 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_535
timestamp 1698431365
transform 1 0 61264 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_543
timestamp 1698431365
transform 1 0 62160 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_2
timestamp 1698431365
transform 1 0 1568 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1698431365
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_37
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_69
timestamp 1698431365
transform 1 0 9072 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_85
timestamp 1698431365
transform 1 0 10864 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_89
timestamp 1698431365
transform 1 0 11312 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_93
timestamp 1698431365
transform 1 0 11760 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_97
timestamp 1698431365
transform 1 0 12208 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_101
timestamp 1698431365
transform 1 0 12656 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_107
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_111
timestamp 1698431365
transform 1 0 13776 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_181
timestamp 1698431365
transform 1 0 21616 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_197
timestamp 1698431365
transform 1 0 23408 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_209
timestamp 1698431365
transform 1 0 24752 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_211
timestamp 1698431365
transform 1 0 24976 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_314
timestamp 1698431365
transform 1 0 36512 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_317
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_321
timestamp 1698431365
transform 1 0 37296 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_325
timestamp 1698431365
transform 1 0 37744 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_329
timestamp 1698431365
transform 1 0 38192 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_333
timestamp 1698431365
transform 1 0 38640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_337
timestamp 1698431365
transform 1 0 39088 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_343
timestamp 1698431365
transform 1 0 39760 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_373
timestamp 1698431365
transform 1 0 43120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_377
timestamp 1698431365
transform 1 0 43568 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_383
timestamp 1698431365
transform 1 0 44240 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_387
timestamp 1698431365
transform 1 0 44688 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_391
timestamp 1698431365
transform 1 0 45136 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_405
timestamp 1698431365
transform 1 0 46704 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_450
timestamp 1698431365
transform 1 0 51744 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_452
timestamp 1698431365
transform 1 0 51968 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_457
timestamp 1698431365
transform 1 0 52528 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_461
timestamp 1698431365
transform 1 0 52976 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_502
timestamp 1698431365
transform 1 0 57568 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_506
timestamp 1698431365
transform 1 0 58016 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_510
timestamp 1698431365
transform 1 0 58464 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_518
timestamp 1698431365
transform 1 0 59360 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_522
timestamp 1698431365
transform 1 0 59808 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_524
timestamp 1698431365
transform 1 0 60032 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_527
timestamp 1698431365
transform 1 0 60368 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_543
timestamp 1698431365
transform 1 0 62160 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_2
timestamp 1698431365
transform 1 0 1568 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_66
timestamp 1698431365
transform 1 0 8736 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_72
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_88
timestamp 1698431365
transform 1 0 11200 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_96
timestamp 1698431365
transform 1 0 12096 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_100
timestamp 1698431365
transform 1 0 12544 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_103
timestamp 1698431365
transform 1 0 12880 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_152
timestamp 1698431365
transform 1 0 18368 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_154
timestamp 1698431365
transform 1 0 18592 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_198
timestamp 1698431365
transform 1 0 23520 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_247
timestamp 1698431365
transform 1 0 29008 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_284
timestamp 1698431365
transform 1 0 33152 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_300
timestamp 1698431365
transform 1 0 34944 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_307
timestamp 1698431365
transform 1 0 35728 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_311
timestamp 1698431365
transform 1 0 36176 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_315
timestamp 1698431365
transform 1 0 36624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_319
timestamp 1698431365
transform 1 0 37072 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_323
timestamp 1698431365
transform 1 0 37520 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_327
timestamp 1698431365
transform 1 0 37968 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_343
timestamp 1698431365
transform 1 0 39760 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_347
timestamp 1698431365
transform 1 0 40208 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_349
timestamp 1698431365
transform 1 0 40432 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_352
timestamp 1698431365
transform 1 0 40768 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_358
timestamp 1698431365
transform 1 0 41440 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_362
timestamp 1698431365
transform 1 0 41888 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_366
timestamp 1698431365
transform 1 0 42336 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_374
timestamp 1698431365
transform 1 0 43232 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_400
timestamp 1698431365
transform 1 0 46144 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_404
timestamp 1698431365
transform 1 0 46592 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_406
timestamp 1698431365
transform 1 0 46816 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_409
timestamp 1698431365
transform 1 0 47152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_411
timestamp 1698431365
transform 1 0 47376 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_422
timestamp 1698431365
transform 1 0 48608 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_426
timestamp 1698431365
transform 1 0 49056 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_429
timestamp 1698431365
transform 1 0 49392 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_437
timestamp 1698431365
transform 1 0 50288 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_441
timestamp 1698431365
transform 1 0 50736 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_489
timestamp 1698431365
transform 1 0 56112 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_492
timestamp 1698431365
transform 1 0 56448 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_496
timestamp 1698431365
transform 1 0 56896 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_528
timestamp 1698431365
transform 1 0 60480 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_544
timestamp 1698431365
transform 1 0 62272 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_2
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698431365
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_101
timestamp 1698431365
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_137
timestamp 1698431365
transform 1 0 16688 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_139
timestamp 1698431365
transform 1 0 16912 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_174
timestamp 1698431365
transform 1 0 20832 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_310
timestamp 1698431365
transform 1 0 36064 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_314
timestamp 1698431365
transform 1 0 36512 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_321
timestamp 1698431365
transform 1 0 37296 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_337
timestamp 1698431365
transform 1 0 39088 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_345
timestamp 1698431365
transform 1 0 39984 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_349
timestamp 1698431365
transform 1 0 40432 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_353
timestamp 1698431365
transform 1 0 40880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_357
timestamp 1698431365
transform 1 0 41328 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_373
timestamp 1698431365
transform 1 0 43120 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_381
timestamp 1698431365
transform 1 0 44016 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_387
timestamp 1698431365
transform 1 0 44688 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_389
timestamp 1698431365
transform 1 0 44912 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_392
timestamp 1698431365
transform 1 0 45248 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_396
timestamp 1698431365
transform 1 0 45696 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_400
timestamp 1698431365
transform 1 0 46144 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_408
timestamp 1698431365
transform 1 0 47040 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_414
timestamp 1698431365
transform 1 0 47712 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_418
timestamp 1698431365
transform 1 0 48160 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_422
timestamp 1698431365
transform 1 0 48608 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_426
timestamp 1698431365
transform 1 0 49056 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_430
timestamp 1698431365
transform 1 0 49504 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_434
timestamp 1698431365
transform 1 0 49952 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_438
timestamp 1698431365
transform 1 0 50400 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_442
timestamp 1698431365
transform 1 0 50848 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_444
timestamp 1698431365
transform 1 0 51072 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_447
timestamp 1698431365
transform 1 0 51408 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_451
timestamp 1698431365
transform 1 0 51856 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_465
timestamp 1698431365
transform 1 0 53424 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_475
timestamp 1698431365
transform 1 0 54544 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_507
timestamp 1698431365
transform 1 0 58128 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_523
timestamp 1698431365
transform 1 0 59920 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_527
timestamp 1698431365
transform 1 0 60368 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_543
timestamp 1698431365
transform 1 0 62160 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_66
timestamp 1698431365
transform 1 0 8736 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_72
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_104
timestamp 1698431365
transform 1 0 12992 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_112
timestamp 1698431365
transform 1 0 13888 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_135
timestamp 1698431365
transform 1 0 16464 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_137
timestamp 1698431365
transform 1 0 16688 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_164
timestamp 1698431365
transform 1 0 19712 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_193
timestamp 1698431365
transform 1 0 22960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_214
timestamp 1698431365
transform 1 0 25312 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_249
timestamp 1698431365
transform 1 0 29232 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_303
timestamp 1698431365
transform 1 0 35280 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_307
timestamp 1698431365
transform 1 0 35728 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_311
timestamp 1698431365
transform 1 0 36176 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_343
timestamp 1698431365
transform 1 0 39760 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_347
timestamp 1698431365
transform 1 0 40208 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_349
timestamp 1698431365
transform 1 0 40432 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_352
timestamp 1698431365
transform 1 0 40768 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_416
timestamp 1698431365
transform 1 0 47936 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_448
timestamp 1698431365
transform 1 0 51520 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_480
timestamp 1698431365
transform 1 0 55104 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_488
timestamp 1698431365
transform 1 0 56000 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_492
timestamp 1698431365
transform 1 0 56448 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_524
timestamp 1698431365
transform 1 0 60032 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_540
timestamp 1698431365
transform 1 0 61824 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_2
timestamp 1698431365
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_36
timestamp 1698431365
transform 1 0 5376 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_70
timestamp 1698431365
transform 1 0 9184 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_104
timestamp 1698431365
transform 1 0 12992 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_164
timestamp 1698431365
transform 1 0 19712 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_172
timestamp 1698431365
transform 1 0 20608 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_198
timestamp 1698431365
transform 1 0 23520 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_206
timestamp 1698431365
transform 1 0 24416 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_208
timestamp 1698431365
transform 1 0 24640 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_237
timestamp 1698431365
transform 1 0 27888 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_246
timestamp 1698431365
transform 1 0 28896 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_269
timestamp 1698431365
transform 1 0 31472 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_271
timestamp 1698431365
transform 1 0 31696 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_294
timestamp 1698431365
transform 1 0 34272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_298
timestamp 1698431365
transform 1 0 34720 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_302
timestamp 1698431365
transform 1 0 35168 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_308
timestamp 1698431365
transform 1 0 35840 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_324
timestamp 1698431365
transform 1 0 37632 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_328
timestamp 1698431365
transform 1 0 38080 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_330
timestamp 1698431365
transform 1 0 38304 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_335
timestamp 1698431365
transform 1 0 38864 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_339
timestamp 1698431365
transform 1 0 39312 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_342
timestamp 1698431365
transform 1 0 39648 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_376
timestamp 1698431365
transform 1 0 43456 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_410
timestamp 1698431365
transform 1 0 47264 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_414
timestamp 1698431365
transform 1 0 47712 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_441
timestamp 1698431365
transform 1 0 50736 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_444
timestamp 1698431365
transform 1 0 51072 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_478
timestamp 1698431365
transform 1 0 54880 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_512
timestamp 1698431365
transform 1 0 58688 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_544
timestamp 1698431365
transform 1 0 62272 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2
timestamp 1698431365
transform -1 0 62384 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 56784 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform 1 0 32256 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform 1 0 33824 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 62384 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698431365
transform -1 0 61824 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input8
timestamp 1698431365
transform -1 0 62384 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 35168 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 62384 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 31136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 30352 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input17
timestamp 1698431365
transform -1 0 34272 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 59472 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform 1 0 59472 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform -1 0 40544 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform -1 0 4480 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform 1 0 16800 0 1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698431365
transform 1 0 26320 0 -1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698431365
transform 1 0 48608 0 -1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698431365
transform 1 0 47824 0 1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_73 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 62608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 62608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 62608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 62608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 62608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 62608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 62608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 62608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 62608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 62608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 62608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 62608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 62608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 62608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 62608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 62608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 62608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 62608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 62608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 62608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 62608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 62608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 62608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 62608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 62608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 62608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 62608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 62608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 62608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 62608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 62608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 62608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 62608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 62608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 62608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 62608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 62608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_110
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 62608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_111
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 62608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_112
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 62608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_113
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 62608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_114
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 62608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_115
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 62608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_116
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 62608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_117
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 62608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_118
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 62608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_119
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 62608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_120
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 62608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_121
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 62608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_122
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 62608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_123
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 62608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_124
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 62608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_125
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 62608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_126
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 62608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_127
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 62608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_128
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 62608 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_129
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 62608 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_130
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 62608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_131
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 62608 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_132
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 62608 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_133
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 62608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_134
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 62608 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_135
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 62608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_136
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 62608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_137
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 62608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_138
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 62608 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_139
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 62608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_140
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 62608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_141
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 62608 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_142
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 62608 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_143
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 62608 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_144
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 62608 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_145
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 62608 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  rotfpga2a_135 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  rotfpga2a_136
timestamp 1698431365
transform 1 0 61936 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  rotfpga2a_137
timestamp 1698431365
transform -1 0 38864 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_150
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_151
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_152
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_153
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_154
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_155
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_156
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_157
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_158
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_159
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_160
timestamp 1698431365
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_161
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_162
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_163
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_164
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_165
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_166
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_167
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_168
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_169
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_170
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_171
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_172
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_173
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_174
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_175
timestamp 1698431365
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_176
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_177
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_178
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_179
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_180
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_181
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_182
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_183
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_184
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_185
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_186
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_187
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_188
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_189
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_190
timestamp 1698431365
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_191
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_192
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_193
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_194
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_195
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_196
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_197
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_198
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_199
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_200
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_201
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_202
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_203
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_204
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_205
timestamp 1698431365
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_206
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_207
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_208
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_209
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_210
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_211
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_212
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_213
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_214
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_215
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_216
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_217
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_218
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_219
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_220
timestamp 1698431365
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_221
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_222
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_223
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_224
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_225
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_226
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_227
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_228
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_229
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_230
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_231
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_232
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_233
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_234
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_235
timestamp 1698431365
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_236
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_237
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_238
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_239
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_240
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_241
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_242
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_243
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_244
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_245
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_246
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_247
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_248
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_249
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_250
timestamp 1698431365
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_251
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_252
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_253
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_254
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_255
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_256
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_257
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_258
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_259
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_260
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_261
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_262
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_263
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_264
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_265
timestamp 1698431365
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_266
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_267
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_268
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_269
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_270
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_271
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_272
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_273
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_274
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_275
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_276
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_277
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_278
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_279
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_280
timestamp 1698431365
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_281
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_282
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_283
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_284
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_285
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_286
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_287
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_288
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_289
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_290
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_291
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_292
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_293
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_294
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_295
timestamp 1698431365
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_296
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_297
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_298
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_299
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_300
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_301
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_302
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_303
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_304
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_305
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_306
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_307
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_308
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_309
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_310
timestamp 1698431365
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_311
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_312
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_313
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_314
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_315
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_316
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_317
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_318
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_319
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_320
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_321
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_322
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_323
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_324
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_325
timestamp 1698431365
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_326
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_327
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_328
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_329
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_330
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_331
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_332
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_333
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_334
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_335
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_336
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_337
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_338
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_339
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_340
timestamp 1698431365
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_341
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_342
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_343
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_344
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_345
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_346
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_347
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_348
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_349
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_350
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_351
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_352
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_353
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_354
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_355
timestamp 1698431365
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_356
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_357
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_358
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_359
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_360
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_361
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_362
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_363
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_364
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_365
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_366
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_367
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_368
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_369
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_370
timestamp 1698431365
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_371
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_372
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_373
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_374
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_375
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_376
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_377
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_378
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_379
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_380
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_381
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_382
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_383
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_384
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_385
timestamp 1698431365
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_386
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_387
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_388
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_389
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_390
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_391
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_392
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_393
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_394
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_395
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_396
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_397
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_398
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_399
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_400
timestamp 1698431365
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_401
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_402
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_403
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_404
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_405
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_406
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_407
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_408
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_409
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_410
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_411
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_412
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_413
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_414
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_415
timestamp 1698431365
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_416
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_417
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_418
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_419
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_420
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_421
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_422
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_423
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_424
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_425
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_426
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_427
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_428
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_429
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_430
timestamp 1698431365
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_431
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_432
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_433
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_434
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_435
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_436
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_437
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_438
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_439
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_440
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_441
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_442
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_443
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_444
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_445
timestamp 1698431365
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_446
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_447
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_448
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_449
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_450
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_451
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_452
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_453
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_454
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_455
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_456
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_457
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_458
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_459
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_460
timestamp 1698431365
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_461
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_462
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_463
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_464
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_465
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_466
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_467
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_468
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_469
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_470
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_471
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_472
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_473
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_474
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_475
timestamp 1698431365
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_476
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_477
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_478
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_479
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_480
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_481
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_482
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_483
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_484
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_485
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_486
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_487
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_488
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_489
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_490
timestamp 1698431365
transform 1 0 60144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_491
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_492
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_493
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_494
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_495
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_496
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_497
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_498
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_499
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_500
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_501
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_502
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_503
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_504
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_505
timestamp 1698431365
transform 1 0 60144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_506
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_507
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_508
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_509
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_510
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_511
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_512
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_513
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_514
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_515
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_516
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_517
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_518
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_519
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_520
timestamp 1698431365
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_521
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_522
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_523
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_524
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_525
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_526
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_527
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_528
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_529
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_530
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_531
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_532
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_533
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_534
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_535
timestamp 1698431365
transform 1 0 60144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_536
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_537
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_538
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_539
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_540
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_541
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_542
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_543
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_544
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_545
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_546
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_547
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_548
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_549
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_550
timestamp 1698431365
transform 1 0 60144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_551
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_552
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_553
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_554
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_555
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_556
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_557
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_558
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_559
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_560
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_561
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_562
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_563
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_564
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_565
timestamp 1698431365
transform 1 0 60144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_566
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_567
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_568
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_569
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_570
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_571
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_572
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_573
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_574
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_575
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_576
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_577
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_578
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_579
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_580
timestamp 1698431365
transform 1 0 60144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_581
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_582
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_583
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_584
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_585
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_586
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_587
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_588
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_589
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_590
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_591
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_592
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_593
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_594
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_595
timestamp 1698431365
transform 1 0 60144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_596
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_597
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_598
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_599
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_600
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_601
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_602
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_603
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_604
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_605
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_606
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_607
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_608
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_609
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_610
timestamp 1698431365
transform 1 0 60144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_611
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_612
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_613
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_614
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_615
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_616
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_617
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_618
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_619
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_620
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_621
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_622
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_623
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_624
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_625
timestamp 1698431365
transform 1 0 60144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_626
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_627
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_628
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_629
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_630
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_631
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_632
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_633
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_634
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_635
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_636
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_637
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_638
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_639
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_640
timestamp 1698431365
transform 1 0 60144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_641
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_642
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_643
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_644
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_645
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_646
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_647
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_648
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_649
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_650
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_651
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_652
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_653
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_654
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_655
timestamp 1698431365
transform 1 0 60144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_656
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_657
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_658
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_659
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_660
timestamp 1698431365
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_661
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_662
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_663
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_664
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_665
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_666
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_667
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_668
timestamp 1698431365
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_669
timestamp 1698431365
transform 1 0 52304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_670
timestamp 1698431365
transform 1 0 60144 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_671
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_672
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_673
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_674
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_675
timestamp 1698431365
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_676
timestamp 1698431365
transform 1 0 48384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_677
timestamp 1698431365
transform 1 0 56224 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_678
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_679
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_680
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_681
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_682
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_683
timestamp 1698431365
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_684
timestamp 1698431365
transform 1 0 52304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_685
timestamp 1698431365
transform 1 0 60144 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_686
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_687
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_688
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_689
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_690
timestamp 1698431365
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_691
timestamp 1698431365
transform 1 0 48384 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_692
timestamp 1698431365
transform 1 0 56224 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_693
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_694
timestamp 1698431365
transform 1 0 8960 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_695
timestamp 1698431365
transform 1 0 12768 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_696
timestamp 1698431365
transform 1 0 16576 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_697
timestamp 1698431365
transform 1 0 20384 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_698
timestamp 1698431365
transform 1 0 24192 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_699
timestamp 1698431365
transform 1 0 28000 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_700
timestamp 1698431365
transform 1 0 31808 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_701
timestamp 1698431365
transform 1 0 35616 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_702
timestamp 1698431365
transform 1 0 39424 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_703
timestamp 1698431365
transform 1 0 43232 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_704
timestamp 1698431365
transform 1 0 47040 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_705
timestamp 1698431365
transform 1 0 50848 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_706
timestamp 1698431365
transform 1 0 54656 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_707
timestamp 1698431365
transform 1 0 58464 0 1 59584
box -86 -86 310 870
<< labels >>
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 54432 800 54544 0 FreeSans 448 0 0 0 in[0]
port 1 nsew signal input
flabel metal3 s 63200 29568 64000 29680 0 FreeSans 448 0 0 0 in[10]
port 2 nsew signal input
flabel metal3 s 63200 30240 64000 30352 0 FreeSans 448 0 0 0 in[11]
port 3 nsew signal input
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 in[12]
port 4 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 in[13]
port 5 nsew signal input
flabel metal3 s 63200 28896 64000 29008 0 FreeSans 448 0 0 0 in[14]
port 6 nsew signal input
flabel metal3 s 63200 27552 64000 27664 0 FreeSans 448 0 0 0 in[15]
port 7 nsew signal input
flabel metal3 s 63200 28224 64000 28336 0 FreeSans 448 0 0 0 in[16]
port 8 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 in[17]
port 9 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 in[18]
port 10 nsew signal input
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 in[1]
port 11 nsew signal input
flabel metal3 s 63200 32928 64000 33040 0 FreeSans 448 0 0 0 in[2]
port 12 nsew signal input
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 in[3]
port 13 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 in[4]
port 14 nsew signal input
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 in[5]
port 15 nsew signal input
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 in[6]
port 16 nsew signal input
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 in[7]
port 17 nsew signal input
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 in[8]
port 18 nsew signal input
flabel metal2 s 29568 63200 29680 64000 0 FreeSans 448 90 0 0 in[9]
port 19 nsew signal input
flabel metal3 s 63200 43008 64000 43120 0 FreeSans 448 0 0 0 out[0]
port 20 nsew signal tristate
flabel metal3 s 63200 58464 64000 58576 0 FreeSans 448 0 0 0 out[10]
port 21 nsew signal tristate
flabel metal2 s 38304 63200 38416 64000 0 FreeSans 448 90 0 0 out[11]
port 22 nsew signal tristate
flabel metal3 s 63200 30912 64000 31024 0 FreeSans 448 0 0 0 out[1]
port 23 nsew signal tristate
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 out[2]
port 24 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 out[3]
port 25 nsew signal tristate
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 out[4]
port 26 nsew signal tristate
flabel metal2 s 16128 63200 16240 64000 0 FreeSans 448 90 0 0 out[5]
port 27 nsew signal tristate
flabel metal2 s 26208 63200 26320 64000 0 FreeSans 448 90 0 0 out[6]
port 28 nsew signal tristate
flabel metal2 s 48384 63200 48496 64000 0 FreeSans 448 90 0 0 out[7]
port 29 nsew signal tristate
flabel metal2 s 47712 63200 47824 64000 0 FreeSans 448 90 0 0 out[8]
port 30 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 out[9]
port 31 nsew signal tristate
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 rst_n
port 32 nsew signal input
flabel metal4 s 4448 3076 4768 60428 0 FreeSans 1280 90 0 0 vdd
port 33 nsew power bidirectional
flabel metal4 s 35168 3076 35488 60428 0 FreeSans 1280 90 0 0 vdd
port 33 nsew power bidirectional
flabel metal4 s 19808 3076 20128 60428 0 FreeSans 1280 90 0 0 vss
port 34 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 60428 0 FreeSans 1280 90 0 0 vss
port 34 nsew ground bidirectional
rlabel metal1 31976 60368 31976 60368 0 vdd
rlabel metal1 31976 59584 31976 59584 0 vss
rlabel metal3 30016 55160 30016 55160 0 _0000_
rlabel metal2 33880 56336 33880 56336 0 _0001_
rlabel metal3 29792 52808 29792 52808 0 _0002_
rlabel metal2 32088 52136 32088 52136 0 _0003_
rlabel metal3 30632 54488 30632 54488 0 _0004_
rlabel metal2 29512 54768 29512 54768 0 _0005_
rlabel metal2 30408 54544 30408 54544 0 _0006_
rlabel metal2 30632 55944 30632 55944 0 _0007_
rlabel metal2 30072 56000 30072 56000 0 _0008_
rlabel metal3 31640 55384 31640 55384 0 _0009_
rlabel metal2 1288 21560 1288 21560 0 _0010_
rlabel metal2 27608 53816 27608 53816 0 _0011_
rlabel metal2 31416 55860 31416 55860 0 _0012_
rlabel metal3 2408 16184 2408 16184 0 _0013_
rlabel metal3 31080 53928 31080 53928 0 _0014_
rlabel metal3 31472 51576 31472 51576 0 _0015_
rlabel metal2 30744 50204 30744 50204 0 _0016_
rlabel metal3 29512 51352 29512 51352 0 _0017_
rlabel metal3 25984 51576 25984 51576 0 _0018_
rlabel metal3 46256 45976 46256 45976 0 _0019_
rlabel metal2 44856 50848 44856 50848 0 _0020_
rlabel metal2 45528 49392 45528 49392 0 _0021_
rlabel metal3 43400 48328 43400 48328 0 _0022_
rlabel metal2 41496 48440 41496 48440 0 _0023_
rlabel metal2 25760 39144 25760 39144 0 _0024_
rlabel metal3 32256 45864 32256 45864 0 _0025_
rlabel metal2 21672 40992 21672 40992 0 _0026_
rlabel metal2 25704 35672 25704 35672 0 _0027_
rlabel metal3 25200 19992 25200 19992 0 _0028_
rlabel metal2 10640 26824 10640 26824 0 _0029_
rlabel metal2 20272 37800 20272 37800 0 _0030_
rlabel metal2 22008 36288 22008 36288 0 _0031_
rlabel metal2 20328 38248 20328 38248 0 _0032_
rlabel metal2 39368 49280 39368 49280 0 _0033_
rlabel metal3 20440 40824 20440 40824 0 _0034_
rlabel metal2 24584 40768 24584 40768 0 _0035_
rlabel metal2 20440 39984 20440 39984 0 _0036_
rlabel metal2 17976 41888 17976 41888 0 _0037_
rlabel metal3 18648 40936 18648 40936 0 _0038_
rlabel metal2 17976 40712 17976 40712 0 _0039_
rlabel metal2 18256 41272 18256 41272 0 _0040_
rlabel metal2 24360 48720 24360 48720 0 _0041_
rlabel metal2 24248 43232 24248 43232 0 _0042_
rlabel metal2 21672 41888 21672 41888 0 _0043_
rlabel metal3 22960 41944 22960 41944 0 _0044_
rlabel metal3 22456 38696 22456 38696 0 _0045_
rlabel metal2 23688 43008 23688 43008 0 _0046_
rlabel metal4 23016 45248 23016 45248 0 _0047_
rlabel metal2 24360 40432 24360 40432 0 _0048_
rlabel metal3 23800 39480 23800 39480 0 _0049_
rlabel metal2 21784 40768 21784 40768 0 _0050_
rlabel metal2 20664 40992 20664 40992 0 _0051_
rlabel metal2 23072 41384 23072 41384 0 _0052_
rlabel metal2 26824 45024 26824 45024 0 _0053_
rlabel metal2 35672 48944 35672 48944 0 _0054_
rlabel metal3 38724 49560 38724 49560 0 _0055_
rlabel metal2 37128 49756 37128 49756 0 _0056_
rlabel metal2 34328 48608 34328 48608 0 _0057_
rlabel metal2 29736 52080 29736 52080 0 _0058_
rlabel metal2 34440 48496 34440 48496 0 _0059_
rlabel metal3 19880 48216 19880 48216 0 _0060_
rlabel metal2 21112 47992 21112 47992 0 _0061_
rlabel metal2 18984 50736 18984 50736 0 _0062_
rlabel metal2 35672 48160 35672 48160 0 _0063_
rlabel metal2 36736 51464 36736 51464 0 _0064_
rlabel metal3 35504 50568 35504 50568 0 _0065_
rlabel metal2 35448 49560 35448 49560 0 _0066_
rlabel metal2 41720 52136 41720 52136 0 _0067_
rlabel metal2 13832 46984 13832 46984 0 _0068_
rlabel metal2 16184 48048 16184 48048 0 _0069_
rlabel metal3 15932 50008 15932 50008 0 _0070_
rlabel metal3 12376 50456 12376 50456 0 _0071_
rlabel metal2 16744 23520 16744 23520 0 _0072_
rlabel metal2 16184 51240 16184 51240 0 _0073_
rlabel metal2 10696 47264 10696 47264 0 _0074_
rlabel metal3 40320 40936 40320 40936 0 _0075_
rlabel metal2 40264 44240 40264 44240 0 _0076_
rlabel metal2 40824 39984 40824 39984 0 _0077_
rlabel metal2 40488 41664 40488 41664 0 _0078_
rlabel metal4 16520 42392 16520 42392 0 _0079_
rlabel metal2 10696 45864 10696 45864 0 _0080_
rlabel metal3 14448 42728 14448 42728 0 _0081_
rlabel metal2 12712 38024 12712 38024 0 _0082_
rlabel metal3 16856 15400 16856 15400 0 _0083_
rlabel metal2 2744 41832 2744 41832 0 _0084_
rlabel metal3 16072 17248 16072 17248 0 _0085_
rlabel metal2 15736 15736 15736 15736 0 _0086_
rlabel metal2 15400 16520 15400 16520 0 _0087_
rlabel metal2 14168 33488 14168 33488 0 _0088_
rlabel metal2 10136 46144 10136 46144 0 _0089_
rlabel metal2 15736 37688 15736 37688 0 _0090_
rlabel metal3 15792 38024 15792 38024 0 _0091_
rlabel metal2 14112 37240 14112 37240 0 _0092_
rlabel metal2 11704 35672 11704 35672 0 _0093_
rlabel metal2 11368 35280 11368 35280 0 _0094_
rlabel metal2 12040 36008 12040 36008 0 _0095_
rlabel metal2 11480 36792 11480 36792 0 _0096_
rlabel metal2 16912 40376 16912 40376 0 _0097_
rlabel metal2 14728 39032 14728 39032 0 _0098_
rlabel metal3 13104 38808 13104 38808 0 _0099_
rlabel metal2 12040 39424 12040 39424 0 _0100_
rlabel metal2 9688 40656 9688 40656 0 _0101_
rlabel metal2 14728 37520 14728 37520 0 _0102_
rlabel metal2 14728 40208 14728 40208 0 _0103_
rlabel metal2 16072 37296 16072 37296 0 _0104_
rlabel metal3 13160 40936 13160 40936 0 _0105_
rlabel metal2 12992 38920 12992 38920 0 _0106_
rlabel metal2 16184 38080 16184 38080 0 _0107_
rlabel metal2 12936 40152 12936 40152 0 _0108_
rlabel metal2 12040 43064 12040 43064 0 _0109_
rlabel metal2 12264 44800 12264 44800 0 _0110_
rlabel metal2 11256 44016 11256 44016 0 _0111_
rlabel metal4 10920 45528 10920 45528 0 _0112_
rlabel metal2 9352 48608 9352 48608 0 _0113_
rlabel metal2 10584 47488 10584 47488 0 _0114_
rlabel metal2 9240 47992 9240 47992 0 _0115_
rlabel metal2 14056 46984 14056 46984 0 _0116_
rlabel metal2 9856 46088 9856 46088 0 _0117_
rlabel metal3 9688 46760 9688 46760 0 _0118_
rlabel metal2 11872 46088 11872 46088 0 _0119_
rlabel metal2 8792 46256 8792 46256 0 _0120_
rlabel metal2 9016 46032 9016 46032 0 _0121_
rlabel metal2 1624 15904 1624 15904 0 _0122_
rlabel metal2 5992 44632 5992 44632 0 _0123_
rlabel metal3 7168 42056 7168 42056 0 _0124_
rlabel metal3 22904 43400 22904 43400 0 _0125_
rlabel metal2 7336 41888 7336 41888 0 _0126_
rlabel metal3 5320 42056 5320 42056 0 _0127_
rlabel metal2 3752 41944 3752 41944 0 _0128_
rlabel metal3 15176 37520 15176 37520 0 _0129_
rlabel metal2 26264 37184 26264 37184 0 _0130_
rlabel metal2 3080 37800 3080 37800 0 _0131_
rlabel metal2 2744 37520 2744 37520 0 _0132_
rlabel metal2 4536 43400 4536 43400 0 _0133_
rlabel metal2 2632 31640 2632 31640 0 _0134_
rlabel metal2 2352 35784 2352 35784 0 _0135_
rlabel metal2 2744 29624 2744 29624 0 _0136_
rlabel metal3 9856 34888 9856 34888 0 _0137_
rlabel metal2 5880 32592 5880 32592 0 _0138_
rlabel metal3 6720 30184 6720 30184 0 _0139_
rlabel metal2 3864 31360 3864 31360 0 _0140_
rlabel metal3 4760 20664 4760 20664 0 _0141_
rlabel metal3 6776 26376 6776 26376 0 _0142_
rlabel metal2 6216 24584 6216 24584 0 _0143_
rlabel metal2 3192 23072 3192 23072 0 _0144_
rlabel metal2 2912 24472 2912 24472 0 _0145_
rlabel metal2 3304 36960 3304 36960 0 _0146_
rlabel metal3 4928 38920 4928 38920 0 _0147_
rlabel metal2 3080 35280 3080 35280 0 _0148_
rlabel metal2 3192 31528 3192 31528 0 _0149_
rlabel metal2 5656 28560 5656 28560 0 _0150_
rlabel metal2 5992 29792 5992 29792 0 _0151_
rlabel metal2 3976 36400 3976 36400 0 _0152_
rlabel metal2 2520 31920 2520 31920 0 _0153_
rlabel metal2 6216 32256 6216 32256 0 _0154_
rlabel metal2 2408 32480 2408 32480 0 _0155_
rlabel metal2 2744 32760 2744 32760 0 _0156_
rlabel metal2 6216 31696 6216 31696 0 _0157_
rlabel metal2 2072 34832 2072 34832 0 _0158_
rlabel metal2 2184 36400 2184 36400 0 _0159_
rlabel metal2 3192 42448 3192 42448 0 _0160_
rlabel metal2 4256 42952 4256 42952 0 _0161_
rlabel metal2 3192 42840 3192 42840 0 _0162_
rlabel metal2 2632 44688 2632 44688 0 _0163_
rlabel metal2 8568 44800 8568 44800 0 _0164_
rlabel metal3 5208 44408 5208 44408 0 _0165_
rlabel metal2 2856 43008 2856 43008 0 _0166_
rlabel metal2 22904 44912 22904 44912 0 _0167_
rlabel metal2 3416 45752 3416 45752 0 _0168_
rlabel metal2 3304 45248 3304 45248 0 _0169_
rlabel metal2 1568 49784 1568 49784 0 _0170_
rlabel metal3 21728 56728 21728 56728 0 _0171_
rlabel metal3 18312 53592 18312 53592 0 _0172_
rlabel metal2 16408 28896 16408 28896 0 _0173_
rlabel metal3 2128 18424 2128 18424 0 _0174_
rlabel metal2 16576 31752 16576 31752 0 _0175_
rlabel metal3 16744 26264 16744 26264 0 _0176_
rlabel metal2 19432 24136 19432 24136 0 _0177_
rlabel metal2 16968 26992 16968 26992 0 _0178_
rlabel metal2 15848 27496 15848 27496 0 _0179_
rlabel metal2 14896 26488 14896 26488 0 _0180_
rlabel metal3 17080 57064 17080 57064 0 _0181_
rlabel metal2 2296 18256 2296 18256 0 _0182_
rlabel metal2 13720 30688 13720 30688 0 _0183_
rlabel metal3 16296 30968 16296 30968 0 _0184_
rlabel metal2 18760 31416 18760 31416 0 _0185_
rlabel metal2 17528 32032 17528 32032 0 _0186_
rlabel metal2 16408 31528 16408 31528 0 _0187_
rlabel metal2 5432 21840 5432 21840 0 _0188_
rlabel metal2 4648 22120 4648 22120 0 _0189_
rlabel metal2 4872 23128 4872 23128 0 _0190_
rlabel metal2 4648 23352 4648 23352 0 _0191_
rlabel metal3 3080 17808 3080 17808 0 _0192_
rlabel metal2 15512 32480 15512 32480 0 _0193_
rlabel metal2 14560 32312 14560 32312 0 _0194_
rlabel metal2 11256 30520 11256 30520 0 _0195_
rlabel metal3 13160 31192 13160 31192 0 _0196_
rlabel metal2 4424 17360 4424 17360 0 _0197_
rlabel metal2 2072 18760 2072 18760 0 _0198_
rlabel metal2 15624 29456 15624 29456 0 _0199_
rlabel metal2 15288 31136 15288 31136 0 _0200_
rlabel metal2 19320 32928 19320 32928 0 _0201_
rlabel metal2 17416 32760 17416 32760 0 _0202_
rlabel metal3 16240 31080 16240 31080 0 _0203_
rlabel metal2 17752 33824 17752 33824 0 _0204_
rlabel metal3 15568 41272 15568 41272 0 _0205_
rlabel metal2 15512 53424 15512 53424 0 _0206_
rlabel metal2 16240 53704 16240 53704 0 _0207_
rlabel metal3 15288 53480 15288 53480 0 _0208_
rlabel metal2 16184 56000 16184 56000 0 _0209_
rlabel metal2 2408 33600 2408 33600 0 _0210_
rlabel metal2 8568 31248 8568 31248 0 _0211_
rlabel metal2 2856 33040 2856 33040 0 _0212_
rlabel metal3 2184 31136 2184 31136 0 _0213_
rlabel metal2 1512 51940 1512 51940 0 _0214_
rlabel metal3 20104 56840 20104 56840 0 _0215_
rlabel metal2 15512 50960 15512 50960 0 _0216_
rlabel metal2 20216 54992 20216 54992 0 _0217_
rlabel metal2 18984 55608 18984 55608 0 _0218_
rlabel metal3 18872 54376 18872 54376 0 _0219_
rlabel metal2 17528 54208 17528 54208 0 _0220_
rlabel metal2 15456 52920 15456 52920 0 _0221_
rlabel metal2 15848 53200 15848 53200 0 _0222_
rlabel metal3 14168 53032 14168 53032 0 _0223_
rlabel metal2 14392 56504 14392 56504 0 _0224_
rlabel metal2 17528 52080 17528 52080 0 _0225_
rlabel metal2 17416 51688 17416 51688 0 _0226_
rlabel metal2 17584 51128 17584 51128 0 _0227_
rlabel metal2 21168 52136 21168 52136 0 _0228_
rlabel metal3 31976 48216 31976 48216 0 _0229_
rlabel metal2 28952 46928 28952 46928 0 _0230_
rlabel metal2 30520 28672 30520 28672 0 _0231_
rlabel metal2 28280 42280 28280 42280 0 _0232_
rlabel metal2 26152 29512 26152 29512 0 _0233_
rlabel metal2 32984 27440 32984 27440 0 _0234_
rlabel metal2 34216 23576 34216 23576 0 _0235_
rlabel metal2 33096 28392 33096 28392 0 _0236_
rlabel metal3 32704 27832 32704 27832 0 _0237_
rlabel metal2 33208 28504 33208 28504 0 _0238_
rlabel metal2 28616 46368 28616 46368 0 _0239_
rlabel metal3 29288 42616 29288 42616 0 _0240_
rlabel metal2 28728 29344 28728 29344 0 _0241_
rlabel metal2 17976 25648 17976 25648 0 _0242_
rlabel metal2 18648 27888 18648 27888 0 _0243_
rlabel metal3 20440 28840 20440 28840 0 _0244_
rlabel metal2 18984 29400 18984 29400 0 _0245_
rlabel metal2 20216 32424 20216 32424 0 _0246_
rlabel metal2 19544 31136 19544 31136 0 _0247_
rlabel metal3 20048 29400 20048 29400 0 _0248_
rlabel metal2 26208 30856 26208 30856 0 _0249_
rlabel metal2 26040 30856 26040 30856 0 _0250_
rlabel metal2 26376 29680 26376 29680 0 _0251_
rlabel metal2 23240 19488 23240 19488 0 _0252_
rlabel metal3 52528 8344 52528 8344 0 _0253_
rlabel metal2 29960 29456 29960 29456 0 _0254_
rlabel metal2 23912 30688 23912 30688 0 _0255_
rlabel metal2 21840 29176 21840 29176 0 _0256_
rlabel metal2 25592 29904 25592 29904 0 _0257_
rlabel metal2 24696 29848 24696 29848 0 _0258_
rlabel metal3 28000 42504 28000 42504 0 _0259_
rlabel metal2 26600 45472 26600 45472 0 _0260_
rlabel metal2 27048 44800 27048 44800 0 _0261_
rlabel metal2 26712 45584 26712 45584 0 _0262_
rlabel metal2 24136 46088 24136 46088 0 _0263_
rlabel metal2 18872 53760 18872 53760 0 _0264_
rlabel metal2 22120 46872 22120 46872 0 _0265_
rlabel metal2 24136 42448 24136 42448 0 _0266_
rlabel metal2 15288 41272 15288 41272 0 _0267_
rlabel metal3 23016 44296 23016 44296 0 _0268_
rlabel metal3 23184 44408 23184 44408 0 _0269_
rlabel metal2 23912 44408 23912 44408 0 _0270_
rlabel metal2 24640 45640 24640 45640 0 _0271_
rlabel metal2 23240 45360 23240 45360 0 _0272_
rlabel metal3 23744 45080 23744 45080 0 _0273_
rlabel metal4 15176 42504 15176 42504 0 _0274_
rlabel metal2 15624 44352 15624 44352 0 _0275_
rlabel metal3 20832 21560 20832 21560 0 _0276_
rlabel metal2 19656 24584 19656 24584 0 _0277_
rlabel metal2 21784 41720 21784 41720 0 _0278_
rlabel metal2 18312 42168 18312 42168 0 _0279_
rlabel metal2 18592 39032 18592 39032 0 _0280_
rlabel metal3 20216 38808 20216 38808 0 _0281_
rlabel via2 17752 45864 17752 45864 0 _0282_
rlabel metal2 17640 43120 17640 43120 0 _0283_
rlabel metal3 21280 18424 21280 18424 0 _0284_
rlabel metal3 1904 39480 1904 39480 0 _0285_
rlabel metal3 19656 18424 19656 18424 0 _0286_
rlabel metal3 20832 16072 20832 16072 0 _0287_
rlabel metal3 20160 16744 20160 16744 0 _0288_
rlabel metal3 19208 16968 19208 16968 0 _0289_
rlabel metal2 18312 17920 18312 17920 0 _0290_
rlabel metal2 18984 44016 18984 44016 0 _0291_
rlabel metal3 19152 21784 19152 21784 0 _0292_
rlabel metal2 20104 19656 20104 19656 0 _0293_
rlabel metal2 12600 20720 12600 20720 0 _0294_
rlabel metal3 12320 22120 12320 22120 0 _0295_
rlabel metal4 12376 20720 12376 20720 0 _0296_
rlabel metal2 13160 20664 13160 20664 0 _0297_
rlabel metal2 12712 22064 12712 22064 0 _0298_
rlabel metal2 17024 26488 17024 26488 0 _0299_
rlabel metal2 17864 21616 17864 21616 0 _0300_
rlabel metal2 16520 20272 16520 20272 0 _0301_
rlabel metal3 18648 19992 18648 19992 0 _0302_
rlabel metal2 15512 17528 15512 17528 0 _0303_
rlabel metal3 16352 17864 16352 17864 0 _0304_
rlabel metal2 18088 21392 18088 21392 0 _0305_
rlabel metal2 23184 3192 23184 3192 0 _0306_
rlabel metal2 19880 18256 19880 18256 0 _0307_
rlabel metal2 16072 18368 16072 18368 0 _0308_
rlabel metal2 16632 20216 16632 20216 0 _0309_
rlabel metal2 17304 20832 17304 20832 0 _0310_
rlabel metal2 17416 21280 17416 21280 0 _0311_
rlabel metal2 17976 36008 17976 36008 0 _0312_
rlabel metal2 17136 41048 17136 41048 0 _0313_
rlabel metal2 16184 42392 16184 42392 0 _0314_
rlabel metal2 16912 40936 16912 40936 0 _0315_
rlabel metal3 17136 39480 17136 39480 0 _0316_
rlabel metal2 24920 42336 24920 42336 0 _0317_
rlabel metal2 15344 41944 15344 41944 0 _0318_
rlabel metal2 14168 40264 14168 40264 0 _0319_
rlabel metal3 10528 39592 10528 39592 0 _0320_
rlabel metal2 13832 40320 13832 40320 0 _0321_
rlabel metal2 14392 40992 14392 40992 0 _0322_
rlabel metal2 15960 40320 15960 40320 0 _0323_
rlabel metal3 16464 40936 16464 40936 0 _0324_
rlabel metal3 16352 41944 16352 41944 0 _0325_
rlabel metal2 15400 42448 15400 42448 0 _0326_
rlabel metal2 14728 42336 14728 42336 0 _0327_
rlabel metal2 15512 40376 15512 40376 0 _0328_
rlabel metal2 15736 39508 15736 39508 0 _0329_
rlabel metal2 18312 36064 18312 36064 0 _0330_
rlabel metal2 15624 35280 15624 35280 0 _0331_
rlabel metal3 7728 34888 7728 34888 0 _0332_
rlabel metal2 7896 20384 7896 20384 0 _0333_
rlabel metal2 11200 16072 11200 16072 0 _0334_
rlabel metal2 10808 15204 10808 15204 0 _0335_
rlabel metal2 10584 8288 10584 8288 0 _0336_
rlabel metal2 9744 15960 9744 15960 0 _0337_
rlabel metal2 8008 16520 8008 16520 0 _0338_
rlabel metal3 9128 38024 9128 38024 0 _0339_
rlabel metal2 11256 21056 11256 21056 0 _0340_
rlabel metal2 9912 16632 9912 16632 0 _0341_
rlabel metal2 9688 18424 9688 18424 0 _0342_
rlabel metal2 4424 21616 4424 21616 0 _0343_
rlabel metal2 6328 21056 6328 21056 0 _0344_
rlabel metal3 11032 19208 11032 19208 0 _0345_
rlabel metal2 8568 20384 8568 20384 0 _0346_
rlabel metal2 6664 22344 6664 22344 0 _0347_
rlabel metal2 7336 19880 7336 19880 0 _0348_
rlabel metal2 5544 16632 5544 16632 0 _0349_
rlabel metal3 8008 17080 8008 17080 0 _0350_
rlabel metal2 7448 17976 7448 17976 0 _0351_
rlabel metal2 9576 19096 9576 19096 0 _0352_
rlabel metal3 9800 20664 9800 20664 0 _0353_
rlabel metal3 9912 22232 9912 22232 0 _0354_
rlabel metal2 6104 20776 6104 20776 0 _0355_
rlabel metal2 6328 19880 6328 19880 0 _0356_
rlabel metal2 9016 20608 9016 20608 0 _0357_
rlabel metal2 8120 22568 8120 22568 0 _0358_
rlabel metal2 10584 22456 10584 22456 0 _0359_
rlabel metal2 8344 31472 8344 31472 0 _0360_
rlabel metal2 9016 41104 9016 41104 0 _0361_
rlabel metal3 7000 40600 7000 40600 0 _0362_
rlabel metal2 10248 32256 10248 32256 0 _0363_
rlabel metal2 8568 32816 8568 32816 0 _0364_
rlabel metal2 12152 40656 12152 40656 0 _0365_
rlabel metal2 7560 34944 7560 34944 0 _0366_
rlabel metal2 2184 34328 2184 34328 0 _0367_
rlabel metal3 8848 33432 8848 33432 0 _0368_
rlabel metal2 9240 32536 9240 32536 0 _0369_
rlabel metal3 9520 33320 9520 33320 0 _0370_
rlabel metal2 8120 31192 8120 31192 0 _0371_
rlabel metal2 8288 30968 8288 30968 0 _0372_
rlabel metal2 2968 31696 2968 31696 0 _0373_
rlabel metal2 6440 31640 6440 31640 0 _0374_
rlabel metal2 7448 31584 7448 31584 0 _0375_
rlabel metal2 16296 32592 16296 32592 0 _0376_
rlabel metal2 16016 29624 16016 29624 0 _0377_
rlabel metal2 15736 30184 15736 30184 0 _0378_
rlabel metal2 16184 29400 16184 29400 0 _0379_
rlabel metal3 16128 25480 16128 25480 0 _0380_
rlabel metal2 16968 29512 16968 29512 0 _0381_
rlabel metal2 14056 34272 14056 34272 0 _0382_
rlabel metal3 12264 30184 12264 30184 0 _0383_
rlabel metal3 17360 34888 17360 34888 0 _0384_
rlabel metal2 12880 34328 12880 34328 0 _0385_
rlabel metal2 22568 33376 22568 33376 0 _0386_
rlabel metal2 23128 55552 23128 55552 0 _0387_
rlabel metal2 23800 32200 23800 32200 0 _0388_
rlabel metal3 29624 34216 29624 34216 0 _0389_
rlabel metal2 24360 27384 24360 27384 0 _0390_
rlabel metal2 24584 25424 24584 25424 0 _0391_
rlabel metal2 44184 28616 44184 28616 0 _0392_
rlabel metal2 47152 26712 47152 26712 0 _0393_
rlabel metal2 23912 18200 23912 18200 0 _0394_
rlabel metal2 44744 28392 44744 28392 0 _0395_
rlabel metal2 30520 25312 30520 25312 0 _0396_
rlabel metal2 27048 33208 27048 33208 0 _0397_
rlabel metal2 27664 27272 27664 27272 0 _0398_
rlabel metal2 26152 26152 26152 26152 0 _0399_
rlabel metal2 27048 24696 27048 24696 0 _0400_
rlabel metal2 30072 23016 30072 23016 0 _0401_
rlabel metal3 32872 23688 32872 23688 0 _0402_
rlabel metal2 30408 23408 30408 23408 0 _0403_
rlabel metal2 28280 21392 28280 21392 0 _0404_
rlabel metal2 21280 20888 21280 20888 0 _0405_
rlabel metal2 20776 23856 20776 23856 0 _0406_
rlabel metal3 22792 24024 22792 24024 0 _0407_
rlabel metal2 25256 22400 25256 22400 0 _0408_
rlabel metal3 25480 22344 25480 22344 0 _0409_
rlabel metal2 27608 24920 27608 24920 0 _0410_
rlabel metal2 24248 25984 24248 25984 0 _0411_
rlabel metal2 22568 25872 22568 25872 0 _0412_
rlabel metal3 25368 27944 25368 27944 0 _0413_
rlabel metal2 25928 26152 25928 26152 0 _0414_
rlabel metal2 25928 24864 25928 24864 0 _0415_
rlabel metal2 29400 22904 29400 22904 0 _0416_
rlabel metal2 25816 26040 25816 26040 0 _0417_
rlabel metal2 25480 23184 25480 23184 0 _0418_
rlabel metal2 25480 27720 25480 27720 0 _0419_
rlabel metal2 24696 32648 24696 32648 0 _0420_
rlabel metal3 25284 33880 25284 33880 0 _0421_
rlabel metal2 23128 29848 23128 29848 0 _0422_
rlabel metal2 25816 30296 25816 30296 0 _0423_
rlabel metal2 23240 30856 23240 30856 0 _0424_
rlabel metal3 23072 30856 23072 30856 0 _0425_
rlabel metal2 22568 31416 22568 31416 0 _0426_
rlabel metal2 16968 34048 16968 34048 0 _0427_
rlabel metal3 20496 33208 20496 33208 0 _0428_
rlabel metal2 22008 33656 22008 33656 0 _0429_
rlabel metal2 25424 33544 25424 33544 0 _0430_
rlabel metal2 24360 31808 24360 31808 0 _0431_
rlabel metal2 62552 21336 62552 21336 0 _0432_
rlabel metal3 23408 31752 23408 31752 0 _0433_
rlabel metal3 22232 22232 22232 22232 0 _0434_
rlabel metal2 23352 22904 23352 22904 0 _0435_
rlabel metal2 22344 23576 22344 23576 0 _0436_
rlabel metal2 23296 27832 23296 27832 0 _0437_
rlabel metal2 22960 37912 22960 37912 0 _0438_
rlabel metal2 2744 15736 2744 15736 0 _0439_
rlabel metal2 33544 19936 33544 19936 0 _0440_
rlabel metal3 24528 19096 24528 19096 0 _0441_
rlabel metal2 25592 18312 25592 18312 0 _0442_
rlabel metal2 37688 18816 37688 18816 0 _0443_
rlabel metal4 54040 13720 54040 13720 0 _0444_
rlabel metal2 44856 18760 44856 18760 0 _0445_
rlabel metal2 39144 19600 39144 19600 0 _0446_
rlabel metal2 36120 17920 36120 17920 0 _0447_
rlabel metal2 35672 17752 35672 17752 0 _0448_
rlabel metal2 23856 34888 23856 34888 0 _0449_
rlabel metal2 24976 26376 24976 26376 0 _0450_
rlabel metal2 28728 19040 28728 19040 0 _0451_
rlabel metal2 26600 14168 26600 14168 0 _0452_
rlabel metal2 23464 12768 23464 12768 0 _0453_
rlabel metal2 26152 14448 26152 14448 0 _0454_
rlabel metal2 26152 15960 26152 15960 0 _0455_
rlabel metal2 26712 16576 26712 16576 0 _0456_
rlabel metal2 33992 22064 33992 22064 0 _0457_
rlabel metal2 28504 18144 28504 18144 0 _0458_
rlabel metal3 26348 16968 26348 16968 0 _0459_
rlabel metal2 27608 16744 27608 16744 0 _0460_
rlabel metal2 29176 16744 29176 16744 0 _0461_
rlabel metal2 29512 17248 29512 17248 0 _0462_
rlabel metal3 25200 19880 25200 19880 0 _0463_
rlabel metal2 26712 19040 26712 19040 0 _0464_
rlabel metal2 26600 20048 26600 20048 0 _0465_
rlabel metal2 26768 17640 26768 17640 0 _0466_
rlabel metal2 26376 17416 26376 17416 0 _0467_
rlabel metal2 25704 19320 25704 19320 0 _0468_
rlabel metal2 25928 20328 25928 20328 0 _0469_
rlabel metal2 3248 16184 3248 16184 0 _0470_
rlabel metal2 13048 24976 13048 24976 0 _0471_
rlabel metal3 15120 24696 15120 24696 0 _0472_
rlabel metal2 14056 23632 14056 23632 0 _0473_
rlabel metal2 22232 29680 22232 29680 0 _0474_
rlabel metal2 22848 28056 22848 28056 0 _0475_
rlabel metal3 16296 19208 16296 19208 0 _0476_
rlabel metal3 16044 19320 16044 19320 0 _0477_
rlabel metal2 14560 22344 14560 22344 0 _0478_
rlabel metal2 13720 24528 13720 24528 0 _0479_
rlabel metal2 16520 24080 16520 24080 0 _0480_
rlabel metal2 2296 16464 2296 16464 0 _0481_
rlabel metal3 12376 24136 12376 24136 0 _0482_
rlabel metal2 12544 24136 12544 24136 0 _0483_
rlabel metal2 11592 23800 11592 23800 0 _0484_
rlabel metal3 23576 16968 23576 16968 0 _0485_
rlabel metal2 15512 20720 15512 20720 0 _0486_
rlabel metal2 15680 20888 15680 20888 0 _0487_
rlabel metal2 16184 22736 16184 22736 0 _0488_
rlabel metal3 18368 20776 18368 20776 0 _0489_
rlabel metal2 20104 21112 20104 21112 0 _0490_
rlabel metal3 11368 16072 11368 16072 0 _0491_
rlabel metal2 12824 41272 12824 41272 0 _0492_
rlabel metal3 14056 25256 14056 25256 0 _0493_
rlabel metal2 14112 15736 14112 15736 0 _0494_
rlabel metal2 16520 11312 16520 11312 0 _0495_
rlabel metal3 18312 5880 18312 5880 0 _0496_
rlabel metal2 42392 7952 42392 7952 0 _0497_
rlabel metal2 22904 7504 22904 7504 0 _0498_
rlabel metal2 50792 5488 50792 5488 0 _0499_
rlabel metal2 23688 8288 23688 8288 0 _0500_
rlabel metal3 22960 8904 22960 8904 0 _0501_
rlabel metal2 17976 14224 17976 14224 0 _0502_
rlabel metal2 21784 11536 21784 11536 0 _0503_
rlabel metal2 21672 9352 21672 9352 0 _0504_
rlabel metal2 20440 9800 20440 9800 0 _0505_
rlabel metal2 15960 9296 15960 9296 0 _0506_
rlabel metal2 16408 8680 16408 8680 0 _0507_
rlabel metal2 15736 9072 15736 9072 0 _0508_
rlabel metal2 16128 9912 16128 9912 0 _0509_
rlabel metal3 24528 14504 24528 14504 0 _0510_
rlabel metal2 18424 13328 18424 13328 0 _0511_
rlabel metal2 19320 9016 19320 9016 0 _0512_
rlabel metal2 18704 10360 18704 10360 0 _0513_
rlabel metal2 16632 9352 16632 9352 0 _0514_
rlabel metal2 16968 7840 16968 7840 0 _0515_
rlabel metal2 17808 11480 17808 11480 0 _0516_
rlabel metal3 20720 7560 20720 7560 0 _0517_
rlabel metal2 17864 11928 17864 11928 0 _0518_
rlabel metal2 18200 9072 18200 9072 0 _0519_
rlabel metal2 20104 7168 20104 7168 0 _0520_
rlabel metal2 19768 9800 19768 9800 0 _0521_
rlabel metal2 16856 12712 16856 12712 0 _0522_
rlabel metal2 14056 14896 14056 14896 0 _0523_
rlabel metal2 13944 15568 13944 15568 0 _0524_
rlabel metal3 7784 20552 7784 20552 0 _0525_
rlabel metal3 8456 19208 8456 19208 0 _0526_
rlabel metal2 8624 19992 8624 19992 0 _0527_
rlabel metal2 12264 18088 12264 18088 0 _0528_
rlabel metal2 14056 21112 14056 21112 0 _0529_
rlabel metal2 12152 17696 12152 17696 0 _0530_
rlabel metal3 12208 16296 12208 16296 0 _0531_
rlabel metal3 42728 25704 42728 25704 0 _0532_
rlabel metal3 16408 13832 16408 13832 0 _0533_
rlabel metal2 12936 15680 12936 15680 0 _0534_
rlabel metal2 12600 15624 12600 15624 0 _0535_
rlabel metal2 8344 21168 8344 21168 0 _0536_
rlabel metal2 5544 20496 5544 20496 0 _0537_
rlabel metal2 8456 19152 8456 19152 0 _0538_
rlabel metal2 5768 19656 5768 19656 0 _0539_
rlabel metal2 1960 20328 1960 20328 0 _0540_
rlabel metal2 1848 21280 1848 21280 0 _0541_
rlabel metal2 3304 32256 3304 32256 0 _0542_
rlabel metal2 7000 26992 7000 26992 0 _0543_
rlabel metal2 9072 16072 9072 16072 0 _0544_
rlabel metal3 6440 15400 6440 15400 0 _0545_
rlabel metal2 8232 12824 8232 12824 0 _0546_
rlabel metal2 14504 9688 14504 9688 0 _0547_
rlabel metal2 15176 9912 15176 9912 0 _0548_
rlabel metal2 8904 11088 8904 11088 0 _0549_
rlabel metal2 7840 12040 7840 12040 0 _0550_
rlabel metal2 25928 11032 25928 11032 0 _0551_
rlabel metal3 27496 6664 27496 6664 0 _0552_
rlabel metal2 27048 10640 27048 10640 0 _0553_
rlabel metal3 25032 9240 25032 9240 0 _0554_
rlabel metal3 16632 9800 16632 9800 0 _0555_
rlabel metal3 5600 25256 5600 25256 0 _0556_
rlabel metal2 4648 16016 4648 16016 0 _0557_
rlabel metal3 5432 15848 5432 15848 0 _0558_
rlabel metal2 7560 12992 7560 12992 0 _0559_
rlabel metal2 5992 10808 5992 10808 0 _0560_
rlabel metal2 6328 11480 6328 11480 0 _0561_
rlabel metal2 2520 12376 2520 12376 0 _0562_
rlabel metal2 10472 11312 10472 11312 0 _0563_
rlabel metal2 7448 11032 7448 11032 0 _0564_
rlabel metal2 8680 12992 8680 12992 0 _0565_
rlabel metal2 6608 16184 6608 16184 0 _0566_
rlabel metal2 8008 11704 8008 11704 0 _0567_
rlabel metal3 7168 14280 7168 14280 0 _0568_
rlabel metal2 5320 15344 5320 15344 0 _0569_
rlabel metal2 6776 21728 6776 21728 0 _0570_
rlabel metal2 7336 26600 7336 26600 0 _0571_
rlabel metal2 6328 25144 6328 25144 0 _0572_
rlabel metal3 8176 26264 8176 26264 0 _0573_
rlabel metal2 9240 21672 9240 21672 0 _0574_
rlabel metal3 8176 24472 8176 24472 0 _0575_
rlabel metal2 6552 24528 6552 24528 0 _0576_
rlabel metal2 7896 25424 7896 25424 0 _0577_
rlabel metal2 7000 24080 7000 24080 0 _0578_
rlabel metal2 8456 25032 8456 25032 0 _0579_
rlabel metal2 16296 28280 16296 28280 0 _0580_
rlabel metal2 18536 25536 18536 25536 0 _0581_
rlabel metal2 41496 27832 41496 27832 0 _0582_
rlabel metal3 40152 29960 40152 29960 0 _0583_
rlabel metal2 41384 25536 41384 25536 0 _0584_
rlabel metal2 47208 41552 47208 41552 0 _0585_
rlabel metal2 41384 28560 41384 28560 0 _0586_
rlabel metal2 40040 28000 40040 28000 0 _0587_
rlabel metal2 16184 25984 16184 25984 0 _0588_
rlabel metal2 40152 26600 40152 26600 0 _0589_
rlabel metal2 39368 25088 39368 25088 0 _0590_
rlabel metal3 45192 21784 45192 21784 0 _0591_
rlabel metal2 44184 21504 44184 21504 0 _0592_
rlabel metal3 45752 24696 45752 24696 0 _0593_
rlabel metal2 43288 22456 43288 22456 0 _0594_
rlabel metal3 44408 22456 44408 22456 0 _0595_
rlabel metal2 31752 5600 31752 5600 0 _0596_
rlabel metal2 33992 5656 33992 5656 0 _0597_
rlabel metal2 33096 5824 33096 5824 0 _0598_
rlabel metal2 30744 5376 30744 5376 0 _0599_
rlabel metal2 40432 23128 40432 23128 0 _0600_
rlabel metal2 41832 23296 41832 23296 0 _0601_
rlabel metal3 40936 25480 40936 25480 0 _0602_
rlabel metal2 11816 15400 11816 15400 0 _0603_
rlabel metal2 38360 25200 38360 25200 0 _0604_
rlabel metal3 40152 27160 40152 27160 0 _0605_
rlabel metal2 40264 27888 40264 27888 0 _0606_
rlabel metal2 40824 21448 40824 21448 0 _0607_
rlabel metal2 40040 23072 40040 23072 0 _0608_
rlabel metal2 40264 25536 40264 25536 0 _0609_
rlabel metal2 39200 24136 39200 24136 0 _0610_
rlabel metal2 37968 27720 37968 27720 0 _0611_
rlabel metal2 18312 25424 18312 25424 0 _0612_
rlabel metal2 18088 24976 18088 24976 0 _0613_
rlabel metal2 17640 23968 17640 23968 0 _0614_
rlabel metal2 21448 23576 21448 23576 0 _0615_
rlabel metal2 10248 13048 10248 13048 0 _0616_
rlabel metal2 6104 12936 6104 12936 0 _0617_
rlabel metal3 8344 12040 8344 12040 0 _0618_
rlabel metal2 8344 8960 8344 8960 0 _0619_
rlabel metal2 2856 17360 2856 17360 0 _0620_
rlabel metal3 24248 23800 24248 23800 0 _0621_
rlabel metal2 23912 22680 23912 22680 0 _0622_
rlabel metal2 24696 24024 24696 24024 0 _0623_
rlabel metal2 24360 24304 24360 24304 0 _0624_
rlabel metal3 22288 23912 22288 23912 0 _0625_
rlabel metal2 17864 23296 17864 23296 0 _0626_
rlabel metal2 18536 24192 18536 24192 0 _0627_
rlabel metal3 18704 23128 18704 23128 0 _0628_
rlabel metal2 22512 21112 22512 21112 0 _0629_
rlabel metal2 24920 20888 24920 20888 0 _0630_
rlabel metal2 20328 23128 20328 23128 0 _0631_
rlabel metal2 29288 25480 29288 25480 0 _0632_
rlabel metal3 27720 26488 27720 26488 0 _0633_
rlabel metal2 22680 22624 22680 22624 0 _0634_
rlabel metal2 24416 17080 24416 17080 0 _0635_
rlabel metal2 32536 27216 32536 27216 0 _0636_
rlabel metal2 31416 24920 31416 24920 0 _0637_
rlabel metal2 52920 24192 52920 24192 0 _0638_
rlabel metal3 54488 22904 54488 22904 0 _0639_
rlabel metal2 49336 21504 49336 21504 0 _0640_
rlabel metal2 54824 26320 54824 26320 0 _0641_
rlabel metal2 53480 23632 53480 23632 0 _0642_
rlabel metal2 51352 25088 51352 25088 0 _0643_
rlabel metal2 34216 25536 34216 25536 0 _0644_
rlabel metal2 58240 12824 58240 12824 0 _0645_
rlabel metal2 50064 24472 50064 24472 0 _0646_
rlabel metal2 46312 19600 46312 19600 0 _0647_
rlabel metal3 44352 20776 44352 20776 0 _0648_
rlabel metal2 47432 20664 47432 20664 0 _0649_
rlabel metal3 48328 20104 48328 20104 0 _0650_
rlabel metal2 45472 21784 45472 21784 0 _0651_
rlabel metal2 44744 23688 44744 23688 0 _0652_
rlabel via2 49000 21560 49000 21560 0 _0653_
rlabel metal2 46648 22064 46648 22064 0 _0654_
rlabel metal2 47936 24696 47936 24696 0 _0655_
rlabel metal2 48328 23912 48328 23912 0 _0656_
rlabel metal2 49672 23520 49672 23520 0 _0657_
rlabel metal2 53592 23688 53592 23688 0 _0658_
rlabel metal2 46872 23744 46872 23744 0 _0659_
rlabel metal2 48888 21952 48888 21952 0 _0660_
rlabel metal3 50456 22232 50456 22232 0 _0661_
rlabel metal3 49560 23912 49560 23912 0 _0662_
rlabel metal2 49336 25144 49336 25144 0 _0663_
rlabel metal3 44296 21224 44296 21224 0 _0664_
rlabel metal2 33096 22792 33096 22792 0 _0665_
rlabel metal2 31640 20664 31640 20664 0 _0666_
rlabel metal2 31976 19656 31976 19656 0 _0667_
rlabel metal2 26040 24808 26040 24808 0 _0668_
rlabel metal2 25704 25200 25704 25200 0 _0669_
rlabel metal2 30856 17192 30856 17192 0 _0670_
rlabel metal2 32032 16632 32032 16632 0 _0671_
rlabel metal2 30744 17192 30744 17192 0 _0672_
rlabel metal2 32536 20104 32536 20104 0 _0673_
rlabel metal2 33544 22176 33544 22176 0 _0674_
rlabel metal3 32928 20888 32928 20888 0 _0675_
rlabel metal3 32872 21784 32872 21784 0 _0676_
rlabel metal2 32648 23128 32648 23128 0 _0677_
rlabel metal2 30800 20104 30800 20104 0 _0678_
rlabel metal3 25144 16072 25144 16072 0 _0679_
rlabel metal2 24752 13832 24752 13832 0 _0680_
rlabel metal2 24192 16856 24192 16856 0 _0681_
rlabel metal3 26264 15176 26264 15176 0 _0682_
rlabel metal2 21672 15064 21672 15064 0 _0683_
rlabel metal2 19096 17976 19096 17976 0 _0684_
rlabel metal3 22176 12264 22176 12264 0 _0685_
rlabel metal2 50680 10136 50680 10136 0 _0686_
rlabel metal3 48776 12824 48776 12824 0 _0687_
rlabel metal3 48160 10584 48160 10584 0 _0688_
rlabel metal2 53144 11312 53144 11312 0 _0689_
rlabel metal2 51240 10416 51240 10416 0 _0690_
rlabel metal2 22792 16072 22792 16072 0 _0691_
rlabel metal2 51688 6832 51688 6832 0 _0692_
rlabel metal3 48776 8904 48776 8904 0 _0693_
rlabel metal2 46424 5936 46424 5936 0 _0694_
rlabel metal2 45976 6720 45976 6720 0 _0695_
rlabel metal3 46144 6664 46144 6664 0 _0696_
rlabel metal2 45416 7504 45416 7504 0 _0697_
rlabel metal2 45864 7168 45864 7168 0 _0698_
rlabel metal2 47488 19768 47488 19768 0 _0699_
rlabel metal2 46536 12096 46536 12096 0 _0700_
rlabel metal2 45080 8512 45080 8512 0 _0701_
rlabel metal2 47992 8904 47992 8904 0 _0702_
rlabel metal2 48776 6272 48776 6272 0 _0703_
rlabel metal2 51688 8512 51688 8512 0 _0704_
rlabel metal2 51016 10248 51016 10248 0 _0705_
rlabel metal2 49336 9744 49336 9744 0 _0706_
rlabel metal2 45976 11088 45976 11088 0 _0707_
rlabel metal2 48888 9072 48888 9072 0 _0708_
rlabel metal2 48216 9464 48216 9464 0 _0709_
rlabel metal3 45528 10024 45528 10024 0 _0710_
rlabel metal2 47208 12320 47208 12320 0 _0711_
rlabel metal2 24360 13048 24360 13048 0 _0712_
rlabel metal2 23688 12040 23688 12040 0 _0713_
rlabel metal2 24584 11256 24584 11256 0 _0714_
rlabel metal2 21112 12544 21112 12544 0 _0715_
rlabel metal2 30296 16968 30296 16968 0 _0716_
rlabel metal2 22680 13104 22680 13104 0 _0717_
rlabel metal3 22344 11368 22344 11368 0 _0718_
rlabel metal2 16800 7224 16800 7224 0 _0719_
rlabel metal2 19096 11480 19096 11480 0 _0720_
rlabel metal2 20888 12152 20888 12152 0 _0721_
rlabel metal3 22120 12152 22120 12152 0 _0722_
rlabel metal2 24360 11088 24360 11088 0 _0723_
rlabel metal2 56952 13104 56952 13104 0 _0724_
rlabel metal3 23072 10584 23072 10584 0 _0725_
rlabel metal2 23800 11480 23800 11480 0 _0726_
rlabel metal2 23128 8344 23128 8344 0 _0727_
rlabel metal2 19600 12264 19600 12264 0 _0728_
rlabel metal2 19768 11648 19768 11648 0 _0729_
rlabel metal3 20776 10808 20776 10808 0 _0730_
rlabel metal3 23688 6552 23688 6552 0 _0731_
rlabel metal2 12432 12152 12432 12152 0 _0732_
rlabel metal2 16968 4704 16968 4704 0 _0733_
rlabel metal3 36288 5992 36288 5992 0 _0734_
rlabel metal2 37688 9856 37688 9856 0 _0735_
rlabel metal2 35448 8288 35448 8288 0 _0736_
rlabel metal3 9408 9240 9408 9240 0 _0737_
rlabel metal2 25592 6776 25592 6776 0 _0738_
rlabel metal2 37800 8904 37800 8904 0 _0739_
rlabel metal2 36344 7728 36344 7728 0 _0740_
rlabel metal2 31640 6048 31640 6048 0 _0741_
rlabel metal2 33544 4312 33544 4312 0 _0742_
rlabel metal2 45304 6384 45304 6384 0 _0743_
rlabel metal2 35672 5432 35672 5432 0 _0744_
rlabel metal2 34328 5488 34328 5488 0 _0745_
rlabel metal2 38808 6664 38808 6664 0 _0746_
rlabel metal2 39928 9296 39928 9296 0 _0747_
rlabel metal2 35504 6104 35504 6104 0 _0748_
rlabel metal3 20944 5768 20944 5768 0 _0749_
rlabel metal2 37016 8512 37016 8512 0 _0750_
rlabel metal2 34440 8288 34440 8288 0 _0751_
rlabel metal2 32424 8512 32424 8512 0 _0752_
rlabel metal3 34944 6552 34944 6552 0 _0753_
rlabel metal2 36344 6160 36344 6160 0 _0754_
rlabel metal2 32536 7168 32536 7168 0 _0755_
rlabel metal3 34272 9800 34272 9800 0 _0756_
rlabel metal2 15288 9184 15288 9184 0 _0757_
rlabel metal2 13160 10304 13160 10304 0 _0758_
rlabel metal2 11032 16072 11032 16072 0 _0759_
rlabel metal3 11144 11592 11144 11592 0 _0760_
rlabel metal3 13664 9240 13664 9240 0 _0761_
rlabel metal2 11928 10472 11928 10472 0 _0762_
rlabel metal2 20328 10696 20328 10696 0 _0763_
rlabel metal3 10696 10584 10696 10584 0 _0764_
rlabel metal2 9800 11648 9800 11648 0 _0765_
rlabel metal2 12264 10976 12264 10976 0 _0766_
rlabel metal3 13384 12264 13384 12264 0 _0767_
rlabel metal3 13496 10584 13496 10584 0 _0768_
rlabel metal2 13048 10696 13048 10696 0 _0769_
rlabel metal2 12824 11088 12824 11088 0 _0770_
rlabel metal2 6216 14224 6216 14224 0 _0771_
rlabel metal3 7112 10808 7112 10808 0 _0772_
rlabel metal2 6328 14336 6328 14336 0 _0773_
rlabel metal2 52136 6272 52136 6272 0 _0774_
rlabel metal3 40656 23352 40656 23352 0 _0775_
rlabel metal3 40992 23688 40992 23688 0 _0776_
rlabel metal2 39928 28728 39928 28728 0 _0777_
rlabel metal3 40824 23912 40824 23912 0 _0778_
rlabel metal2 41944 22736 41944 22736 0 _0779_
rlabel metal2 41496 19768 41496 19768 0 _0780_
rlabel metal2 40600 21784 40600 21784 0 _0781_
rlabel metal3 37688 24696 37688 24696 0 _0782_
rlabel metal2 38864 23464 38864 23464 0 _0783_
rlabel metal2 35896 22624 35896 22624 0 _0784_
rlabel metal2 46088 26040 46088 26040 0 _0785_
rlabel metal2 26712 27328 26712 27328 0 _0786_
rlabel metal2 25648 26936 25648 26936 0 _0787_
rlabel metal2 45416 27440 45416 27440 0 _0788_
rlabel metal2 46760 28896 46760 28896 0 _0789_
rlabel metal2 56952 30688 56952 30688 0 _0790_
rlabel metal2 62216 28504 62216 28504 0 _0791_
rlabel metal2 61712 32648 61712 32648 0 _0792_
rlabel metal2 58408 30520 58408 30520 0 _0793_
rlabel metal2 45640 28504 45640 28504 0 _0794_
rlabel metal3 44968 35952 44968 35952 0 _0795_
rlabel metal2 61096 32256 61096 32256 0 _0796_
rlabel metal2 58800 27832 58800 27832 0 _0797_
rlabel metal2 61208 22288 61208 22288 0 _0798_
rlabel metal2 59080 22848 59080 22848 0 _0799_
rlabel metal2 57288 21728 57288 21728 0 _0800_
rlabel metal2 57288 25312 57288 25312 0 _0801_
rlabel metal3 57512 24808 57512 24808 0 _0802_
rlabel metal2 53312 29400 53312 29400 0 _0803_
rlabel metal2 51296 28840 51296 28840 0 _0804_
rlabel metal3 55048 29400 55048 29400 0 _0805_
rlabel metal2 58520 25256 58520 25256 0 _0806_
rlabel metal2 60200 26544 60200 26544 0 _0807_
rlabel metal2 58856 25312 58856 25312 0 _0808_
rlabel metal2 56616 29232 56616 29232 0 _0809_
rlabel metal2 58240 27832 58240 27832 0 _0810_
rlabel metal3 56952 28504 56952 28504 0 _0811_
rlabel metal2 61320 30912 61320 30912 0 _0812_
rlabel metal2 57736 28336 57736 28336 0 _0813_
rlabel metal2 58632 26040 58632 26040 0 _0814_
rlabel metal2 61208 28952 61208 28952 0 _0815_
rlabel metal2 60424 26208 60424 26208 0 _0816_
rlabel metal2 55384 30240 55384 30240 0 _0817_
rlabel metal2 50120 27608 50120 27608 0 _0818_
rlabel metal3 47712 27272 47712 27272 0 _0819_
rlabel metal2 47544 24360 47544 24360 0 _0820_
rlabel metal2 49784 20384 49784 20384 0 _0821_
rlabel metal2 47880 22848 47880 22848 0 _0822_
rlabel metal2 45976 23352 45976 23352 0 _0823_
rlabel metal2 45416 25760 45416 25760 0 _0824_
rlabel metal2 42504 24920 42504 24920 0 _0825_
rlabel metal2 45640 25928 45640 25928 0 _0826_
rlabel metal3 47320 26936 47320 26936 0 _0827_
rlabel metal2 47208 28448 47208 28448 0 _0828_
rlabel metal2 47320 26376 47320 26376 0 _0829_
rlabel metal2 47096 25816 47096 25816 0 _0830_
rlabel metal2 47880 20776 47880 20776 0 _0831_
rlabel metal3 49560 24640 49560 24640 0 _0832_
rlabel metal2 47992 20944 47992 20944 0 _0833_
rlabel metal2 48496 17528 48496 17528 0 _0834_
rlabel metal3 44520 17640 44520 17640 0 _0835_
rlabel metal2 35840 19208 35840 19208 0 _0836_
rlabel metal2 42840 18480 42840 18480 0 _0837_
rlabel metal2 55720 18704 55720 18704 0 _0838_
rlabel metal2 54544 17528 54544 17528 0 _0839_
rlabel metal2 55496 16856 55496 16856 0 _0840_
rlabel metal2 56168 21616 56168 21616 0 _0841_
rlabel metal2 53928 19936 53928 19936 0 _0842_
rlabel metal2 39480 19320 39480 19320 0 _0843_
rlabel metal2 54544 9240 54544 9240 0 _0844_
rlabel metal3 53928 18424 53928 18424 0 _0845_
rlabel metal3 52976 13720 52976 13720 0 _0846_
rlabel metal2 54488 13720 54488 13720 0 _0847_
rlabel metal2 49896 15232 49896 15232 0 _0848_
rlabel metal2 55384 16016 55384 16016 0 _0849_
rlabel metal2 54936 16072 54936 16072 0 _0850_
rlabel metal3 60816 21000 60816 21000 0 _0851_
rlabel metal2 55832 14868 55832 14868 0 _0852_
rlabel metal2 56056 14504 56056 14504 0 _0853_
rlabel metal2 55832 18032 55832 18032 0 _0854_
rlabel metal2 62216 18200 62216 18200 0 _0855_
rlabel metal2 54040 18480 54040 18480 0 _0856_
rlabel metal2 53368 18312 53368 18312 0 _0857_
rlabel metal2 56280 19936 56280 19936 0 _0858_
rlabel metal2 57064 18256 57064 18256 0 _0859_
rlabel metal2 55272 14812 55272 14812 0 _0860_
rlabel metal2 55048 14448 55048 14448 0 _0861_
rlabel metal2 57400 18088 57400 18088 0 _0862_
rlabel metal2 52360 18088 52360 18088 0 _0863_
rlabel metal2 43176 18312 43176 18312 0 _0864_
rlabel metal2 44800 17864 44800 17864 0 _0865_
rlabel metal3 45528 18984 45528 18984 0 _0866_
rlabel metal2 45192 17976 45192 17976 0 _0867_
rlabel metal2 48664 24584 48664 24584 0 _0868_
rlabel metal2 45640 18984 45640 18984 0 _0869_
rlabel metal2 48440 6776 48440 6776 0 _0870_
rlabel metal3 46200 9016 46200 9016 0 _0871_
rlabel metal2 46200 11816 46200 11816 0 _0872_
rlabel metal2 45080 17864 45080 17864 0 _0873_
rlabel metal3 46200 19096 46200 19096 0 _0874_
rlabel metal2 40040 18088 40040 18088 0 _0875_
rlabel metal2 40208 17640 40208 17640 0 _0876_
rlabel metal2 40152 15624 40152 15624 0 _0877_
rlabel metal3 46368 9128 46368 9128 0 _0878_
rlabel metal3 46256 9576 46256 9576 0 _0879_
rlabel metal2 48944 12152 48944 12152 0 _0880_
rlabel metal2 45752 8792 45752 8792 0 _0881_
rlabel metal2 47544 6944 47544 6944 0 _0882_
rlabel metal2 59584 12376 59584 12376 0 _0883_
rlabel metal2 47208 6272 47208 6272 0 _0884_
rlabel metal2 40096 9016 40096 9016 0 _0885_
rlabel metal3 17248 11592 17248 11592 0 _0886_
rlabel metal2 55048 9128 55048 9128 0 _0887_
rlabel metal2 41496 9296 41496 9296 0 _0888_
rlabel metal3 41776 8008 41776 8008 0 _0889_
rlabel metal2 41720 12208 41720 12208 0 _0890_
rlabel metal2 43680 14392 43680 14392 0 _0891_
rlabel metal2 43288 18872 43288 18872 0 _0892_
rlabel metal3 43008 17528 43008 17528 0 _0893_
rlabel metal2 42504 6496 42504 6496 0 _0894_
rlabel metal3 43624 15288 43624 15288 0 _0895_
rlabel metal2 42616 17192 42616 17192 0 _0896_
rlabel metal2 43176 16744 43176 16744 0 _0897_
rlabel metal3 37912 14504 37912 14504 0 _0898_
rlabel metal3 40432 13608 40432 13608 0 _0899_
rlabel metal2 39984 15512 39984 15512 0 _0900_
rlabel metal2 38920 13664 38920 13664 0 _0901_
rlabel metal2 39256 12992 39256 12992 0 _0902_
rlabel metal2 39928 15148 39928 15148 0 _0903_
rlabel metal3 56280 13720 56280 13720 0 _0904_
rlabel metal3 53928 14448 53928 14448 0 _0905_
rlabel metal3 44912 13720 44912 13720 0 _0906_
rlabel metal2 42616 14000 42616 14000 0 _0907_
rlabel metal2 41888 15736 41888 15736 0 _0908_
rlabel metal2 41440 13944 41440 13944 0 _0909_
rlabel metal2 42560 12040 42560 12040 0 _0910_
rlabel metal2 42952 16016 42952 16016 0 _0911_
rlabel metal2 47600 16856 47600 16856 0 _0912_
rlabel metal2 42168 13720 42168 13720 0 _0913_
rlabel metal2 42000 16184 42000 16184 0 _0914_
rlabel metal2 48160 16856 48160 16856 0 _0915_
rlabel metal2 42392 11424 42392 11424 0 _0916_
rlabel metal2 41048 10752 41048 10752 0 _0917_
rlabel metal2 41720 9688 41720 9688 0 _0918_
rlabel metal2 34776 8064 34776 8064 0 _0919_
rlabel metal2 39032 8176 39032 8176 0 _0920_
rlabel metal2 38696 8904 38696 8904 0 _0921_
rlabel metal2 39816 7784 39816 7784 0 _0922_
rlabel metal2 44184 9296 44184 9296 0 _0923_
rlabel metal2 41552 7672 41552 7672 0 _0924_
rlabel metal2 41328 7672 41328 7672 0 _0925_
rlabel metal2 42784 9016 42784 9016 0 _0926_
rlabel metal2 40152 9520 40152 9520 0 _0927_
rlabel metal3 52864 7672 52864 7672 0 _0928_
rlabel metal2 40320 9800 40320 9800 0 _0929_
rlabel metal2 32984 7392 32984 7392 0 _0930_
rlabel metal2 35784 7168 35784 7168 0 _0931_
rlabel metal2 39256 7784 39256 7784 0 _0932_
rlabel metal2 39592 6776 39592 6776 0 _0933_
rlabel metal2 40152 5488 40152 5488 0 _0934_
rlabel metal2 25704 10528 25704 10528 0 _0935_
rlabel metal2 25032 9520 25032 9520 0 _0936_
rlabel metal2 25816 12264 25816 12264 0 _0937_
rlabel metal2 26880 9128 26880 9128 0 _0938_
rlabel metal2 25368 10696 25368 10696 0 _0939_
rlabel metal2 38472 14224 38472 14224 0 _0940_
rlabel metal2 34440 13608 34440 13608 0 _0941_
rlabel metal2 33096 14896 33096 14896 0 _0942_
rlabel metal2 30856 14000 30856 14000 0 _0943_
rlabel metal2 31752 33376 31752 33376 0 _0944_
rlabel metal2 25704 5264 25704 5264 0 _0945_
rlabel metal2 26040 11480 26040 11480 0 _0946_
rlabel metal2 28616 10752 28616 10752 0 _0947_
rlabel metal2 28056 11816 28056 11816 0 _0948_
rlabel metal3 29512 11592 29512 11592 0 _0949_
rlabel metal2 25256 9576 25256 9576 0 _0950_
rlabel metal2 25536 9240 25536 9240 0 _0951_
rlabel metal2 30520 10696 30520 10696 0 _0952_
rlabel metal3 34832 12824 34832 12824 0 _0953_
rlabel metal2 30968 15540 30968 15540 0 _0954_
rlabel metal2 34552 12992 34552 12992 0 _0955_
rlabel metal2 28280 11312 28280 11312 0 _0956_
rlabel metal2 29624 14616 29624 14616 0 _0957_
rlabel metal2 26824 11648 26824 11648 0 _0958_
rlabel metal2 29848 9464 29848 9464 0 _0959_
rlabel metal2 28392 9352 28392 9352 0 _0960_
rlabel metal2 30520 7168 30520 7168 0 _0961_
rlabel metal2 28280 6944 28280 6944 0 _0962_
rlabel metal2 29960 7616 29960 7616 0 _0963_
rlabel metal2 34328 7728 34328 7728 0 _0964_
rlabel metal2 30296 7280 30296 7280 0 _0965_
rlabel metal2 28504 6664 28504 6664 0 _0966_
rlabel metal2 30072 8232 30072 8232 0 _0967_
rlabel metal3 29232 8904 29232 8904 0 _0968_
rlabel metal2 29176 18424 29176 18424 0 _0969_
rlabel metal2 52024 28000 52024 28000 0 _0970_
rlabel metal2 47992 43848 47992 43848 0 _0971_
rlabel metal2 50176 40936 50176 40936 0 _0972_
rlabel metal2 39816 28168 39816 28168 0 _0973_
rlabel metal3 43176 27664 43176 27664 0 _0974_
rlabel metal2 50456 29736 50456 29736 0 _0975_
rlabel metal2 52696 29064 52696 29064 0 _0976_
rlabel metal2 30184 14056 30184 14056 0 _0977_
rlabel metal2 32312 11760 32312 11760 0 _0978_
rlabel metal3 32536 13720 32536 13720 0 _0979_
rlabel metal2 29344 13048 29344 13048 0 _0980_
rlabel metal2 57848 13216 57848 13216 0 _0981_
rlabel metal3 59248 26600 59248 26600 0 _0982_
rlabel metal2 56784 29176 56784 29176 0 _0983_
rlabel metal2 56840 27216 56840 27216 0 _0984_
rlabel metal2 55272 28056 55272 28056 0 _0985_
rlabel metal3 54152 27720 54152 27720 0 _0986_
rlabel metal3 51800 27048 51800 27048 0 _0987_
rlabel metal2 62384 51240 62384 51240 0 _0988_
rlabel metal2 53648 27048 53648 27048 0 _0989_
rlabel metal3 52360 26824 52360 26824 0 _0990_
rlabel metal2 52080 27272 52080 27272 0 _0991_
rlabel metal2 50904 30464 50904 30464 0 _0992_
rlabel metal2 61096 14672 61096 14672 0 _0993_
rlabel metal3 56448 29512 56448 29512 0 _0994_
rlabel metal2 55832 29288 55832 29288 0 _0995_
rlabel metal2 56000 29176 56000 29176 0 _0996_
rlabel metal2 62888 24696 62888 24696 0 _0997_
rlabel metal3 59752 21560 59752 21560 0 _0998_
rlabel metal2 54600 28112 54600 28112 0 _0999_
rlabel metal2 55048 21784 55048 21784 0 _1000_
rlabel metal2 53368 24640 53368 24640 0 _1001_
rlabel metal2 55272 21616 55272 21616 0 _1002_
rlabel metal3 57624 20160 57624 20160 0 _1003_
rlabel metal3 59584 26488 59584 26488 0 _1004_
rlabel metal2 61040 23912 61040 23912 0 _1005_
rlabel metal2 58520 20440 58520 20440 0 _1006_
rlabel metal3 59472 17640 59472 17640 0 _1007_
rlabel metal3 57456 19208 57456 19208 0 _1008_
rlabel metal2 57680 18648 57680 18648 0 _1009_
rlabel metal3 58520 21000 58520 21000 0 _1010_
rlabel metal2 53928 21112 53928 21112 0 _1011_
rlabel metal3 56280 20776 56280 20776 0 _1012_
rlabel metal3 59920 20776 59920 20776 0 _1013_
rlabel metal2 60536 21392 60536 21392 0 _1014_
rlabel metal3 56784 16968 56784 16968 0 _1015_
rlabel metal2 57736 17192 57736 17192 0 _1016_
rlabel metal2 57400 14504 57400 14504 0 _1017_
rlabel metal2 56616 13216 56616 13216 0 _1018_
rlabel metal2 50064 13720 50064 13720 0 _1019_
rlabel metal3 60312 14000 60312 14000 0 _1020_
rlabel metal2 48888 17248 48888 17248 0 _1021_
rlabel metal2 48776 11816 48776 11816 0 _1022_
rlabel metal2 49280 16296 49280 16296 0 _1023_
rlabel metal2 49560 14056 49560 14056 0 _1024_
rlabel metal3 60088 17864 60088 17864 0 _1025_
rlabel metal3 50260 15400 50260 15400 0 _1026_
rlabel metal2 47432 16576 47432 16576 0 _1027_
rlabel metal2 42224 16856 42224 16856 0 _1028_
rlabel metal3 45360 15960 45360 15960 0 _1029_
rlabel metal2 48664 13944 48664 13944 0 _1030_
rlabel metal2 49616 15176 49616 15176 0 _1031_
rlabel metal2 50288 13832 50288 13832 0 _1032_
rlabel metal2 49168 15288 49168 15288 0 _1033_
rlabel metal2 49336 15568 49336 15568 0 _1034_
rlabel metal2 49560 16240 49560 16240 0 _1035_
rlabel metal2 41328 16072 41328 16072 0 _1036_
rlabel metal2 41552 16856 41552 16856 0 _1037_
rlabel metal3 40544 16856 40544 16856 0 _1038_
rlabel metal2 59304 12992 59304 12992 0 _1039_
rlabel metal2 38920 16688 38920 16688 0 _1040_
rlabel metal2 35336 16744 35336 16744 0 _1041_
rlabel metal2 34104 10248 34104 10248 0 _1042_
rlabel metal2 35000 15904 35000 15904 0 _1043_
rlabel metal2 51800 5852 51800 5852 0 _1044_
rlabel metal3 50540 13944 50540 13944 0 _1045_
rlabel metal2 35000 17920 35000 17920 0 _1046_
rlabel metal2 35560 17136 35560 17136 0 _1047_
rlabel metal2 47320 14784 47320 14784 0 _1048_
rlabel metal2 36680 13440 36680 13440 0 _1049_
rlabel metal2 35672 13328 35672 13328 0 _1050_
rlabel metal3 34272 14728 34272 14728 0 _1051_
rlabel metal2 36120 15988 36120 15988 0 _1052_
rlabel metal2 34328 15288 34328 15288 0 _1053_
rlabel metal3 35840 15848 35840 15848 0 _1054_
rlabel metal2 34328 14672 34328 14672 0 _1055_
rlabel metal2 33544 15624 33544 15624 0 _1056_
rlabel metal2 25424 12376 25424 12376 0 _1057_
rlabel metal2 28616 14392 28616 14392 0 _1058_
rlabel metal2 28504 15176 28504 15176 0 _1059_
rlabel metal2 54824 41720 54824 41720 0 _1060_
rlabel metal2 56672 46760 56672 46760 0 _1061_
rlabel metal2 56840 46872 56840 46872 0 _1062_
rlabel metal2 52696 41552 52696 41552 0 _1063_
rlabel metal2 55496 40768 55496 40768 0 _1064_
rlabel metal2 55608 43848 55608 43848 0 _1065_
rlabel metal2 48104 45360 48104 45360 0 _1066_
rlabel metal2 53928 43400 53928 43400 0 _1067_
rlabel metal2 52024 40152 52024 40152 0 _1068_
rlabel metal3 62188 47320 62188 47320 0 _1069_
rlabel metal2 57400 31248 57400 31248 0 _1070_
rlabel metal2 61992 47936 61992 47936 0 _1071_
rlabel metal2 58968 49280 58968 49280 0 _1072_
rlabel metal2 57288 46480 57288 46480 0 _1073_
rlabel metal3 56896 42952 56896 42952 0 _1074_
rlabel metal3 55776 46872 55776 46872 0 _1075_
rlabel metal3 56672 41384 56672 41384 0 _1076_
rlabel metal2 58240 41944 58240 41944 0 _1077_
rlabel metal2 62272 46648 62272 46648 0 _1078_
rlabel metal2 57904 42168 57904 42168 0 _1079_
rlabel metal2 54936 41888 54936 41888 0 _1080_
rlabel metal3 57512 43736 57512 43736 0 _1081_
rlabel metal2 53928 46984 53928 46984 0 _1082_
rlabel metal2 60760 42000 60760 42000 0 _1083_
rlabel metal3 57568 41160 57568 41160 0 _1084_
rlabel metal2 61656 36288 61656 36288 0 _1085_
rlabel metal3 58688 37352 58688 37352 0 _1086_
rlabel metal2 56616 37632 56616 37632 0 _1087_
rlabel metal3 55608 37240 55608 37240 0 _1088_
rlabel metal2 53536 38584 53536 38584 0 _1089_
rlabel metal2 53928 33432 53928 33432 0 _1090_
rlabel metal2 51800 18200 51800 18200 0 _1091_
rlabel metal2 52752 19432 52752 19432 0 _1092_
rlabel metal2 48440 44576 48440 44576 0 _1093_
rlabel metal2 54936 34552 54936 34552 0 _1094_
rlabel metal2 53256 34216 53256 34216 0 _1095_
rlabel metal2 55608 34216 55608 34216 0 _1096_
rlabel metal2 52360 34776 52360 34776 0 _1097_
rlabel metal2 46424 36344 46424 36344 0 _1098_
rlabel metal2 52808 36008 52808 36008 0 _1099_
rlabel metal2 53592 35336 53592 35336 0 _1100_
rlabel metal2 61992 36512 61992 36512 0 _1101_
rlabel via2 55496 35224 55496 35224 0 _1102_
rlabel metal2 55944 34496 55944 34496 0 _1103_
rlabel metal2 53592 33712 53592 33712 0 _1104_
rlabel metal2 53368 34440 53368 34440 0 _1105_
rlabel metal2 46648 38080 46648 38080 0 _1106_
rlabel metal2 48104 36736 48104 36736 0 _1107_
rlabel metal2 48272 36456 48272 36456 0 _1108_
rlabel metal2 47768 36456 47768 36456 0 _1109_
rlabel metal2 46088 38416 46088 38416 0 _1110_
rlabel metal2 42000 39592 42000 39592 0 _1111_
rlabel metal2 41832 12096 41832 12096 0 _1112_
rlabel metal3 42728 23800 42728 23800 0 _1113_
rlabel metal2 41384 40488 41384 40488 0 _1114_
rlabel metal3 42112 38248 42112 38248 0 _1115_
rlabel metal3 44968 38024 44968 38024 0 _1116_
rlabel metal2 43848 37912 43848 37912 0 _1117_
rlabel metal2 39928 36176 39928 36176 0 _1118_
rlabel metal2 40936 34944 40936 34944 0 _1119_
rlabel metal2 42392 36120 42392 36120 0 _1120_
rlabel metal3 43344 35560 43344 35560 0 _1121_
rlabel metal2 46872 37240 46872 37240 0 _1122_
rlabel metal3 44464 36568 44464 36568 0 _1123_
rlabel metal2 44184 37856 44184 37856 0 _1124_
rlabel metal3 42560 38808 42560 38808 0 _1125_
rlabel metal2 41832 38528 41832 38528 0 _1126_
rlabel metal2 40152 36008 40152 36008 0 _1127_
rlabel metal2 40096 40040 40096 40040 0 _1128_
rlabel metal2 39928 40376 39928 40376 0 _1129_
rlabel metal2 40600 40376 40600 40376 0 _1130_
rlabel metal2 40488 33040 40488 33040 0 _1131_
rlabel metal3 31864 31640 31864 31640 0 _1132_
rlabel metal2 26712 10864 26712 10864 0 _1133_
rlabel metal3 30800 31528 30800 31528 0 _1134_
rlabel metal2 33208 36344 33208 36344 0 _1135_
rlabel metal2 33656 34048 33656 34048 0 _1136_
rlabel metal3 34104 32536 34104 32536 0 _1137_
rlabel metal2 36120 32928 36120 32928 0 _1138_
rlabel metal2 42952 36064 42952 36064 0 _1139_
rlabel metal2 35784 31640 35784 31640 0 _1140_
rlabel metal2 36008 31808 36008 31808 0 _1141_
rlabel metal2 35896 32368 35896 32368 0 _1142_
rlabel metal3 33992 30184 33992 30184 0 _1143_
rlabel metal2 34216 30408 34216 30408 0 _1144_
rlabel metal2 34552 28728 34552 28728 0 _1145_
rlabel metal2 34888 30184 34888 30184 0 _1146_
rlabel metal2 36064 29400 36064 29400 0 _1147_
rlabel metal2 39032 29176 39032 29176 0 _1148_
rlabel metal2 36680 28504 36680 28504 0 _1149_
rlabel metal2 34888 28392 34888 28392 0 _1150_
rlabel metal2 33208 26684 33208 26684 0 _1151_
rlabel metal2 33880 28392 33880 28392 0 _1152_
rlabel metal3 41720 55272 41720 55272 0 _1153_
rlabel metal2 45080 55048 45080 55048 0 _1154_
rlabel metal2 44744 54936 44744 54936 0 _1155_
rlabel metal2 43400 54656 43400 54656 0 _1156_
rlabel metal2 51576 49672 51576 49672 0 _1157_
rlabel metal2 51408 49224 51408 49224 0 _1158_
rlabel metal2 51128 48048 51128 48048 0 _1159_
rlabel metal2 53256 45024 53256 45024 0 _1160_
rlabel metal3 43512 40600 43512 40600 0 _1161_
rlabel metal2 42616 42448 42616 42448 0 _1162_
rlabel metal2 42728 40992 42728 40992 0 _1163_
rlabel metal2 42504 40656 42504 40656 0 _1164_
rlabel metal2 32984 40320 32984 40320 0 _1165_
rlabel metal3 31024 41832 31024 41832 0 _1166_
rlabel metal2 32536 41440 32536 41440 0 _1167_
rlabel metal2 32200 41328 32200 41328 0 _1168_
rlabel metal2 29680 55384 29680 55384 0 _1169_
rlabel metal3 30968 56056 30968 56056 0 _1170_
rlabel metal2 32088 56504 32088 56504 0 _1171_
rlabel metal3 31304 55496 31304 55496 0 _1172_
rlabel metal2 31304 46424 31304 46424 0 _1173_
rlabel metal2 37688 48832 37688 48832 0 _1174_
rlabel metal2 36792 48552 36792 48552 0 _1175_
rlabel metal3 37240 48160 37240 48160 0 _1176_
rlabel metal2 12152 49336 12152 49336 0 _1177_
rlabel metal2 13272 47264 13272 47264 0 _1178_
rlabel metal2 13160 46928 13160 46928 0 _1179_
rlabel metal2 11256 45360 11256 45360 0 _1180_
rlabel metal2 2408 36568 2408 36568 0 _1181_
rlabel metal2 2632 37520 2632 37520 0 _1182_
rlabel metal3 7616 43288 7616 43288 0 _1183_
rlabel metal2 5208 44744 5208 44744 0 _1184_
rlabel metal2 2744 44968 2744 44968 0 _1185_
rlabel metal3 1400 38920 1400 38920 0 _1186_
rlabel metal2 14392 52472 14392 52472 0 _1187_
rlabel metal2 15400 55552 15400 55552 0 _1188_
rlabel metal2 15008 54712 15008 54712 0 _1189_
rlabel metal3 17220 57512 17220 57512 0 _1190_
rlabel metal2 28168 43456 28168 43456 0 _1191_
rlabel metal3 24136 43512 24136 43512 0 _1192_
rlabel metal2 26488 43904 26488 43904 0 _1193_
rlabel metal2 27720 45584 27720 45584 0 _1194_
rlabel metal2 17472 35896 17472 35896 0 _1195_
rlabel metal2 14056 40376 14056 40376 0 _1196_
rlabel metal3 17472 38920 17472 38920 0 _1197_
rlabel metal2 17864 41944 17864 41944 0 _1198_
rlabel metal2 2520 34608 2520 34608 0 _1199_
rlabel metal2 5880 35672 5880 35672 0 _1200_
rlabel metal3 7280 27160 7280 27160 0 _1201_
rlabel metal2 7616 38808 7616 38808 0 _1202_
rlabel metal2 7952 38584 7952 38584 0 _1203_
rlabel metal2 20888 31808 20888 31808 0 _1204_
rlabel metal2 16576 34664 16576 34664 0 _1205_
rlabel metal2 18424 34440 18424 34440 0 _1206_
rlabel metal2 23408 32760 23408 32760 0 _1207_
rlabel metal2 24136 18424 24136 18424 0 _1208_
rlabel metal2 14056 22848 14056 22848 0 _1209_
rlabel metal3 18648 25144 18648 25144 0 _1210_
rlabel metal2 22456 26180 22456 26180 0 _1211_
rlabel metal3 13216 18648 13216 18648 0 _1212_
rlabel metal2 14280 21448 14280 21448 0 _1213_
rlabel metal3 14112 18424 14112 18424 0 _1214_
rlabel metal2 13944 17808 13944 17808 0 _1215_
rlabel metal2 5712 15512 5712 15512 0 _1216_
rlabel metal2 5992 25816 5992 25816 0 _1217_
rlabel metal2 8792 22176 8792 22176 0 _1218_
rlabel metal2 7672 22680 7672 22680 0 _1219_
rlabel metal3 8456 24136 8456 24136 0 _1220_
rlabel metal2 6440 25816 6440 25816 0 _1221_
rlabel metal2 16296 20328 16296 20328 0 _1222_
rlabel metal3 23240 23184 23240 23184 0 _1223_
rlabel metal2 18032 24136 18032 24136 0 _1224_
rlabel metal2 17416 29064 17416 29064 0 _1225_
rlabel metal2 49672 24304 49672 24304 0 _1226_
rlabel metal2 29960 21112 29960 21112 0 _1227_
rlabel metal2 31640 24696 31640 24696 0 _1228_
rlabel metal3 31472 24696 31472 24696 0 _1229_
rlabel metal3 22400 12712 22400 12712 0 _1230_
rlabel metal2 19432 13048 19432 13048 0 _1231_
rlabel metal2 21672 12880 21672 12880 0 _1232_
rlabel metal3 20272 13720 20272 13720 0 _1233_
rlabel metal2 9688 7504 9688 7504 0 _1234_
rlabel metal2 8344 7784 8344 7784 0 _1235_
rlabel metal3 11872 9128 11872 9128 0 _1236_
rlabel metal2 7448 15736 7448 15736 0 _1237_
rlabel metal2 8232 7672 8232 7672 0 _1238_
rlabel metal3 45752 23352 45752 23352 0 _1239_
rlabel metal2 41720 21784 41720 21784 0 _1240_
rlabel metal2 44968 24640 44968 24640 0 _1241_
rlabel metal3 43680 26936 43680 26936 0 _1242_
rlabel metal2 43064 19376 43064 19376 0 _1243_
rlabel metal2 44520 18200 44520 18200 0 _1244_
rlabel metal2 44072 18536 44072 18536 0 _1245_
rlabel metal2 42392 19880 42392 19880 0 _1246_
rlabel metal2 43736 8176 43736 8176 0 _1247_
rlabel metal2 44744 7672 44744 7672 0 _1248_
rlabel metal3 43960 7560 43960 7560 0 _1249_
rlabel metal2 42952 7504 42952 7504 0 _1250_
rlabel metal3 27664 9016 27664 9016 0 _1251_
rlabel metal2 26152 9688 26152 9688 0 _1252_
rlabel metal2 32648 8568 32648 8568 0 _1253_
rlabel metal2 31528 7728 31528 7728 0 _1254_
rlabel metal2 30856 7784 30856 7784 0 _1255_
rlabel metal2 25928 8904 25928 8904 0 _1256_
rlabel metal2 47432 30632 47432 30632 0 _1257_
rlabel metal2 48216 42840 48216 42840 0 _1258_
rlabel metal2 47880 31080 47880 31080 0 _1259_
rlabel metal2 55608 27608 55608 27608 0 _1260_
rlabel metal3 49308 30968 49308 30968 0 _1261_
rlabel metal2 54264 23072 54264 23072 0 _1262_
rlabel metal2 54600 26264 54600 26264 0 _1263_
rlabel metal2 56728 24528 56728 24528 0 _1264_
rlabel metal2 61544 20776 61544 20776 0 _1265_
rlabel metal2 57064 23856 57064 23856 0 _1266_
rlabel metal2 49224 12432 49224 12432 0 _1267_
rlabel metal2 49336 17192 49336 17192 0 _1268_
rlabel metal3 50400 12824 50400 12824 0 _1269_
rlabel metal2 48104 14840 48104 14840 0 _1270_
rlabel metal2 51016 13328 51016 13328 0 _1271_
rlabel metal2 33320 11648 33320 11648 0 _1272_
rlabel metal2 33544 11704 33544 11704 0 _1273_
rlabel metal3 34216 10808 34216 10808 0 _1274_
rlabel metal2 33992 15932 33992 15932 0 _1275_
rlabel metal3 33544 11144 33544 11144 0 _1276_
rlabel metal2 60536 47376 60536 47376 0 _1277_
rlabel metal2 56952 46424 56952 46424 0 _1278_
rlabel metal2 57624 47096 57624 47096 0 _1279_
rlabel metal2 60872 45808 60872 45808 0 _1280_
rlabel metal2 61656 47124 61656 47124 0 _1281_
rlabel metal2 54208 34888 54208 34888 0 _1282_
rlabel metal3 58184 36344 58184 36344 0 _1283_
rlabel metal3 53592 36456 53592 36456 0 _1284_
rlabel metal2 54600 34832 54600 34832 0 _1285_
rlabel metal2 54544 33544 54544 33544 0 _1286_
rlabel metal2 41440 34328 41440 34328 0 _1287_
rlabel metal2 42952 35112 42952 35112 0 _1288_
rlabel metal2 42728 34440 42728 34440 0 _1289_
rlabel metal2 41944 34384 41944 34384 0 _1290_
rlabel metal2 43568 32760 43568 32760 0 _1291_
rlabel metal2 37128 33712 37128 33712 0 _1292_
rlabel metal2 37968 33544 37968 33544 0 _1293_
rlabel metal2 32200 33656 32200 33656 0 _1294_
rlabel metal2 33208 38668 33208 38668 0 _1295_
rlabel metal2 31416 34048 31416 34048 0 _1296_
rlabel metal2 35224 28784 35224 28784 0 _1297_
rlabel metal2 36456 29120 36456 29120 0 _1298_
rlabel metal2 48888 43848 48888 43848 0 _1299_
rlabel metal3 49672 45080 49672 45080 0 _1300_
rlabel metal2 50344 53704 50344 53704 0 _1301_
rlabel metal2 49168 53704 49168 53704 0 _1302_
rlabel metal2 45640 55552 45640 55552 0 _1303_
rlabel metal2 49336 55048 49336 55048 0 _1304_
rlabel metal2 49560 53592 49560 53592 0 _1305_
rlabel metal4 49224 50904 49224 50904 0 _1306_
rlabel metal2 48720 26488 48720 26488 0 _1307_
rlabel metal2 46984 29904 46984 29904 0 _1308_
rlabel metal2 49336 29904 49336 29904 0 _1309_
rlabel metal2 50344 47096 50344 47096 0 _1310_
rlabel metal2 50120 47432 50120 47432 0 _1311_
rlabel metal2 51016 44968 51016 44968 0 _1312_
rlabel metal2 54824 47936 54824 47936 0 _1313_
rlabel metal2 60928 47544 60928 47544 0 _1314_
rlabel metal2 54152 44520 54152 44520 0 _1315_
rlabel metal2 57064 42168 57064 42168 0 _1316_
rlabel metal3 57232 44184 57232 44184 0 _1317_
rlabel metal2 52024 43064 52024 43064 0 _1318_
rlabel metal2 39704 31472 39704 31472 0 _1319_
rlabel metal2 33432 31472 33432 31472 0 _1320_
rlabel metal2 38696 31780 38696 31780 0 _1321_
rlabel metal2 39480 33040 39480 33040 0 _1322_
rlabel metal3 39648 31752 39648 31752 0 _1323_
rlabel metal2 44184 40824 44184 40824 0 _1324_
rlabel metal2 58520 47600 58520 47600 0 _1325_
rlabel metal2 51800 44016 51800 44016 0 _1326_
rlabel metal2 48888 41272 48888 41272 0 _1327_
rlabel metal2 49784 44016 49784 44016 0 _1328_
rlabel metal2 50120 44464 50120 44464 0 _1329_
rlabel metal2 50008 47488 50008 47488 0 _1330_
rlabel metal2 49672 44576 49672 44576 0 _1331_
rlabel metal2 53144 44352 53144 44352 0 _1332_
rlabel metal2 49560 47096 49560 47096 0 _1333_
rlabel metal2 49224 44240 49224 44240 0 _1334_
rlabel metal2 49336 47656 49336 47656 0 _1335_
rlabel metal2 46536 53200 46536 53200 0 _1336_
rlabel metal2 20664 56560 20664 56560 0 _1337_
rlabel metal2 20216 56112 20216 56112 0 _1338_
rlabel metal3 21056 58520 21056 58520 0 _1339_
rlabel metal2 16128 59752 16128 59752 0 _1340_
rlabel metal2 16072 56896 16072 56896 0 _1341_
rlabel metal2 17192 57512 17192 57512 0 _1342_
rlabel metal2 15960 58688 15960 58688 0 _1343_
rlabel metal2 22008 57512 22008 57512 0 _1344_
rlabel metal2 48776 54992 48776 54992 0 _1345_
rlabel metal2 22792 56728 22792 56728 0 _1346_
rlabel metal3 24528 56056 24528 56056 0 _1347_
rlabel metal3 32816 59752 32816 59752 0 _1348_
rlabel metal2 31192 58016 31192 58016 0 _1349_
rlabel metal2 30184 58352 30184 58352 0 _1350_
rlabel metal2 27720 58744 27720 58744 0 _1351_
rlabel metal2 6104 47656 6104 47656 0 _1352_
rlabel metal2 2464 46648 2464 46648 0 _1353_
rlabel metal2 2744 46368 2744 46368 0 _1354_
rlabel metal2 5096 48496 5096 48496 0 _1355_
rlabel metal2 16968 58408 16968 58408 0 _1356_
rlabel metal2 26824 58352 26824 58352 0 _1357_
rlabel metal2 25760 57624 25760 57624 0 _1358_
rlabel metal2 18648 44800 18648 44800 0 _1359_
rlabel metal2 28168 58688 28168 58688 0 _1360_
rlabel metal2 20776 57176 20776 57176 0 _1361_
rlabel metal2 15512 57120 15512 57120 0 _1362_
rlabel metal2 24136 57120 24136 57120 0 _1363_
rlabel metal2 24416 56168 24416 56168 0 _1364_
rlabel metal2 31304 58576 31304 58576 0 _1365_
rlabel metal2 28056 57680 28056 57680 0 _1366_
rlabel metal2 24024 57792 24024 57792 0 _1367_
rlabel metal2 23464 56224 23464 56224 0 _1368_
rlabel metal3 41384 56728 41384 56728 0 _1369_
rlabel metal3 43232 53704 43232 53704 0 _1370_
rlabel metal3 47432 53032 47432 53032 0 _1371_
rlabel metal3 47040 53144 47040 53144 0 _1372_
rlabel metal2 46704 54488 46704 54488 0 _1373_
rlabel metal2 28728 40656 28728 40656 0 _1374_
rlabel metal2 30072 39368 30072 39368 0 _1375_
rlabel metal3 25760 38920 25760 38920 0 _1376_
rlabel metal2 34328 44016 34328 44016 0 _1377_
rlabel metal3 33992 42616 33992 42616 0 _1378_
rlabel metal2 34440 44744 34440 44744 0 _1379_
rlabel metal2 34216 44184 34216 44184 0 _1380_
rlabel metal2 30352 40488 30352 40488 0 _1381_
rlabel metal3 28560 39592 28560 39592 0 _1382_
rlabel metal2 29288 39088 29288 39088 0 _1383_
rlabel metal2 6328 38668 6328 38668 0 _1384_
rlabel metal3 2352 42616 2352 42616 0 _1385_
rlabel metal2 3920 40712 3920 40712 0 _1386_
rlabel metal3 5040 39368 5040 39368 0 _1387_
rlabel metal2 22680 35728 22680 35728 0 _1388_
rlabel metal2 29960 33040 29960 33040 0 _1389_
rlabel metal2 30072 32312 30072 32312 0 _1390_
rlabel metal2 31528 33320 31528 33320 0 _1391_
rlabel metal2 29624 34552 29624 34552 0 _1392_
rlabel metal2 28056 36792 28056 36792 0 _1393_
rlabel metal2 29288 35336 29288 35336 0 _1394_
rlabel metal3 27664 40264 27664 40264 0 _1395_
rlabel metal2 28616 39368 28616 39368 0 _1396_
rlabel metal2 31192 40544 31192 40544 0 _1397_
rlabel metal3 29176 39816 29176 39816 0 _1398_
rlabel metal2 31080 39760 31080 39760 0 _1399_
rlabel metal2 31640 35728 31640 35728 0 _1400_
rlabel metal2 31192 39872 31192 39872 0 _1401_
rlabel metal2 29064 40320 29064 40320 0 _1402_
rlabel metal2 45080 52752 45080 52752 0 _1403_
rlabel metal3 52136 53592 52136 53592 0 _1404_
rlabel metal2 55944 54152 55944 54152 0 _1405_
rlabel metal3 62440 15512 62440 15512 0 _1406_
rlabel metal2 60704 42952 60704 42952 0 _1407_
rlabel metal2 61208 46060 61208 46060 0 _1408_
rlabel metal2 62776 50232 62776 50232 0 _1409_
rlabel metal3 36288 56056 36288 56056 0 _1410_
rlabel metal2 39032 55496 39032 55496 0 _1411_
rlabel metal2 38808 55412 38808 55412 0 _1412_
rlabel metal2 31304 56224 31304 56224 0 _1413_
rlabel metal2 37856 56056 37856 56056 0 _1414_
rlabel metal2 38472 56728 38472 56728 0 _1415_
rlabel metal2 55720 53312 55720 53312 0 _1416_
rlabel metal2 50456 55160 50456 55160 0 _1417_
rlabel metal2 49224 55216 49224 55216 0 _1418_
rlabel metal3 49560 54880 49560 54880 0 _1419_
rlabel metal3 52472 54600 52472 54600 0 _1420_
rlabel metal2 53032 52136 53032 52136 0 _1421_
rlabel metal2 54824 50204 54824 50204 0 _1422_
rlabel metal2 53592 54432 53592 54432 0 _1423_
rlabel metal2 53480 54768 53480 54768 0 _1424_
rlabel metal3 54264 54488 54264 54488 0 _1425_
rlabel metal2 54264 52752 54264 52752 0 _1426_
rlabel metal2 54488 55944 54488 55944 0 _1427_
rlabel metal2 52080 53704 52080 53704 0 _1428_
rlabel metal2 40600 56560 40600 56560 0 _1429_
rlabel metal2 55160 55776 55160 55776 0 _1430_
rlabel metal2 53816 57680 53816 57680 0 _1431_
rlabel metal3 55944 53704 55944 53704 0 _1432_
rlabel metal2 53928 53088 53928 53088 0 _1433_
rlabel metal2 58968 54320 58968 54320 0 _1434_
rlabel metal2 53144 57456 53144 57456 0 _1435_
rlabel metal2 46872 53928 46872 53928 0 _1436_
rlabel metal2 47432 54656 47432 54656 0 _1437_
rlabel metal2 23688 27160 23688 27160 0 _1438_
rlabel metal3 35616 25480 35616 25480 0 _1439_
rlabel metal2 24808 20048 24808 20048 0 _1440_
rlabel metal2 48832 48104 48832 48104 0 _1441_
rlabel metal2 43960 53648 43960 53648 0 _1442_
rlabel metal2 45584 53704 45584 53704 0 _1443_
rlabel metal2 37352 25816 37352 25816 0 _1444_
rlabel metal2 42728 46088 42728 46088 0 _1445_
rlabel metal2 44968 52584 44968 52584 0 _1446_
rlabel metal2 48888 56952 48888 56952 0 _1447_
rlabel metal3 55496 52808 55496 52808 0 _1448_
rlabel metal2 56840 54152 56840 54152 0 _1449_
rlabel metal3 56392 52696 56392 52696 0 _1450_
rlabel metal2 41496 29736 41496 29736 0 _1451_
rlabel metal2 41832 33040 41832 33040 0 _1452_
rlabel metal2 59416 51072 59416 51072 0 _1453_
rlabel metal2 62664 49336 62664 49336 0 _1454_
rlabel metal2 61880 38808 61880 38808 0 _1455_
rlabel metal2 58520 48160 58520 48160 0 _1456_
rlabel metal2 53816 49280 53816 49280 0 _1457_
rlabel metal3 56896 47432 56896 47432 0 _1458_
rlabel metal2 57848 48552 57848 48552 0 _1459_
rlabel metal4 54264 44016 54264 44016 0 _1460_
rlabel metal3 55160 23912 55160 23912 0 _1461_
rlabel metal2 55160 25032 55160 25032 0 _1462_
rlabel metal2 55496 24976 55496 24976 0 _1463_
rlabel metal2 55272 25844 55272 25844 0 _1464_
rlabel metal2 54600 40600 54600 40600 0 _1465_
rlabel metal2 57960 39256 57960 39256 0 _1466_
rlabel metal2 58296 34776 58296 34776 0 _1467_
rlabel metal2 52808 32872 52808 32872 0 _1468_
rlabel metal2 58408 36512 58408 36512 0 _1469_
rlabel metal2 59640 34832 59640 34832 0 _1470_
rlabel metal2 60984 36400 60984 36400 0 _1471_
rlabel metal2 60648 36792 60648 36792 0 _1472_
rlabel metal2 58968 44184 58968 44184 0 _1473_
rlabel metal2 58632 41440 58632 41440 0 _1474_
rlabel metal2 61096 37352 61096 37352 0 _1475_
rlabel metal2 59080 39312 59080 39312 0 _1476_
rlabel metal2 56560 41048 56560 41048 0 _1477_
rlabel metal2 56168 41496 56168 41496 0 _1478_
rlabel metal3 58744 13048 58744 13048 0 _1479_
rlabel metal2 57400 49672 57400 49672 0 _1480_
rlabel metal2 54824 39704 54824 39704 0 _1481_
rlabel metal3 56504 41048 56504 41048 0 _1482_
rlabel metal2 57624 39564 57624 39564 0 _1483_
rlabel metal2 59640 38864 59640 38864 0 _1484_
rlabel metal2 57288 40208 57288 40208 0 _1485_
rlabel metal2 53704 45136 53704 45136 0 _1486_
rlabel metal2 54096 48440 54096 48440 0 _1487_
rlabel metal2 31080 47880 31080 47880 0 _1488_
rlabel metal2 49448 47712 49448 47712 0 _1489_
rlabel metal3 32368 49896 32368 49896 0 _1490_
rlabel metal2 23352 47096 23352 47096 0 _1491_
rlabel metal2 25816 45808 25816 45808 0 _1492_
rlabel metal2 29400 47376 29400 47376 0 _1493_
rlabel metal2 29176 47320 29176 47320 0 _1494_
rlabel metal2 29624 47152 29624 47152 0 _1495_
rlabel metal2 56392 48104 56392 48104 0 _1496_
rlabel metal2 38920 54264 38920 54264 0 _1497_
rlabel metal2 31528 48440 31528 48440 0 _1498_
rlabel metal2 35000 51632 35000 51632 0 _1499_
rlabel metal2 34776 50092 34776 50092 0 _1500_
rlabel metal2 33992 52192 33992 52192 0 _1501_
rlabel metal3 32928 51352 32928 51352 0 _1502_
rlabel metal3 29736 57624 29736 57624 0 _1503_
rlabel metal2 30632 52864 30632 52864 0 _1504_
rlabel metal2 30408 52752 30408 52752 0 _1505_
rlabel metal2 31304 50204 31304 50204 0 _1506_
rlabel metal2 32984 49896 32984 49896 0 _1507_
rlabel metal2 33432 50288 33432 50288 0 _1508_
rlabel metal2 49896 48216 49896 48216 0 _1509_
rlabel metal2 28168 47432 28168 47432 0 _1510_
rlabel metal2 30968 48272 30968 48272 0 _1511_
rlabel metal3 30296 49224 30296 49224 0 _1512_
rlabel metal3 32760 52024 32760 52024 0 _1513_
rlabel metal2 32256 52136 32256 52136 0 _1514_
rlabel metal2 36232 48216 36232 48216 0 _1515_
rlabel metal2 40264 47376 40264 47376 0 _1516_
rlabel metal3 50512 52920 50512 52920 0 _1517_
rlabel metal3 53872 51016 53872 51016 0 _1518_
rlabel metal2 52136 48916 52136 48916 0 _1519_
rlabel metal2 50792 49392 50792 49392 0 _1520_
rlabel metal2 52024 53200 52024 53200 0 _1521_
rlabel metal2 50344 50792 50344 50792 0 _1522_
rlabel metal2 47768 49056 47768 49056 0 _1523_
rlabel metal2 45864 47376 45864 47376 0 _1524_
rlabel metal2 56616 21672 56616 21672 0 _1525_
rlabel metal2 56392 20832 56392 20832 0 _1526_
rlabel metal2 56056 33040 56056 33040 0 _1527_
rlabel metal2 45640 47544 45640 47544 0 _1528_
rlabel metal2 39872 51576 39872 51576 0 _1529_
rlabel metal2 39592 49308 39592 49308 0 _1530_
rlabel metal2 39256 52808 39256 52808 0 _1531_
rlabel metal2 41048 49336 41048 49336 0 _1532_
rlabel metal3 41832 49784 41832 49784 0 _1533_
rlabel metal2 41160 49784 41160 49784 0 _1534_
rlabel metal2 47096 46984 47096 46984 0 _1535_
rlabel metal2 45976 49056 45976 49056 0 _1536_
rlabel metal3 55944 50008 55944 50008 0 _1537_
rlabel metal2 48776 47432 48776 47432 0 _1538_
rlabel metal3 47432 45864 47432 45864 0 _1539_
rlabel metal2 44408 43848 44408 43848 0 _1540_
rlabel metal2 47992 46816 47992 46816 0 _1541_
rlabel metal2 46648 46984 46648 46984 0 _1542_
rlabel metal2 46760 47376 46760 47376 0 _1543_
rlabel metal2 46984 49392 46984 49392 0 _1544_
rlabel metal3 45024 48216 45024 48216 0 _1545_
rlabel metal3 46760 49000 46760 49000 0 _1546_
rlabel metal2 49000 49336 49000 49336 0 _1547_
rlabel metal2 43624 47712 43624 47712 0 _1548_
rlabel metal2 44184 48944 44184 48944 0 _1549_
rlabel metal2 47768 48160 47768 48160 0 _1550_
rlabel metal3 47936 47432 47936 47432 0 _1551_
rlabel metal3 45864 46760 45864 46760 0 _1552_
rlabel metal2 46088 48496 46088 48496 0 _1553_
rlabel metal2 49784 49952 49784 49952 0 _1554_
rlabel metal2 50904 49336 50904 49336 0 _1555_
rlabel metal2 51744 47656 51744 47656 0 _1556_
rlabel metal2 49784 50428 49784 50428 0 _1557_
rlabel metal2 50792 50960 50792 50960 0 _1558_
rlabel metal2 49224 50456 49224 50456 0 _1559_
rlabel metal2 51464 50176 51464 50176 0 _1560_
rlabel metal2 43008 49112 43008 49112 0 _1561_
rlabel metal2 43008 47544 43008 47544 0 _1562_
rlabel metal2 42224 50344 42224 50344 0 _1563_
rlabel metal2 45304 31640 45304 31640 0 _1564_
rlabel metal2 42840 46872 42840 46872 0 _1565_
rlabel metal2 42280 47712 42280 47712 0 _1566_
rlabel metal2 62216 42616 62216 42616 0 _1567_
rlabel metal2 47544 37464 47544 37464 0 _1568_
rlabel metal2 46872 40544 46872 40544 0 _1569_
rlabel metal3 48664 39480 48664 39480 0 _1570_
rlabel metal2 48776 39816 48776 39816 0 _1571_
rlabel metal2 51800 39144 51800 39144 0 _1572_
rlabel metal2 52920 11088 52920 11088 0 _1573_
rlabel metal2 52696 11032 52696 11032 0 _1574_
rlabel metal2 50904 10528 50904 10528 0 _1575_
rlabel metal2 50568 11872 50568 11872 0 _1576_
rlabel metal3 61824 40376 61824 40376 0 _1577_
rlabel metal2 49448 39144 49448 39144 0 _1578_
rlabel metal2 51912 34888 51912 34888 0 _1579_
rlabel metal2 47768 34608 47768 34608 0 _1580_
rlabel metal2 43736 37576 43736 37576 0 _1581_
rlabel metal2 46256 34888 46256 34888 0 _1582_
rlabel metal2 45024 36456 45024 36456 0 _1583_
rlabel metal2 48216 34608 48216 34608 0 _1584_
rlabel metal2 51016 35168 51016 35168 0 _1585_
rlabel metal2 56056 35168 56056 35168 0 _1586_
rlabel metal2 50456 34608 50456 34608 0 _1587_
rlabel metal4 45192 35560 45192 35560 0 _1588_
rlabel metal2 50120 35224 50120 35224 0 _1589_
rlabel metal3 48608 33880 48608 33880 0 _1590_
rlabel metal2 52248 34216 52248 34216 0 _1591_
rlabel metal2 50344 38808 50344 38808 0 _1592_
rlabel metal2 42840 40712 42840 40712 0 _1593_
rlabel metal2 48104 37968 48104 37968 0 _1594_
rlabel metal3 47656 37352 47656 37352 0 _1595_
rlabel metal2 49112 35728 49112 35728 0 _1596_
rlabel metal2 48720 36456 48720 36456 0 _1597_
rlabel metal2 48776 36848 48776 36848 0 _1598_
rlabel metal3 48216 38920 48216 38920 0 _1599_
rlabel metal3 47936 45192 47936 45192 0 _1600_
rlabel metal2 20664 43456 20664 43456 0 _1601_
rlabel metal2 22008 46256 22008 46256 0 _1602_
rlabel metal2 16632 47544 16632 47544 0 _1603_
rlabel metal2 20552 44800 20552 44800 0 _1604_
rlabel metal3 21896 45080 21896 45080 0 _1605_
rlabel metal2 21784 45920 21784 45920 0 _1606_
rlabel metal3 20328 46760 20328 46760 0 _1607_
rlabel metal2 47320 41664 47320 41664 0 _1608_
rlabel metal3 19824 46536 19824 46536 0 _1609_
rlabel metal2 19880 47880 19880 47880 0 _1610_
rlabel metal2 12824 47880 12824 47880 0 _1611_
rlabel metal2 14280 48608 14280 48608 0 _1612_
rlabel metal2 13608 47880 13608 47880 0 _1613_
rlabel metal2 15400 48888 15400 48888 0 _1614_
rlabel metal2 14840 49280 14840 49280 0 _1615_
rlabel metal2 34216 51240 34216 51240 0 _1616_
rlabel metal2 19768 49224 19768 49224 0 _1617_
rlabel metal2 18536 49280 18536 49280 0 _1618_
rlabel metal2 18144 48216 18144 48216 0 _1619_
rlabel metal2 21336 49448 21336 49448 0 _1620_
rlabel metal2 17304 49560 17304 49560 0 _1621_
rlabel metal2 17416 45416 17416 45416 0 _1622_
rlabel metal2 17640 37688 17640 37688 0 _1623_
rlabel metal2 19768 46816 19768 46816 0 _1624_
rlabel metal2 21448 46872 21448 46872 0 _1625_
rlabel metal2 16744 48384 16744 48384 0 _1626_
rlabel metal3 17976 49000 17976 49000 0 _1627_
rlabel metal2 17976 48216 17976 48216 0 _1628_
rlabel metal2 44408 46984 44408 46984 0 _1629_
rlabel metal2 44744 44632 44744 44632 0 _1630_
rlabel metal3 46144 45080 46144 45080 0 _1631_
rlabel metal3 45752 42168 45752 42168 0 _1632_
rlabel metal2 44072 45192 44072 45192 0 _1633_
rlabel metal2 48104 49896 48104 49896 0 _1634_
rlabel metal3 45640 47768 45640 47768 0 _1635_
rlabel metal3 43008 41944 43008 41944 0 _1636_
rlabel metal3 39872 46760 39872 46760 0 _1637_
rlabel metal2 53704 8848 53704 8848 0 _1638_
rlabel metal2 58856 14000 58856 14000 0 _1639_
rlabel metal2 42392 30184 42392 30184 0 _1640_
rlabel metal2 42168 42952 42168 42952 0 _1641_
rlabel metal3 15148 45864 15148 45864 0 _1642_
rlabel metal2 14728 44520 14728 44520 0 _1643_
rlabel metal2 13608 45584 13608 45584 0 _1644_
rlabel metal3 11368 43512 11368 43512 0 _1645_
rlabel metal2 14168 43624 14168 43624 0 _1646_
rlabel metal2 41384 44632 41384 44632 0 _1647_
rlabel metal3 40600 44408 40600 44408 0 _1648_
rlabel metal2 48328 44968 48328 44968 0 _1649_
rlabel metal2 40376 45136 40376 45136 0 _1650_
rlabel metal3 34328 45304 34328 45304 0 _1651_
rlabel metal2 33768 46312 33768 46312 0 _1652_
rlabel metal2 39368 45024 39368 45024 0 _1653_
rlabel metal2 39424 41272 39424 41272 0 _1654_
rlabel metal2 38752 41384 38752 41384 0 _1655_
rlabel metal2 40824 43120 40824 43120 0 _1656_
rlabel metal2 16296 44800 16296 44800 0 _1657_
rlabel metal3 34160 45192 34160 45192 0 _1658_
rlabel metal2 41160 43288 41160 43288 0 _1659_
rlabel metal3 43960 44632 43960 44632 0 _1660_
rlabel metal2 36568 44856 36568 44856 0 _1661_
rlabel metal2 40936 42784 40936 42784 0 _1662_
rlabel metal2 42952 42504 42952 42504 0 _1663_
rlabel metal2 44296 43624 44296 43624 0 _1664_
rlabel metal2 44072 41944 44072 41944 0 _1665_
rlabel metal3 44072 44296 44072 44296 0 _1666_
rlabel metal2 43400 44856 43400 44856 0 _1667_
rlabel metal2 42504 44520 42504 44520 0 _1668_
rlabel metal2 39704 44744 39704 44744 0 _1669_
rlabel metal2 38024 44296 38024 44296 0 _1670_
rlabel metal2 40264 45360 40264 45360 0 _1671_
rlabel metal2 41160 45136 41160 45136 0 _1672_
rlabel metal2 39816 36064 39816 36064 0 _1673_
rlabel metal2 33768 42112 33768 42112 0 _1674_
rlabel metal2 36008 39144 36008 39144 0 _1675_
rlabel metal2 32760 41328 32760 41328 0 _1676_
rlabel metal2 37464 40656 37464 40656 0 _1677_
rlabel metal2 37072 39816 37072 39816 0 _1678_
rlabel metal3 36568 11480 36568 11480 0 _1679_
rlabel metal3 36680 9800 36680 9800 0 _1680_
rlabel metal2 36960 9576 36960 9576 0 _1681_
rlabel metal2 37688 11592 37688 11592 0 _1682_
rlabel metal2 43568 34328 43568 34328 0 _1683_
rlabel metal2 36456 38724 36456 38724 0 _1684_
rlabel metal2 36680 35952 36680 35952 0 _1685_
rlabel metal2 39704 32816 39704 32816 0 _1686_
rlabel metal2 39816 33040 39816 33040 0 _1687_
rlabel metal2 38696 36512 38696 36512 0 _1688_
rlabel metal2 45416 35952 45416 35952 0 _1689_
rlabel metal3 42728 35784 42728 35784 0 _1690_
rlabel metal2 41384 33656 41384 33656 0 _1691_
rlabel metal2 37464 36064 37464 36064 0 _1692_
rlabel metal3 40880 38920 40880 38920 0 _1693_
rlabel metal2 36344 36456 36344 36456 0 _1694_
rlabel metal3 45360 9240 45360 9240 0 _1695_
rlabel metal2 37464 37968 37464 37968 0 _1696_
rlabel metal2 39704 37184 39704 37184 0 _1697_
rlabel metal2 40600 34160 40600 34160 0 _1698_
rlabel metal2 41048 35448 41048 35448 0 _1699_
rlabel metal2 40656 35112 40656 35112 0 _1700_
rlabel metal2 33544 39928 33544 39928 0 _1701_
rlabel metal2 31864 42392 31864 42392 0 _1702_
rlabel metal2 7112 41720 7112 41720 0 _1703_
rlabel metal3 21336 43120 21336 43120 0 _1704_
rlabel metal2 5768 42728 5768 42728 0 _1705_
rlabel metal3 7392 39592 7392 39592 0 _1706_
rlabel metal2 10024 38752 10024 38752 0 _1707_
rlabel metal2 10360 38024 10360 38024 0 _1708_
rlabel metal2 8848 39032 8848 39032 0 _1709_
rlabel metal2 10024 39032 10024 39032 0 _1710_
rlabel metal2 33824 40936 33824 40936 0 _1711_
rlabel metal3 10080 41160 10080 41160 0 _1712_
rlabel metal2 8680 43624 8680 43624 0 _1713_
rlabel metal2 6216 47768 6216 47768 0 _1714_
rlabel metal2 2632 46144 2632 46144 0 _1715_
rlabel metal3 11256 50344 11256 50344 0 _1716_
rlabel metal2 7448 46760 7448 46760 0 _1717_
rlabel metal2 7336 46760 7336 46760 0 _1718_
rlabel metal2 7672 44968 7672 44968 0 _1719_
rlabel metal3 5376 47208 5376 47208 0 _1720_
rlabel metal3 8288 42728 8288 42728 0 _1721_
rlabel metal3 2520 41944 2520 41944 0 _1722_
rlabel metal2 8008 42168 8008 42168 0 _1723_
rlabel metal2 8120 43624 8120 43624 0 _1724_
rlabel metal2 6328 42504 6328 42504 0 _1725_
rlabel metal2 6664 45976 6664 45976 0 _1726_
rlabel metal2 8344 44352 8344 44352 0 _1727_
rlabel metal3 7672 45080 7672 45080 0 _1728_
rlabel metal3 7840 43512 7840 43512 0 _1729_
rlabel metal2 20552 43232 20552 43232 0 _1730_
rlabel metal3 28616 43512 28616 43512 0 _1731_
rlabel metal2 32088 43120 32088 43120 0 _1732_
rlabel metal2 31696 42840 31696 42840 0 _1733_
rlabel metal2 30632 43568 30632 43568 0 _1734_
rlabel metal2 41552 43288 41552 43288 0 _1735_
rlabel metal2 31360 42056 31360 42056 0 _1736_
rlabel metal2 30968 40544 30968 40544 0 _1737_
rlabel metal2 30968 42224 30968 42224 0 _1738_
rlabel metal2 31304 42896 31304 42896 0 _1739_
rlabel metal2 29848 43288 29848 43288 0 _1740_
rlabel metal2 30072 43232 30072 43232 0 _1741_
rlabel metal2 19880 38724 19880 38724 0 _1742_
rlabel metal3 16240 49672 16240 49672 0 _1743_
rlabel metal2 29232 42952 29232 42952 0 _1744_
rlabel metal2 22400 49672 22400 49672 0 _1745_
rlabel metal3 2996 17080 2996 17080 0 _1746_
rlabel metal3 1512 17752 1512 17752 0 _1747_
rlabel metal2 26992 37016 26992 37016 0 _1748_
rlabel metal3 28280 40600 28280 40600 0 _1749_
rlabel metal2 26600 38024 26600 38024 0 _1750_
rlabel metal3 16296 53032 16296 53032 0 _1751_
rlabel metal2 24472 57456 24472 57456 0 _1752_
rlabel metal2 24584 58352 24584 58352 0 _1753_
rlabel metal2 30520 56392 30520 56392 0 _1754_
rlabel metal3 26348 53144 26348 53144 0 _1755_
rlabel metal2 22736 18424 22736 18424 0 _1756_
rlabel metal2 3304 42280 3304 42280 0 _1757_
rlabel metal2 26488 53200 26488 53200 0 _1758_
rlabel metal2 24360 59528 24360 59528 0 _1759_
rlabel metal2 25256 56560 25256 56560 0 _1760_
rlabel metal3 24920 56168 24920 56168 0 _1761_
rlabel metal2 21392 56952 21392 56952 0 _1762_
rlabel metal3 32928 55272 32928 55272 0 _1763_
rlabel metal2 58744 49504 58744 49504 0 _1764_
rlabel metal2 56056 55720 56056 55720 0 _1765_
rlabel metal2 58296 49280 58296 49280 0 _1766_
rlabel metal2 58408 54376 58408 54376 0 _1767_
rlabel metal3 39984 55944 39984 55944 0 _1768_
rlabel metal2 33656 56504 33656 56504 0 _1769_
rlabel metal2 24248 55216 24248 55216 0 _1770_
rlabel metal2 22568 54208 22568 54208 0 _1771_
rlabel metal2 26264 32200 26264 32200 0 _1772_
rlabel metal2 1624 44352 1624 44352 0 _1773_
rlabel metal2 25760 49784 25760 49784 0 _1774_
rlabel metal2 25816 32312 25816 32312 0 _1775_
rlabel metal2 25200 49784 25200 49784 0 _1776_
rlabel metal3 25144 50008 25144 50008 0 _1777_
rlabel metal2 36288 54712 36288 54712 0 _1778_
rlabel metal2 25144 54096 25144 54096 0 _1779_
rlabel metal2 24584 52864 24584 52864 0 _1780_
rlabel metal2 23408 52248 23408 52248 0 _1781_
rlabel metal2 22792 49392 22792 49392 0 _1782_
rlabel metal2 24136 48328 24136 48328 0 _1783_
rlabel metal2 21448 50064 21448 50064 0 _1784_
rlabel metal3 21224 50456 21224 50456 0 _1785_
rlabel metal2 20888 54936 20888 54936 0 _1786_
rlabel metal3 17248 56056 17248 56056 0 _1787_
rlabel metal2 17528 56728 17528 56728 0 _1788_
rlabel metal2 22176 54488 22176 54488 0 _1789_
rlabel metal2 21840 50232 21840 50232 0 _1790_
rlabel metal2 23072 52360 23072 52360 0 _1791_
rlabel metal3 19376 54488 19376 54488 0 _1792_
rlabel metal2 24360 55160 24360 55160 0 _1793_
rlabel metal2 23912 54936 23912 54936 0 _1794_
rlabel metal2 24360 51464 24360 51464 0 _1795_
rlabel metal2 21896 55720 21896 55720 0 _1796_
rlabel metal2 22568 49896 22568 49896 0 _1797_
rlabel metal2 17472 52808 17472 52808 0 _1798_
rlabel metal2 19096 53200 19096 53200 0 _1799_
rlabel metal2 26600 54600 26600 54600 0 _1800_
rlabel metal2 37968 31752 37968 31752 0 g.bi_l\[0\]\[0\]
rlabel metal2 35112 33096 35112 33096 0 g.bi_l\[0\]\[1\]
rlabel metal2 52920 14280 52920 14280 0 g.bi_l\[11\]\[0\]
rlabel metal2 55048 12656 55048 12656 0 g.bi_l\[11\]\[1\]
rlabel metal2 62216 21448 62216 21448 0 g.bi_l\[13\]\[0\]
rlabel metal3 60816 24136 60816 24136 0 g.bi_l\[13\]\[1\]
rlabel metal3 47656 29288 47656 29288 0 g.bi_l\[15\]\[0\]
rlabel metal2 49896 29176 49896 29176 0 g.bi_l\[15\]\[1\]
rlabel metal2 24696 8512 24696 8512 0 g.bi_l\[16\]\[0\]
rlabel metal2 27608 6496 27608 6496 0 g.bi_l\[16\]\[1\]
rlabel metal2 44856 6216 44856 6216 0 g.bi_l\[18\]\[0\]
rlabel metal2 44968 5880 44968 5880 0 g.bi_l\[18\]\[1\]
rlabel metal3 45136 17864 45136 17864 0 g.bi_l\[20\]\[0\]
rlabel metal2 42056 20104 42056 20104 0 g.bi_l\[20\]\[1\]
rlabel metal2 42952 26544 42952 26544 0 g.bi_l\[22\]\[0\]
rlabel metal2 46760 24304 46760 24304 0 g.bi_l\[22\]\[1\]
rlabel metal2 13832 10024 13832 10024 0 g.bi_l\[25\]\[0\]
rlabel metal3 11760 8232 11760 8232 0 g.bi_l\[25\]\[1\]
rlabel metal3 23688 15176 23688 15176 0 g.bi_l\[27\]\[0\]
rlabel metal2 21560 14504 21560 14504 0 g.bi_l\[27\]\[1\]
rlabel metal3 32872 26264 32872 26264 0 g.bi_l\[29\]\[0\]
rlabel metal2 35168 24136 35168 24136 0 g.bi_l\[29\]\[1\]
rlabel metal3 43456 36456 43456 36456 0 g.bi_l\[2\]\[0\]
rlabel metal3 44968 33320 44968 33320 0 g.bi_l\[2\]\[1\]
rlabel metal2 21336 24752 21336 24752 0 g.bi_l\[31\]\[0\]
rlabel metal3 19992 25704 19992 25704 0 g.bi_l\[31\]\[1\]
rlabel metal2 2632 23576 2632 23576 0 g.bi_l\[32\]\[0\]
rlabel metal2 4816 26040 4816 26040 0 g.bi_l\[32\]\[1\]
rlabel metal2 15960 16128 15960 16128 0 g.bi_l\[34\]\[0\]
rlabel metal2 12992 17528 12992 17528 0 g.bi_l\[34\]\[1\]
rlabel metal2 16464 25704 16464 25704 0 g.bi_l\[36\]\[0\]
rlabel metal2 12488 27272 12488 27272 0 g.bi_l\[36\]\[1\]
rlabel metal2 20776 33208 20776 33208 0 g.bi_l\[38\]\[0\]
rlabel metal2 21448 34720 21448 34720 0 g.bi_l\[38\]\[1\]
rlabel metal2 8344 38668 8344 38668 0 g.bi_l\[41\]\[0\]
rlabel metal2 7448 36512 7448 36512 0 g.bi_l\[41\]\[1\]
rlabel metal2 16240 40264 16240 40264 0 g.bi_l\[43\]\[0\]
rlabel metal2 19208 40880 19208 40880 0 g.bi_l\[43\]\[1\]
rlabel metal2 23800 48272 23800 48272 0 g.bi_l\[45\]\[0\]
rlabel metal2 26096 47320 26096 47320 0 g.bi_l\[45\]\[1\]
rlabel metal2 16632 56560 16632 56560 0 g.bi_l\[47\]\[0\]
rlabel metal2 16464 57624 16464 57624 0 g.bi_l\[47\]\[1\]
rlabel metal3 5096 49112 5096 49112 0 g.bi_l\[48\]\[0\]
rlabel metal2 3192 41216 3192 41216 0 g.bi_l\[48\]\[1\]
rlabel metal2 55496 35504 55496 35504 0 g.bi_l\[4\]\[0\]
rlabel metal2 58800 33880 58800 33880 0 g.bi_l\[4\]\[1\]
rlabel metal3 10192 49112 10192 49112 0 g.bi_l\[50\]\[0\]
rlabel metal3 13720 50568 13720 50568 0 g.bi_l\[50\]\[1\]
rlabel metal2 40040 49784 40040 49784 0 g.bi_l\[52\]\[0\]
rlabel metal2 38416 50008 38416 50008 0 g.bi_l\[52\]\[1\]
rlabel metal2 32760 57064 32760 57064 0 g.bi_l\[54\]\[0\]
rlabel metal2 33544 58856 33544 58856 0 g.bi_l\[54\]\[1\]
rlabel metal3 36120 41160 36120 41160 0 g.bi_l\[57\]\[0\]
rlabel metal2 35168 42168 35168 42168 0 g.bi_l\[57\]\[1\]
rlabel metal2 46816 41944 46816 41944 0 g.bi_l\[59\]\[0\]
rlabel metal2 44968 41552 44968 41552 0 g.bi_l\[59\]\[1\]
rlabel metal3 54096 50008 54096 50008 0 g.bi_l\[61\]\[0\]
rlabel metal2 54040 49000 54040 49000 0 g.bi_l\[61\]\[1\]
rlabel metal2 49392 54376 49392 54376 0 g.bi_l\[63\]\[0\]
rlabel metal2 45304 55776 45304 55776 0 g.bi_l\[63\]\[1\]
rlabel metal2 61768 17640 61768 17640 0 g.bi_l\[6\]\[0\]
rlabel metal3 61320 47544 61320 47544 0 g.bi_l\[6\]\[1\]
rlabel metal2 37016 11872 37016 11872 0 g.bi_l\[9\]\[0\]
rlabel metal2 39704 12264 39704 12264 0 g.bi_l\[9\]\[1\]
rlabel metal2 37128 31136 37128 31136 0 g.g_y\[0\].g_x\[0\].t.out_sc
rlabel metal2 32312 31248 32312 31248 0 g.g_y\[0\].g_x\[0\].t.r_d
rlabel metal3 36848 31640 36848 31640 0 g.g_y\[0\].g_x\[0\].t.r_h
rlabel metal2 31864 32928 31864 32928 0 g.g_y\[0\].g_x\[0\].t.r_v
rlabel metal2 36232 33040 36232 33040 0 g.g_y\[0\].g_x\[0\].t.w_dh
rlabel metal2 33432 34272 33432 34272 0 g.g_y\[0\].g_x\[0\].t.w_na
rlabel metal2 34328 30408 34328 30408 0 g.g_y\[0\].g_x\[0\].t.w_si
rlabel metal2 40040 39760 40040 39760 0 g.g_y\[0\].g_x\[1\].t.out_sc
rlabel metal2 41552 36456 41552 36456 0 g.g_y\[0\].g_x\[1\].t.r_d
rlabel metal2 42840 34384 42840 34384 0 g.g_y\[0\].g_x\[1\].t.r_h
rlabel metal3 36680 40488 36680 40488 0 g.g_y\[0\].g_x\[1\].t.r_v
rlabel metal2 37912 38360 37912 38360 0 g.g_y\[0\].g_x\[1\].t.w_si
rlabel metal3 46424 38808 46424 38808 0 g.g_y\[0\].g_x\[2\].t.out_sc
rlabel metal2 45976 31416 45976 31416 0 g.g_y\[0\].g_x\[2\].t.r_d
rlabel metal3 45696 34104 45696 34104 0 g.g_y\[0\].g_x\[2\].t.r_h
rlabel metal3 44184 31864 44184 31864 0 g.g_y\[0\].g_x\[2\].t.r_v
rlabel metal2 43960 37240 43960 37240 0 g.g_y\[0\].g_x\[2\].t.w_dh
rlabel metal2 42280 33600 42280 33600 0 g.g_y\[0\].g_x\[2\].t.w_na
rlabel metal3 42112 38696 42112 38696 0 g.g_y\[0\].g_x\[2\].t.w_si
rlabel metal3 48440 33208 48440 33208 0 g.g_y\[0\].g_x\[3\].t.out_sc
rlabel metal2 51016 33544 51016 33544 0 g.g_y\[0\].g_x\[3\].t.r_d
rlabel metal3 51464 33320 51464 33320 0 g.g_y\[0\].g_x\[3\].t.r_h
rlabel metal2 46424 37296 46424 37296 0 g.g_y\[0\].g_x\[3\].t.r_v
rlabel metal2 46648 38668 46648 38668 0 g.g_y\[0\].g_x\[3\].t.w_si
rlabel metal3 58128 32424 58128 32424 0 g.g_y\[0\].g_x\[4\].t.out_sc
rlabel metal3 59472 33320 59472 33320 0 g.g_y\[0\].g_x\[4\].t.r_d
rlabel metal3 58352 33880 58352 33880 0 g.g_y\[0\].g_x\[4\].t.r_h
rlabel metal2 55720 32088 55720 32088 0 g.g_y\[0\].g_x\[4\].t.r_v
rlabel metal2 55384 32760 55384 32760 0 g.g_y\[0\].g_x\[4\].t.w_dh
rlabel metal2 57064 34384 57064 34384 0 g.g_y\[0\].g_x\[4\].t.w_na
rlabel metal2 52024 33320 52024 33320 0 g.g_y\[0\].g_x\[4\].t.w_si
rlabel metal2 62216 38192 62216 38192 0 g.g_y\[0\].g_x\[5\].t.out_sc
rlabel metal3 58352 38808 58352 38808 0 g.g_y\[0\].g_x\[5\].t.r_d
rlabel metal2 58072 42168 58072 42168 0 g.g_y\[0\].g_x\[5\].t.r_h
rlabel metal2 55384 41160 55384 41160 0 g.g_y\[0\].g_x\[5\].t.r_v
rlabel metal2 59584 35784 59584 35784 0 g.g_y\[0\].g_x\[5\].t.w_si
rlabel metal2 61936 46872 61936 46872 0 g.g_y\[0\].g_x\[6\].t.out_sc
rlabel metal2 61376 48104 61376 48104 0 g.g_y\[0\].g_x\[6\].t.r_d
rlabel metal2 59808 44520 59808 44520 0 g.g_y\[0\].g_x\[6\].t.r_h
rlabel metal2 62440 37744 62440 37744 0 g.g_y\[0\].g_x\[6\].t.r_v
rlabel metal2 56952 45248 56952 45248 0 g.g_y\[0\].g_x\[6\].t.w_dh
rlabel metal2 59640 47152 59640 47152 0 g.g_y\[0\].g_x\[6\].t.w_na
rlabel metal2 61096 41552 61096 41552 0 g.g_y\[0\].g_x\[6\].t.w_si
rlabel metal2 50344 39984 50344 39984 0 g.g_y\[0\].g_x\[7\].t.out_sc
rlabel metal2 52024 41552 52024 41552 0 g.g_y\[0\].g_x\[7\].t.r_d
rlabel metal3 54376 47768 54376 47768 0 g.g_y\[0\].g_x\[7\].t.r_h
rlabel metal2 49448 46816 49448 46816 0 g.g_y\[0\].g_x\[7\].t.r_v
rlabel metal2 52472 40544 52472 40544 0 g.g_y\[0\].g_x\[7\].t.w_si
rlabel metal2 30800 15512 30800 15512 0 g.g_y\[1\].g_x\[0\].t.out_sc
rlabel metal2 28112 16184 28112 16184 0 g.g_y\[1\].g_x\[0\].t.r_d
rlabel metal2 31920 16072 31920 16072 0 g.g_y\[1\].g_x\[0\].t.r_h
rlabel metal2 26376 11928 26376 11928 0 g.g_y\[1\].g_x\[0\].t.r_v
rlabel metal2 27888 15512 27888 15512 0 g.g_y\[1\].g_x\[0\].t.w_si
rlabel metal2 38808 11144 38808 11144 0 g.g_y\[1\].g_x\[1\].t.out_sc
rlabel metal2 37632 12824 37632 12824 0 g.g_y\[1\].g_x\[1\].t.r_d
rlabel metal3 37912 15512 37912 15512 0 g.g_y\[1\].g_x\[1\].t.r_h
rlabel metal2 36792 10976 36792 10976 0 g.g_y\[1\].g_x\[1\].t.r_v
rlabel metal2 35672 15400 35672 15400 0 g.g_y\[1\].g_x\[1\].t.w_dh
rlabel metal2 33432 11872 33432 11872 0 g.g_y\[1\].g_x\[1\].t.w_na
rlabel metal2 34384 15512 34384 15512 0 g.g_y\[1\].g_x\[1\].t.w_si
rlabel metal3 44016 16184 44016 16184 0 g.g_y\[1\].g_x\[2\].t.out_sc
rlabel metal3 43568 14728 43568 14728 0 g.g_y\[1\].g_x\[2\].t.r_d
rlabel metal3 48328 15400 48328 15400 0 g.g_y\[1\].g_x\[2\].t.r_h
rlabel metal3 44800 12152 44800 12152 0 g.g_y\[1\].g_x\[2\].t.r_v
rlabel metal2 39368 16240 39368 16240 0 g.g_y\[1\].g_x\[2\].t.w_si
rlabel metal2 57008 12264 57008 12264 0 g.g_y\[1\].g_x\[3\].t.out_sc
rlabel metal2 55272 12880 55272 12880 0 g.g_y\[1\].g_x\[3\].t.r_d
rlabel metal3 54600 15176 54600 15176 0 g.g_y\[1\].g_x\[3\].t.r_h
rlabel metal2 51800 12152 51800 12152 0 g.g_y\[1\].g_x\[3\].t.r_v
rlabel metal2 49784 14168 49784 14168 0 g.g_y\[1\].g_x\[3\].t.w_dh
rlabel metal2 53368 12488 53368 12488 0 g.g_y\[1\].g_x\[3\].t.w_na
rlabel metal2 50848 16184 50848 16184 0 g.g_y\[1\].g_x\[3\].t.w_si
rlabel metal2 59976 18816 59976 18816 0 g.g_y\[1\].g_x\[4\].t.out_sc
rlabel metal2 58744 14868 58744 14868 0 g.g_y\[1\].g_x\[4\].t.r_d
rlabel metal2 57624 16016 57624 16016 0 g.g_y\[1\].g_x\[4\].t.r_h
rlabel metal2 57176 17528 57176 17528 0 g.g_y\[1\].g_x\[4\].t.r_v
rlabel metal2 57624 14868 57624 14868 0 g.g_y\[1\].g_x\[4\].t.w_si
rlabel metal2 61208 17752 61208 17752 0 g.g_y\[1\].g_x\[5\].t.out_sc
rlabel metal3 60536 21336 60536 21336 0 g.g_y\[1\].g_x\[5\].t.r_d
rlabel metal2 62048 21000 62048 21000 0 g.g_y\[1\].g_x\[5\].t.r_h
rlabel metal2 55888 21560 55888 21560 0 g.g_y\[1\].g_x\[5\].t.r_v
rlabel metal2 54264 21224 54264 21224 0 g.g_y\[1\].g_x\[5\].t.w_dh
rlabel metal2 58184 23912 58184 23912 0 g.g_y\[1\].g_x\[5\].t.w_na
rlabel metal2 59024 20104 59024 20104 0 g.g_y\[1\].g_x\[5\].t.w_si
rlabel metal2 62272 24584 62272 24584 0 g.g_y\[1\].g_x\[6\].t.out_sc
rlabel metal3 60760 28616 60760 28616 0 g.g_y\[1\].g_x\[6\].t.r_d
rlabel metal2 60200 27328 60200 27328 0 g.g_y\[1\].g_x\[6\].t.r_h
rlabel metal2 56616 31192 56616 31192 0 g.g_y\[1\].g_x\[6\].t.r_v
rlabel metal3 60368 28840 60368 28840 0 g.g_y\[1\].g_x\[6\].t.w_si
rlabel metal2 53816 26516 53816 26516 0 g.g_y\[1\].g_x\[7\].t.out_sc
rlabel metal2 48888 28728 48888 28728 0 g.g_y\[1\].g_x\[7\].t.r_d
rlabel metal3 53872 30184 53872 30184 0 g.g_y\[1\].g_x\[7\].t.r_h
rlabel metal2 47208 29568 47208 29568 0 g.g_y\[1\].g_x\[7\].t.r_v
rlabel metal2 50344 28336 50344 28336 0 g.g_y\[1\].g_x\[7\].t.w_dh
rlabel metal2 47992 29680 47992 29680 0 g.g_y\[1\].g_x\[7\].t.w_na
rlabel metal2 51688 26628 51688 26628 0 g.g_y\[1\].g_x\[7\].t.w_si
rlabel metal2 28280 5712 28280 5712 0 g.g_y\[2\].g_x\[0\].t.out_sc
rlabel metal2 27776 5880 27776 5880 0 g.g_y\[2\].g_x\[0\].t.r_d
rlabel metal2 31640 5376 31640 5376 0 g.g_y\[2\].g_x\[0\].t.r_h
rlabel metal2 24472 8512 24472 8512 0 g.g_y\[2\].g_x\[0\].t.r_v
rlabel metal2 29624 5320 29624 5320 0 g.g_y\[2\].g_x\[0\].t.w_dh
rlabel metal2 25984 7560 25984 7560 0 g.g_y\[2\].g_x\[0\].t.w_na
rlabel metal2 29904 8344 29904 8344 0 g.g_y\[2\].g_x\[0\].t.w_si
rlabel metal2 39368 6552 39368 6552 0 g.g_y\[2\].g_x\[1\].t.out_sc
rlabel metal2 36904 5544 36904 5544 0 g.g_y\[2\].g_x\[1\].t.r_d
rlabel metal2 38920 8456 38920 8456 0 g.g_y\[2\].g_x\[1\].t.r_h
rlabel metal2 33432 8708 33432 8708 0 g.g_y\[2\].g_x\[1\].t.r_v
rlabel metal2 39144 5488 39144 5488 0 g.g_y\[2\].g_x\[1\].t.w_si
rlabel metal2 42728 3976 42728 3976 0 g.g_y\[2\].g_x\[2\].t.out_sc
rlabel metal2 42336 9016 42336 9016 0 g.g_y\[2\].g_x\[2\].t.r_d
rlabel metal2 40600 5992 40600 5992 0 g.g_y\[2\].g_x\[2\].t.r_h
rlabel metal3 40600 7224 40600 7224 0 g.g_y\[2\].g_x\[2\].t.r_v
rlabel metal2 41776 6552 41776 6552 0 g.g_y\[2\].g_x\[2\].t.w_dh
rlabel metal2 43344 5992 43344 5992 0 g.g_y\[2\].g_x\[2\].t.w_na
rlabel metal2 40544 3640 40544 3640 0 g.g_y\[2\].g_x\[2\].t.w_si
rlabel metal2 50344 7336 50344 7336 0 g.g_y\[2\].g_x\[3\].t.out_sc
rlabel metal3 48552 7336 48552 7336 0 g.g_y\[2\].g_x\[3\].t.r_d
rlabel metal2 45192 11032 45192 11032 0 g.g_y\[2\].g_x\[3\].t.r_h
rlabel metal2 51464 8372 51464 8372 0 g.g_y\[2\].g_x\[3\].t.r_v
rlabel metal2 47488 5208 47488 5208 0 g.g_y\[2\].g_x\[3\].t.w_si
rlabel metal2 40376 18928 40376 18928 0 g.g_y\[2\].g_x\[4\].t.out_sc
rlabel metal2 43008 20216 43008 20216 0 g.g_y\[2\].g_x\[4\].t.r_d
rlabel metal3 46312 19992 46312 19992 0 g.g_y\[2\].g_x\[4\].t.r_h
rlabel metal2 38248 17136 38248 17136 0 g.g_y\[2\].g_x\[4\].t.r_v
rlabel metal2 47208 18424 47208 18424 0 g.g_y\[2\].g_x\[4\].t.w_dh
rlabel metal2 40264 19208 40264 19208 0 g.g_y\[2\].g_x\[4\].t.w_na
rlabel metal2 39592 18088 39592 18088 0 g.g_y\[2\].g_x\[4\].t.w_si
rlabel metal2 51072 20664 51072 20664 0 g.g_y\[2\].g_x\[5\].t.out_sc
rlabel metal2 51688 20160 51688 20160 0 g.g_y\[2\].g_x\[5\].t.r_d
rlabel metal2 45976 20776 45976 20776 0 g.g_y\[2\].g_x\[5\].t.r_h
rlabel metal2 52640 20776 52640 20776 0 g.g_y\[2\].g_x\[5\].t.r_v
rlabel metal2 48384 17752 48384 17752 0 g.g_y\[2\].g_x\[5\].t.w_si
rlabel metal2 46648 25816 46648 25816 0 g.g_y\[2\].g_x\[6\].t.out_sc
rlabel metal3 46648 25368 46648 25368 0 g.g_y\[2\].g_x\[6\].t.r_d
rlabel metal2 45752 22344 45752 22344 0 g.g_y\[2\].g_x\[6\].t.r_h
rlabel metal3 47208 28784 47208 28784 0 g.g_y\[2\].g_x\[6\].t.r_v
rlabel metal2 44856 27272 44856 27272 0 g.g_y\[2\].g_x\[6\].t.w_dh
rlabel metal2 42672 23800 42672 23800 0 g.g_y\[2\].g_x\[6\].t.w_na
rlabel metal2 48776 25872 48776 25872 0 g.g_y\[2\].g_x\[6\].t.w_si
rlabel metal2 36344 25592 36344 25592 0 g.g_y\[2\].g_x\[7\].t.out_sc
rlabel metal2 37688 25760 37688 25760 0 g.g_y\[2\].g_x\[7\].t.r_d
rlabel metal2 39032 22848 39032 22848 0 g.g_y\[2\].g_x\[7\].t.r_h
rlabel metal2 37688 24920 37688 24920 0 g.g_y\[2\].g_x\[7\].t.r_v
rlabel metal3 38920 21560 38920 21560 0 g.g_y\[2\].g_x\[7\].t.w_si
rlabel metal2 9912 12936 9912 12936 0 g.g_y\[3\].g_x\[0\].t.out_sc
rlabel metal2 4648 13160 4648 13160 0 g.g_y\[3\].g_x\[0\].t.r_d
rlabel metal2 5768 11312 5768 11312 0 g.g_y\[3\].g_x\[0\].t.r_h
rlabel metal2 15624 13384 15624 13384 0 g.g_y\[3\].g_x\[0\].t.r_v
rlabel metal2 11984 13048 11984 13048 0 g.g_y\[3\].g_x\[0\].t.w_si
rlabel metal2 15624 7168 15624 7168 0 g.g_y\[3\].g_x\[1\].t.out_sc
rlabel metal3 12600 6664 12600 6664 0 g.g_y\[3\].g_x\[1\].t.r_d
rlabel metal2 15288 7728 15288 7728 0 g.g_y\[3\].g_x\[1\].t.r_h
rlabel metal2 15512 10304 15512 10304 0 g.g_y\[3\].g_x\[1\].t.r_v
rlabel metal2 15176 11424 15176 11424 0 g.g_y\[3\].g_x\[1\].t.w_dh
rlabel metal2 8568 7896 8568 7896 0 g.g_y\[3\].g_x\[1\].t.w_na
rlabel metal2 13440 7560 13440 7560 0 g.g_y\[3\].g_x\[1\].t.w_si
rlabel metal2 23072 6552 23072 6552 0 g.g_y\[3\].g_x\[2\].t.out_sc
rlabel metal2 20440 6328 20440 6328 0 g.g_y\[3\].g_x\[2\].t.r_d
rlabel metal2 19880 8736 19880 8736 0 g.g_y\[3\].g_x\[2\].t.r_h
rlabel metal2 17976 12096 17976 12096 0 g.g_y\[3\].g_x\[2\].t.r_v
rlabel metal2 22120 9408 22120 9408 0 g.g_y\[3\].g_x\[2\].t.w_si
rlabel metal3 25368 12936 25368 12936 0 g.g_y\[3\].g_x\[3\].t.out_sc
rlabel metal2 20664 14056 20664 14056 0 g.g_y\[3\].g_x\[3\].t.r_d
rlabel metal3 22008 15288 22008 15288 0 g.g_y\[3\].g_x\[3\].t.r_h
rlabel metal3 18536 14168 18536 14168 0 g.g_y\[3\].g_x\[3\].t.r_v
rlabel metal2 24696 11144 24696 11144 0 g.g_y\[3\].g_x\[3\].t.w_dh
rlabel metal2 21336 13160 21336 13160 0 g.g_y\[3\].g_x\[3\].t.w_na
rlabel metal2 23072 11256 23072 11256 0 g.g_y\[3\].g_x\[3\].t.w_si
rlabel metal2 24920 18088 24920 18088 0 g.g_y\[3\].g_x\[4\].t.out_sc
rlabel metal2 23800 18704 23800 18704 0 g.g_y\[3\].g_x\[4\].t.r_d
rlabel metal3 31696 18424 31696 18424 0 g.g_y\[3\].g_x\[4\].t.r_h
rlabel metal2 35000 19656 35000 19656 0 g.g_y\[3\].g_x\[4\].t.r_v
rlabel metal3 23408 16744 23408 16744 0 g.g_y\[3\].g_x\[4\].t.w_si
rlabel metal3 36064 23688 36064 23688 0 g.g_y\[3\].g_x\[5\].t.out_sc
rlabel metal2 35448 23576 35448 23576 0 g.g_y\[3\].g_x\[5\].t.r_d
rlabel metal3 32200 21448 32200 21448 0 g.g_y\[3\].g_x\[5\].t.r_h
rlabel metal2 32200 26208 32200 26208 0 g.g_y\[3\].g_x\[5\].t.r_v
rlabel metal2 31752 22064 31752 22064 0 g.g_y\[3\].g_x\[5\].t.w_dh
rlabel metal3 32760 24808 32760 24808 0 g.g_y\[3\].g_x\[5\].t.w_na
rlabel metal2 33040 20888 33040 20888 0 g.g_y\[3\].g_x\[5\].t.w_si
rlabel metal2 24696 21336 24696 21336 0 g.g_y\[3\].g_x\[6\].t.out_sc
rlabel metal3 23464 21560 23464 21560 0 g.g_y\[3\].g_x\[6\].t.r_d
rlabel metal2 25256 24024 25256 24024 0 g.g_y\[3\].g_x\[6\].t.r_h
rlabel metal2 24528 26040 24528 26040 0 g.g_y\[3\].g_x\[6\].t.r_v
rlabel metal2 22568 20944 22568 20944 0 g.g_y\[3\].g_x\[6\].t.w_si
rlabel metal2 20552 22120 20552 22120 0 g.g_y\[3\].g_x\[7\].t.out_sc
rlabel metal2 19656 25256 19656 25256 0 g.g_y\[3\].g_x\[7\].t.r_d
rlabel metal2 23128 23632 23128 23632 0 g.g_y\[3\].g_x\[7\].t.r_h
rlabel metal2 15904 24696 15904 24696 0 g.g_y\[3\].g_x\[7\].t.r_v
rlabel metal2 17304 23464 17304 23464 0 g.g_y\[3\].g_x\[7\].t.w_dh
rlabel metal2 17976 27832 17976 27832 0 g.g_y\[3\].g_x\[7\].t.w_na
rlabel metal2 18424 22904 18424 22904 0 g.g_y\[3\].g_x\[7\].t.w_si
rlabel metal2 4984 25536 4984 25536 0 g.g_y\[4\].g_x\[0\].t.out_sc
rlabel metal2 5880 24864 5880 24864 0 g.g_y\[4\].g_x\[0\].t.r_d
rlabel metal3 3864 21672 3864 21672 0 g.g_y\[4\].g_x\[0\].t.r_h
rlabel metal2 2856 23632 2856 23632 0 g.g_y\[4\].g_x\[0\].t.r_v
rlabel metal2 3528 22568 3528 22568 0 g.g_y\[4\].g_x\[0\].t.w_dh
rlabel metal2 2968 26040 2968 26040 0 g.g_y\[4\].g_x\[0\].t.w_na
rlabel metal2 7560 25144 7560 25144 0 g.g_y\[4\].g_x\[0\].t.w_si
rlabel metal2 2968 19432 2968 19432 0 g.g_y\[4\].g_x\[1\].t.out_sc
rlabel metal3 5656 17416 5656 17416 0 g.g_y\[4\].g_x\[1\].t.r_d
rlabel metal3 10416 20104 10416 20104 0 g.g_y\[4\].g_x\[1\].t.r_h
rlabel metal2 10248 22904 10248 22904 0 g.g_y\[4\].g_x\[1\].t.r_v
rlabel metal3 2352 20328 2352 20328 0 g.g_y\[4\].g_x\[1\].t.w_si
rlabel metal2 11536 19096 11536 19096 0 g.g_y\[4\].g_x\[2\].t.out_sc
rlabel metal2 14168 17192 14168 17192 0 g.g_y\[4\].g_x\[2\].t.r_d
rlabel metal2 12040 21168 12040 21168 0 g.g_y\[4\].g_x\[2\].t.r_h
rlabel metal3 17024 13720 17024 13720 0 g.g_y\[4\].g_x\[2\].t.r_v
rlabel metal2 14840 15624 14840 15624 0 g.g_y\[4\].g_x\[2\].t.w_dh
rlabel metal2 11368 18480 11368 18480 0 g.g_y\[4\].g_x\[2\].t.w_na
rlabel metal2 12376 13776 12376 13776 0 g.g_y\[4\].g_x\[2\].t.w_si
rlabel metal3 17864 22120 17864 22120 0 g.g_y\[4\].g_x\[3\].t.out_sc
rlabel metal2 15512 18424 15512 18424 0 g.g_y\[4\].g_x\[3\].t.r_d
rlabel metal2 15568 22344 15568 22344 0 g.g_y\[4\].g_x\[3\].t.r_h
rlabel metal3 17416 17640 17416 17640 0 g.g_y\[4\].g_x\[3\].t.r_v
rlabel metal3 21392 20104 21392 20104 0 g.g_y\[4\].g_x\[3\].t.w_si
rlabel metal2 12040 25592 12040 25592 0 g.g_y\[4\].g_x\[4\].t.out_sc
rlabel metal3 11984 27944 11984 27944 0 g.g_y\[4\].g_x\[4\].t.r_d
rlabel metal2 17640 25760 17640 25760 0 g.g_y\[4\].g_x\[4\].t.r_h
rlabel metal3 22008 36456 22008 36456 0 g.g_y\[4\].g_x\[4\].t.r_v
rlabel metal2 14728 25144 14728 25144 0 g.g_y\[4\].g_x\[4\].t.w_dh
rlabel metal2 22792 26040 22792 26040 0 g.g_y\[4\].g_x\[4\].t.w_na
rlabel metal2 11816 24360 11816 24360 0 g.g_y\[4\].g_x\[4\].t.w_si
rlabel metal2 26264 28224 26264 28224 0 g.g_y\[4\].g_x\[5\].t.out_sc
rlabel metal2 28504 30296 28504 30296 0 g.g_y\[4\].g_x\[5\].t.r_d
rlabel metal2 24248 30240 24248 30240 0 g.g_y\[4\].g_x\[5\].t.r_h
rlabel metal2 31416 28336 31416 28336 0 g.g_y\[4\].g_x\[5\].t.r_v
rlabel metal2 22680 28280 22680 28280 0 g.g_y\[4\].g_x\[5\].t.w_si
rlabel metal2 28056 32424 28056 32424 0 g.g_y\[4\].g_x\[6\].t.out_sc
rlabel metal3 24080 32648 24080 32648 0 g.g_y\[4\].g_x\[6\].t.r_d
rlabel metal2 20272 31192 20272 31192 0 g.g_y\[4\].g_x\[6\].t.r_h
rlabel metal2 26712 33656 26712 33656 0 g.g_y\[4\].g_x\[6\].t.r_v
rlabel metal2 23240 33600 23240 33600 0 g.g_y\[4\].g_x\[6\].t.w_dh
rlabel metal2 18312 34384 18312 34384 0 g.g_y\[4\].g_x\[6\].t.w_na
rlabel metal3 25256 31640 25256 31640 0 g.g_y\[4\].g_x\[6\].t.w_si
rlabel metal2 11312 32760 11312 32760 0 g.g_y\[4\].g_x\[7\].t.out_sc
rlabel metal2 12152 31360 12152 31360 0 g.g_y\[4\].g_x\[7\].t.r_d
rlabel metal2 13384 33376 13384 33376 0 g.g_y\[4\].g_x\[7\].t.r_h
rlabel metal2 12376 29848 12376 29848 0 g.g_y\[4\].g_x\[7\].t.r_v
rlabel metal2 16408 29848 16408 29848 0 g.g_y\[4\].g_x\[7\].t.w_si
rlabel metal2 1736 28784 1736 28784 0 g.g_y\[5\].g_x\[0\].t.out_sc
rlabel metal2 3080 28504 3080 28504 0 g.g_y\[5\].g_x\[0\].t.r_d
rlabel metal2 3192 28672 3192 28672 0 g.g_y\[5\].g_x\[0\].t.r_h
rlabel metal2 2408 30184 2408 30184 0 g.g_y\[5\].g_x\[0\].t.r_v
rlabel metal2 3920 29512 3920 29512 0 g.g_y\[5\].g_x\[0\].t.w_si
rlabel metal2 9128 29064 9128 29064 0 g.g_y\[5\].g_x\[1\].t.out_sc
rlabel metal3 6888 36680 6888 36680 0 g.g_y\[5\].g_x\[1\].t.r_d
rlabel metal2 9688 33824 9688 33824 0 g.g_y\[5\].g_x\[1\].t.r_h
rlabel metal2 8568 39144 8568 39144 0 g.g_y\[5\].g_x\[1\].t.r_v
rlabel metal2 9744 32760 9744 32760 0 g.g_y\[5\].g_x\[1\].t.w_dh
rlabel metal3 7392 37464 7392 37464 0 g.g_y\[5\].g_x\[1\].t.w_na
rlabel metal2 7056 28728 7056 28728 0 g.g_y\[5\].g_x\[1\].t.w_si
rlabel metal2 15176 41048 15176 41048 0 g.g_y\[5\].g_x\[2\].t.out_sc
rlabel metal3 10640 37016 10640 37016 0 g.g_y\[5\].g_x\[2\].t.r_d
rlabel metal2 12040 41664 12040 41664 0 g.g_y\[5\].g_x\[2\].t.r_h
rlabel metal2 12824 42672 12824 42672 0 g.g_y\[5\].g_x\[2\].t.r_v
rlabel metal2 18480 35896 18480 35896 0 g.g_y\[5\].g_x\[2\].t.w_si
rlabel metal2 16632 43960 16632 43960 0 g.g_y\[5\].g_x\[3\].t.out_sc
rlabel metal2 20328 42224 20328 42224 0 g.g_y\[5\].g_x\[3\].t.r_d
rlabel metal3 19656 39480 19656 39480 0 g.g_y\[5\].g_x\[3\].t.r_h
rlabel metal3 17528 46088 17528 46088 0 g.g_y\[5\].g_x\[3\].t.r_v
rlabel metal2 16632 42392 16632 42392 0 g.g_y\[5\].g_x\[3\].t.w_dh
rlabel metal2 17584 40488 17584 40488 0 g.g_y\[5\].g_x\[3\].t.w_na
rlabel metal2 14728 43120 14728 43120 0 g.g_y\[5\].g_x\[3\].t.w_si
rlabel metal3 20496 38024 20496 38024 0 g.g_y\[5\].g_x\[4\].t.out_sc
rlabel metal2 20832 41272 20832 41272 0 g.g_y\[5\].g_x\[4\].t.r_d
rlabel metal3 24192 42728 24192 42728 0 g.g_y\[5\].g_x\[4\].t.r_h
rlabel metal2 22568 39032 22568 39032 0 g.g_y\[5\].g_x\[4\].t.r_v
rlabel metal2 18648 38024 18648 38024 0 g.g_y\[5\].g_x\[4\].t.w_si
rlabel metal2 24248 48188 24248 48188 0 g.g_y\[5\].g_x\[5\].t.out_sc
rlabel metal2 24808 48048 24808 48048 0 g.g_y\[5\].g_x\[5\].t.r_d
rlabel metal2 24024 48328 24024 48328 0 g.g_y\[5\].g_x\[5\].t.r_h
rlabel metal3 24808 47992 24808 47992 0 g.g_y\[5\].g_x\[5\].t.r_v
rlabel metal3 25088 46760 25088 46760 0 g.g_y\[5\].g_x\[5\].t.w_dh
rlabel metal2 28168 44800 28168 44800 0 g.g_y\[5\].g_x\[5\].t.w_na
rlabel metal2 22120 45472 22120 45472 0 g.g_y\[5\].g_x\[5\].t.w_si
rlabel metal2 18200 54376 18200 54376 0 g.g_y\[5\].g_x\[6\].t.out_sc
rlabel metal2 20104 53144 20104 53144 0 g.g_y\[5\].g_x\[6\].t.r_d
rlabel metal2 21112 57120 21112 57120 0 g.g_y\[5\].g_x\[6\].t.r_h
rlabel metal2 25704 55776 25704 55776 0 g.g_y\[5\].g_x\[6\].t.r_v
rlabel metal2 19768 52528 19768 52528 0 g.g_y\[5\].g_x\[6\].t.w_si
rlabel metal2 12936 56336 12936 56336 0 g.g_y\[5\].g_x\[7\].t.out_sc
rlabel metal2 16184 58576 16184 58576 0 g.g_y\[5\].g_x\[7\].t.r_d
rlabel metal2 19544 54544 19544 54544 0 g.g_y\[5\].g_x\[7\].t.r_h
rlabel metal2 19488 58968 19488 58968 0 g.g_y\[5\].g_x\[7\].t.r_v
rlabel metal2 16408 54544 16408 54544 0 g.g_y\[5\].g_x\[7\].t.w_dh
rlabel metal2 14616 58296 14616 58296 0 g.g_y\[5\].g_x\[7\].t.w_na
rlabel metal3 15148 52696 15148 52696 0 g.g_y\[5\].g_x\[7\].t.w_si
rlabel metal2 4984 48664 4984 48664 0 g.g_y\[6\].g_x\[0\].t.out_sc
rlabel metal2 1792 45640 1792 45640 0 g.g_y\[6\].g_x\[0\].t.r_d
rlabel metal3 5320 49000 5320 49000 0 g.g_y\[6\].g_x\[0\].t.r_h
rlabel metal3 5712 38808 5712 38808 0 g.g_y\[6\].g_x\[0\].t.r_v
rlabel metal3 2352 42952 2352 42952 0 g.g_y\[6\].g_x\[0\].t.w_dh
rlabel metal2 2184 38780 2184 38780 0 g.g_y\[6\].g_x\[0\].t.w_na
rlabel metal2 2520 47096 2520 47096 0 g.g_y\[6\].g_x\[0\].t.w_si
rlabel metal3 5768 47320 5768 47320 0 g.g_y\[6\].g_x\[1\].t.out_sc
rlabel metal3 5712 41944 5712 41944 0 g.g_y\[6\].g_x\[1\].t.r_d
rlabel metal2 8624 47656 8624 47656 0 g.g_y\[6\].g_x\[1\].t.r_h
rlabel metal2 6552 40376 6552 40376 0 g.g_y\[6\].g_x\[1\].t.r_v
rlabel metal2 3976 41496 3976 41496 0 g.g_y\[6\].g_x\[1\].t.w_si
rlabel metal2 10136 49756 10136 49756 0 g.g_y\[6\].g_x\[2\].t.out_sc
rlabel metal2 13608 47152 13608 47152 0 g.g_y\[6\].g_x\[2\].t.r_d
rlabel metal2 10696 48832 10696 48832 0 g.g_y\[6\].g_x\[2\].t.r_h
rlabel metal2 9744 46648 9744 46648 0 g.g_y\[6\].g_x\[2\].t.r_v
rlabel metal2 10752 48328 10752 48328 0 g.g_y\[6\].g_x\[2\].t.w_dh
rlabel metal2 11368 49756 11368 49756 0 g.g_y\[6\].g_x\[2\].t.w_na
rlabel metal2 8456 46816 8456 46816 0 g.g_y\[6\].g_x\[2\].t.w_si
rlabel metal2 17304 51800 17304 51800 0 g.g_y\[6\].g_x\[3\].t.out_sc
rlabel metal3 17640 49784 17640 49784 0 g.g_y\[6\].g_x\[3\].t.r_d
rlabel metal2 20328 49952 20328 49952 0 g.g_y\[6\].g_x\[3\].t.r_h
rlabel metal3 16632 46760 16632 46760 0 g.g_y\[6\].g_x\[3\].t.r_v
rlabel metal2 15848 50960 15848 50960 0 g.g_y\[6\].g_x\[3\].t.w_si
rlabel metal2 38024 53648 38024 53648 0 g.g_y\[6\].g_x\[4\].t.out_sc
rlabel metal2 39032 53256 39032 53256 0 g.g_y\[6\].g_x\[4\].t.r_d
rlabel metal2 34552 53200 34552 53200 0 g.g_y\[6\].g_x\[4\].t.r_h
rlabel metal2 39704 49112 39704 49112 0 g.g_y\[6\].g_x\[4\].t.r_v
rlabel metal2 37352 50792 37352 50792 0 g.g_y\[6\].g_x\[4\].t.w_dh
rlabel metal2 36624 49896 36624 49896 0 g.g_y\[6\].g_x\[4\].t.w_na
rlabel metal2 34776 51352 34776 51352 0 g.g_y\[6\].g_x\[4\].t.w_si
rlabel metal2 28168 53368 28168 53368 0 g.g_y\[6\].g_x\[5\].t.out_sc
rlabel metal2 28952 51800 28952 51800 0 g.g_y\[6\].g_x\[5\].t.r_d
rlabel metal2 29288 54096 29288 54096 0 g.g_y\[6\].g_x\[5\].t.r_h
rlabel metal2 29848 48328 29848 48328 0 g.g_y\[6\].g_x\[5\].t.r_v
rlabel metal2 26600 51352 26600 51352 0 g.g_y\[6\].g_x\[5\].t.w_si
rlabel metal2 35672 57624 35672 57624 0 g.g_y\[6\].g_x\[6\].t.out_sc
rlabel metal2 33768 58968 33768 58968 0 g.g_y\[6\].g_x\[6\].t.r_d
rlabel metal3 32144 59864 32144 59864 0 g.g_y\[6\].g_x\[6\].t.r_h
rlabel via2 36680 55272 36680 55272 0 g.g_y\[6\].g_x\[6\].t.r_v
rlabel metal2 33432 55552 33432 55552 0 g.g_y\[6\].g_x\[6\].t.w_dh
rlabel metal2 30856 58128 30856 58128 0 g.g_y\[6\].g_x\[6\].t.w_na
rlabel metal2 31864 54096 31864 54096 0 g.g_y\[6\].g_x\[6\].t.w_si
rlabel metal2 22120 59696 22120 59696 0 g.g_y\[6\].g_x\[7\].t.out_sc
rlabel metal2 22568 59136 22568 59136 0 g.g_y\[6\].g_x\[7\].t.r_d
rlabel metal3 25088 59192 25088 59192 0 g.g_y\[6\].g_x\[7\].t.r_h
rlabel metal2 20552 56504 20552 56504 0 g.g_y\[6\].g_x\[7\].t.r_v
rlabel metal2 25928 53480 25928 53480 0 g.g_y\[6\].g_x\[7\].t.w_si
rlabel metal2 29400 36008 29400 36008 0 g.g_y\[7\].g_x\[0\].t.out_sc
rlabel metal2 26152 39144 26152 39144 0 g.g_y\[7\].g_x\[0\].t.r_d
rlabel metal3 28336 41160 28336 41160 0 g.g_y\[7\].g_x\[0\].t.r_h
rlabel metal2 30632 36456 30632 36456 0 g.g_y\[7\].g_x\[0\].t.r_v
rlabel metal2 25984 39480 25984 39480 0 g.g_y\[7\].g_x\[0\].t.w_si
rlabel metal2 32200 45360 32200 45360 0 g.g_y\[7\].g_x\[1\].t.out_sc
rlabel metal3 34048 41832 34048 41832 0 g.g_y\[7\].g_x\[1\].t.r_d
rlabel metal2 33432 44408 33432 44408 0 g.g_y\[7\].g_x\[1\].t.r_h
rlabel metal2 34328 43120 34328 43120 0 g.g_y\[7\].g_x\[1\].t.r_v
rlabel metal2 31528 43960 31528 43960 0 g.g_y\[7\].g_x\[1\].t.w_dh
rlabel metal2 33432 41664 33432 41664 0 g.g_y\[7\].g_x\[1\].t.w_na
rlabel metal2 30072 44352 30072 44352 0 g.g_y\[7\].g_x\[1\].t.w_si
rlabel metal3 37688 49000 37688 49000 0 g.g_y\[7\].g_x\[2\].t.out_sc
rlabel metal2 37688 47656 37688 47656 0 g.g_y\[7\].g_x\[2\].t.r_d
rlabel metal2 40488 47208 40488 47208 0 g.g_y\[7\].g_x\[2\].t.r_h
rlabel metal2 40152 40936 40152 40936 0 g.g_y\[7\].g_x\[2\].t.r_v
rlabel metal2 40880 45304 40880 45304 0 g.g_y\[7\].g_x\[2\].t.w_si
rlabel metal2 44296 45808 44296 45808 0 g.g_y\[7\].g_x\[3\].t.out_sc
rlabel metal2 45416 41496 45416 41496 0 g.g_y\[7\].g_x\[3\].t.r_d
rlabel metal2 46816 45304 46816 45304 0 g.g_y\[7\].g_x\[3\].t.r_h
rlabel metal2 49112 39480 49112 39480 0 g.g_y\[7\].g_x\[3\].t.r_v
rlabel metal2 44520 42056 44520 42056 0 g.g_y\[7\].g_x\[3\].t.w_dh
rlabel metal2 42616 40656 42616 40656 0 g.g_y\[7\].g_x\[3\].t.w_na
rlabel metal2 42728 44408 42728 44408 0 g.g_y\[7\].g_x\[3\].t.w_si
rlabel metal3 45752 52248 45752 52248 0 g.g_y\[7\].g_x\[4\].t.out_sc
rlabel metal2 43848 52024 43848 52024 0 g.g_y\[7\].g_x\[4\].t.r_d
rlabel metal3 47936 50344 47936 50344 0 g.g_y\[7\].g_x\[4\].t.r_h
rlabel metal3 43456 51576 43456 51576 0 g.g_y\[7\].g_x\[4\].t.r_v
rlabel metal2 43064 51240 43064 51240 0 g.g_y\[7\].g_x\[4\].t.w_si
rlabel metal2 58744 50792 58744 50792 0 g.g_y\[7\].g_x\[5\].t.out_sc
rlabel metal3 56896 50568 56896 50568 0 g.g_y\[7\].g_x\[5\].t.r_d
rlabel metal3 58016 49784 58016 49784 0 g.g_y\[7\].g_x\[5\].t.r_h
rlabel metal2 55496 48608 55496 48608 0 g.g_y\[7\].g_x\[5\].t.r_v
rlabel metal2 51744 46760 51744 46760 0 g.g_y\[7\].g_x\[5\].t.w_dh
rlabel metal2 52472 47936 52472 47936 0 g.g_y\[7\].g_x\[5\].t.w_na
rlabel metal3 49896 50680 49896 50680 0 g.g_y\[7\].g_x\[5\].t.w_si
rlabel metal2 59976 53200 59976 53200 0 g.g_y\[7\].g_x\[6\].t.out_sc
rlabel metal2 55832 57344 55832 57344 0 g.g_y\[7\].g_x\[6\].t.r_d
rlabel metal2 53256 54488 53256 54488 0 g.g_y\[7\].g_x\[6\].t.r_h
rlabel metal2 59640 53200 59640 53200 0 g.g_y\[7\].g_x\[6\].t.r_v
rlabel metal2 59192 50848 59192 50848 0 g.g_y\[7\].g_x\[6\].t.w_si
rlabel metal2 46760 56840 46760 56840 0 g.g_y\[7\].g_x\[7\].t.r_d
rlabel metal2 51464 57344 51464 57344 0 g.g_y\[7\].g_x\[7\].t.r_h
rlabel metal3 51016 54264 51016 54264 0 g.g_y\[7\].g_x\[7\].t.r_v
rlabel metal2 46536 53648 46536 53648 0 g.g_y\[7\].g_x\[7\].t.w_dh
rlabel metal2 42952 55776 42952 55776 0 g.g_y\[7\].g_x\[7\].t.w_na
rlabel metal2 44968 54152 44968 54152 0 g.g_y\[7\].g_x\[7\].t.w_si
rlabel metal2 1736 54824 1736 54824 0 in[0]
rlabel metal2 62272 18984 62272 18984 0 in[10]
rlabel metal3 63154 30296 63154 30296 0 in[11]
rlabel metal2 32368 3416 32368 3416 0 in[12]
rlabel metal3 30016 3752 30016 3752 0 in[13]
rlabel metal2 62160 14392 62160 14392 0 in[14]
rlabel metal3 63154 27608 63154 27608 0 in[15]
rlabel metal2 60200 19096 60200 19096 0 in[16]
rlabel metal2 47992 4144 47992 4144 0 in[1]
rlabel metal4 61656 31528 61656 31528 0 in[2]
rlabel metal2 31640 1246 31640 1246 0 in[3]
rlabel metal2 29624 2058 29624 2058 0 in[4]
rlabel metal2 1736 11816 1736 11816 0 in[5]
rlabel metal2 1736 24080 1736 24080 0 in[6]
rlabel metal2 1736 26600 1736 26600 0 in[7]
rlabel metal3 2072 44296 2072 44296 0 in[8]
rlabel metal3 31808 59976 31808 59976 0 in[9]
rlabel metal2 2072 53032 2072 53032 0 net1
rlabel metal2 41160 33992 41160 33992 0 net10
rlabel metal2 45752 40320 45752 40320 0 net100
rlabel metal2 43400 46648 43400 46648 0 net101
rlabel metal2 46032 52136 46032 52136 0 net102
rlabel metal2 45864 51856 45864 51856 0 net103
rlabel metal3 53760 49224 53760 49224 0 net104
rlabel metal3 57736 50456 57736 50456 0 net105
rlabel metal2 53816 56504 53816 56504 0 net106
rlabel metal2 45192 57120 45192 57120 0 net107
rlabel metal2 45528 56560 45528 56560 0 net108
rlabel metal2 47712 56728 47712 56728 0 net109
rlabel metal2 31528 15736 31528 15736 0 net11
rlabel metal2 2184 24136 2184 24136 0 net110
rlabel metal2 2072 16240 2072 16240 0 net111
rlabel metal2 17640 22288 17640 22288 0 net112
rlabel metal2 16632 23856 16632 23856 0 net113
rlabel metal2 22344 11648 22344 11648 0 net114
rlabel metal2 2856 24248 2856 24248 0 net115
rlabel metal2 14112 51352 14112 51352 0 net116
rlabel metal2 2800 48888 2800 48888 0 net117
rlabel metal2 21448 45640 21448 45640 0 net118
rlabel metal2 25256 34608 25256 34608 0 net119
rlabel metal2 29512 6440 29512 6440 0 net12
rlabel metal3 17640 54936 17640 54936 0 net120
rlabel metal2 2464 21560 2464 21560 0 net121
rlabel metal2 58072 13608 58072 13608 0 net122
rlabel metal2 35000 21112 35000 21112 0 net123
rlabel metal2 52976 10024 52976 10024 0 net124
rlabel metal2 51128 6216 51128 6216 0 net125
rlabel metal2 59416 14448 59416 14448 0 net126
rlabel metal2 41384 54152 41384 54152 0 net127
rlabel metal2 40656 47432 40656 47432 0 net128
rlabel metal2 47096 32368 47096 32368 0 net129
rlabel metal2 2072 11424 2072 11424 0 net13
rlabel metal2 50064 39256 50064 39256 0 net130
rlabel metal2 61544 50792 61544 50792 0 net131
rlabel metal2 47656 57680 47656 57680 0 net132
rlabel metal2 46200 18144 46200 18144 0 net133
rlabel metal2 3080 51240 3080 51240 0 net134
rlabel metal2 7448 2030 7448 2030 0 net135
rlabel metal2 62216 58912 62216 58912 0 net136
rlabel metal2 38360 62734 38360 62734 0 net137
rlabel metal2 7672 23800 7672 23800 0 net14
rlabel metal2 2072 28056 2072 28056 0 net15
rlabel metal3 2744 44184 2744 44184 0 net16
rlabel metal2 29176 50400 29176 50400 0 net17
rlabel metal2 52192 39816 52192 39816 0 net18
rlabel metal2 51800 31024 51800 31024 0 net19
rlabel metal2 47992 25900 47992 25900 0 net2
rlabel metal2 40264 4368 40264 4368 0 net20
rlabel metal3 19992 21616 19992 21616 0 net21
rlabel metal2 4088 33376 4088 33376 0 net22
rlabel metal2 17080 58352 17080 58352 0 net23
rlabel metal2 21504 56728 21504 56728 0 net24
rlabel metal2 48216 58520 48216 58520 0 net25
rlabel metal2 44240 54376 44240 54376 0 net26
rlabel metal2 34328 33096 34328 33096 0 net27
rlabel metal2 38808 31136 38808 31136 0 net28
rlabel metal2 45192 32536 45192 32536 0 net29
rlabel metal2 34944 25592 34944 25592 0 net3
rlabel metal2 45472 34216 45472 34216 0 net30
rlabel metal2 53368 39032 53368 39032 0 net31
rlabel metal3 60088 34216 60088 34216 0 net32
rlabel metal2 58744 43848 58744 43848 0 net33
rlabel metal2 58744 45976 58744 45976 0 net34
rlabel metal3 32368 15960 32368 15960 0 net35
rlabel metal2 39144 12376 39144 12376 0 net36
rlabel metal2 38808 16240 38808 16240 0 net37
rlabel metal2 54264 12152 54264 12152 0 net38
rlabel metal3 54992 15400 54992 15400 0 net39
rlabel metal2 31416 23632 31416 23632 0 net4
rlabel metal2 61488 22232 61488 22232 0 net40
rlabel metal4 60984 20944 60984 20944 0 net41
rlabel metal3 46704 29400 46704 29400 0 net42
rlabel metal2 59808 14280 59808 14280 0 net43
rlabel metal2 26824 7448 26824 7448 0 net44
rlabel metal2 26040 5824 26040 5824 0 net45
rlabel metal2 43400 5040 43400 5040 0 net46
rlabel metal2 45752 4480 45752 4480 0 net47
rlabel metal2 43624 10752 43624 10752 0 net48
rlabel metal2 41216 18200 41216 18200 0 net49
rlabel metal2 33096 26600 33096 26600 0 net5
rlabel metal2 41720 20384 41720 20384 0 net50
rlabel metal2 42504 22232 42504 22232 0 net51
rlabel metal2 47264 26600 47264 26600 0 net52
rlabel metal3 12264 6776 12264 6776 0 net53
rlabel metal2 25256 6216 25256 6216 0 net54
rlabel metal2 21336 7056 21336 7056 0 net55
rlabel metal2 20216 15260 20216 15260 0 net56
rlabel metal2 25368 15848 25368 15848 0 net57
rlabel metal3 24136 18536 24136 18536 0 net58
rlabel via3 24808 17080 24808 17080 0 net59
rlabel metal2 48160 31528 48160 31528 0 net6
rlabel metal3 32928 25256 32928 25256 0 net60
rlabel metal2 23464 21896 23464 21896 0 net61
rlabel metal3 20552 25368 20552 25368 0 net62
rlabel metal2 21896 23744 21896 23744 0 net63
rlabel metal2 2408 24584 2408 24584 0 net64
rlabel metal2 2520 23352 2520 23352 0 net65
rlabel metal2 11144 19824 11144 19824 0 net66
rlabel metal2 17248 20216 17248 20216 0 net67
rlabel metal2 17304 22344 17304 22344 0 net68
rlabel metal2 11368 28280 11368 28280 0 net69
rlabel metal2 61320 17920 61320 17920 0 net7
rlabel metal2 23576 32312 23576 32312 0 net70
rlabel metal2 22232 32480 22232 32480 0 net71
rlabel metal2 19880 33936 19880 33936 0 net72
rlabel metal2 27384 34552 27384 34552 0 net73
rlabel metal2 9464 28560 9464 28560 0 net74
rlabel metal2 15400 35000 15400 35000 0 net75
rlabel metal3 11032 34328 11032 34328 0 net76
rlabel metal3 18368 41720 18368 41720 0 net77
rlabel metal3 17640 43624 17640 43624 0 net78
rlabel metal2 19544 38136 19544 38136 0 net79
rlabel metal2 38920 17304 38920 17304 0 net8
rlabel metal2 25032 47488 25032 47488 0 net80
rlabel metal2 27272 48664 27272 48664 0 net81
rlabel metal2 18536 54656 18536 54656 0 net82
rlabel metal2 15736 57120 15736 57120 0 net83
rlabel metal2 14168 59528 14168 59528 0 net84
rlabel metal2 2408 39872 2408 39872 0 net85
rlabel metal2 3080 47040 3080 47040 0 net86
rlabel metal2 11704 51968 11704 51968 0 net87
rlabel metal2 12992 52024 12992 52024 0 net88
rlabel metal2 18424 49504 18424 49504 0 net89
rlabel metal2 34216 25984 34216 25984 0 net9
rlabel metal3 39032 53032 39032 53032 0 net90
rlabel metal2 25368 53704 25368 53704 0 net91
rlabel metal2 29848 59416 29848 59416 0 net92
rlabel metal2 35168 57736 35168 57736 0 net93
rlabel metal2 27720 41776 27720 41776 0 net94
rlabel metal2 27216 39032 27216 39032 0 net95
rlabel metal2 33488 42504 33488 42504 0 net96
rlabel metal3 33376 45640 33376 45640 0 net97
rlabel metal2 39032 43568 39032 43568 0 net98
rlabel metal3 40880 47320 40880 47320 0 net99
rlabel metal3 61992 43176 61992 43176 0 out[0]
rlabel metal3 62734 30968 62734 30968 0 out[1]
rlabel metal2 38360 1246 38360 1246 0 out[2]
rlabel metal3 1358 24248 1358 24248 0 out[3]
rlabel metal3 1848 33544 1848 33544 0 out[4]
rlabel metal3 17080 60200 17080 60200 0 out[5]
rlabel metal2 26264 61362 26264 61362 0 out[6]
rlabel metal3 49112 59416 49112 59416 0 out[7]
rlabel metal3 48384 60200 48384 60200 0 out[8]
<< properties >>
string FIXED_BBOX 0 0 64000 64000
<< end >>
