magic
tech gf180mcuD
magscale 1 5
timestamp 1702353082
<< obsm1 >>
rect 672 1538 19400 18454
<< metal2 >>
rect 7392 19600 7448 20000
rect 7728 19600 7784 20000
rect 8064 19600 8120 20000
rect 8400 19600 8456 20000
rect 8736 19600 8792 20000
rect 9072 19600 9128 20000
rect 9408 19600 9464 20000
rect 9744 19600 9800 20000
rect 10080 19600 10136 20000
rect 10416 19600 10472 20000
rect 10752 19600 10808 20000
rect 11088 19600 11144 20000
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12096 0 12152 400
<< obsm2 >>
rect 854 19570 7362 19600
rect 7478 19570 7698 19600
rect 7814 19570 8034 19600
rect 8150 19570 8370 19600
rect 8486 19570 8706 19600
rect 8822 19570 9042 19600
rect 9158 19570 9378 19600
rect 9494 19570 9714 19600
rect 9830 19570 10050 19600
rect 10166 19570 10386 19600
rect 10502 19570 10722 19600
rect 10838 19570 11058 19600
rect 11174 19570 19386 19600
rect 854 430 19386 19570
rect 854 400 6354 430
rect 6470 400 6690 430
rect 6806 400 7026 430
rect 7142 400 7362 430
rect 7478 400 7698 430
rect 7814 400 8034 430
rect 8150 400 8370 430
rect 8486 400 8706 430
rect 8822 400 9042 430
rect 9158 400 9378 430
rect 9494 400 9714 430
rect 9830 400 10050 430
rect 10166 400 10386 430
rect 10502 400 10722 430
rect 10838 400 11058 430
rect 11174 400 11394 430
rect 11510 400 11730 430
rect 11846 400 12066 430
rect 12182 400 19386 430
<< metal3 >>
rect 0 12768 400 12824
rect 0 12432 400 12488
rect 0 12096 400 12152
rect 19600 12096 20000 12152
rect 0 11760 400 11816
rect 19600 11760 20000 11816
rect 0 11424 400 11480
rect 19600 11424 20000 11480
rect 0 11088 400 11144
rect 19600 11088 20000 11144
rect 0 10752 400 10808
rect 19600 10752 20000 10808
rect 0 10416 400 10472
rect 19600 10416 20000 10472
rect 0 10080 400 10136
rect 19600 10080 20000 10136
rect 0 9744 400 9800
rect 19600 9744 20000 9800
rect 0 9408 400 9464
rect 19600 9408 20000 9464
rect 0 9072 400 9128
rect 19600 9072 20000 9128
rect 0 8736 400 8792
rect 19600 8736 20000 8792
rect 0 8400 400 8456
rect 19600 8400 20000 8456
rect 0 8064 400 8120
rect 19600 8064 20000 8120
rect 0 7728 400 7784
rect 19600 7728 20000 7784
rect 19600 7392 20000 7448
rect 19600 7056 20000 7112
<< obsm3 >>
rect 400 12854 19600 18438
rect 430 12738 19600 12854
rect 400 12518 19600 12738
rect 430 12402 19600 12518
rect 400 12182 19600 12402
rect 430 12066 19570 12182
rect 400 11846 19600 12066
rect 430 11730 19570 11846
rect 400 11510 19600 11730
rect 430 11394 19570 11510
rect 400 11174 19600 11394
rect 430 11058 19570 11174
rect 400 10838 19600 11058
rect 430 10722 19570 10838
rect 400 10502 19600 10722
rect 430 10386 19570 10502
rect 400 10166 19600 10386
rect 430 10050 19570 10166
rect 400 9830 19600 10050
rect 430 9714 19570 9830
rect 400 9494 19600 9714
rect 430 9378 19570 9494
rect 400 9158 19600 9378
rect 430 9042 19570 9158
rect 400 8822 19600 9042
rect 430 8706 19570 8822
rect 400 8486 19600 8706
rect 430 8370 19570 8486
rect 400 8150 19600 8370
rect 430 8034 19570 8150
rect 400 7814 19600 8034
rect 430 7698 19570 7814
rect 400 7478 19600 7698
rect 400 7362 19570 7478
rect 400 7142 19600 7362
rect 400 7026 19570 7142
rect 400 1554 19600 7026
<< metal4 >>
rect 2923 1538 3083 18454
rect 5254 1538 5414 18454
rect 7585 1538 7745 18454
rect 9916 1538 10076 18454
rect 12247 1538 12407 18454
rect 14578 1538 14738 18454
rect 16909 1538 17069 18454
rect 19240 1538 19400 18454
<< labels >>
rlabel metal3 s 19600 7056 20000 7112 6 out[0]
port 1 nsew signal output
rlabel metal3 s 0 9744 400 9800 6 out[10]
port 2 nsew signal output
rlabel metal2 s 7392 19600 7448 20000 6 out[11]
port 3 nsew signal output
rlabel metal3 s 19600 7728 20000 7784 6 out[1]
port 4 nsew signal output
rlabel metal3 s 19600 12096 20000 12152 6 out[2]
port 5 nsew signal output
rlabel metal3 s 19600 10752 20000 10808 6 out[3]
port 6 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 out[4]
port 7 nsew signal output
rlabel metal2 s 12096 0 12152 400 6 out[5]
port 8 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 out[6]
port 9 nsew signal output
rlabel metal2 s 6384 0 6440 400 6 out[7]
port 10 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 out[8]
port 11 nsew signal output
rlabel metal2 s 8400 19600 8456 20000 6 out[9]
port 12 nsew signal output
rlabel metal3 s 19600 9408 20000 9464 6 proj_out[0]
port 13 nsew signal input
rlabel metal3 s 0 9072 400 9128 6 proj_out[10]
port 14 nsew signal input
rlabel metal2 s 9408 19600 9464 20000 6 proj_out[11]
port 15 nsew signal input
rlabel metal3 s 19600 10080 20000 10136 6 proj_out[12]
port 16 nsew signal input
rlabel metal3 s 19600 8736 20000 8792 6 proj_out[13]
port 17 nsew signal input
rlabel metal3 s 19600 11088 20000 11144 6 proj_out[14]
port 18 nsew signal input
rlabel metal3 s 19600 11760 20000 11816 6 proj_out[15]
port 19 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 proj_out[16]
port 20 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 proj_out[17]
port 21 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 proj_out[18]
port 22 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 proj_out[19]
port 23 nsew signal input
rlabel metal3 s 19600 8400 20000 8456 6 proj_out[1]
port 24 nsew signal input
rlabel metal3 s 0 10752 400 10808 6 proj_out[20]
port 25 nsew signal input
rlabel metal2 s 9072 19600 9128 20000 6 proj_out[21]
port 26 nsew signal input
rlabel metal3 s 0 10080 400 10136 6 proj_out[22]
port 27 nsew signal input
rlabel metal2 s 8736 19600 8792 20000 6 proj_out[23]
port 28 nsew signal input
rlabel metal3 s 19600 9744 20000 9800 6 proj_out[24]
port 29 nsew signal input
rlabel metal3 s 19600 9072 20000 9128 6 proj_out[25]
port 30 nsew signal input
rlabel metal2 s 10416 19600 10472 20000 6 proj_out[26]
port 31 nsew signal input
rlabel metal2 s 10080 19600 10136 20000 6 proj_out[27]
port 32 nsew signal input
rlabel metal3 s 0 7728 400 7784 6 proj_out[28]
port 33 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 proj_out[29]
port 34 nsew signal input
rlabel metal3 s 19600 11424 20000 11480 6 proj_out[2]
port 35 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 proj_out[30]
port 36 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 proj_out[31]
port 37 nsew signal input
rlabel metal3 s 0 11088 400 11144 6 proj_out[32]
port 38 nsew signal input
rlabel metal3 s 0 12096 400 12152 6 proj_out[33]
port 39 nsew signal input
rlabel metal3 s 0 12432 400 12488 6 proj_out[34]
port 40 nsew signal input
rlabel metal3 s 0 11760 400 11816 6 proj_out[35]
port 41 nsew signal input
rlabel metal3 s 19600 7392 20000 7448 6 proj_out[36]
port 42 nsew signal input
rlabel metal3 s 19600 8064 20000 8120 6 proj_out[37]
port 43 nsew signal input
rlabel metal2 s 11088 19600 11144 20000 6 proj_out[38]
port 44 nsew signal input
rlabel metal2 s 10752 19600 10808 20000 6 proj_out[39]
port 45 nsew signal input
rlabel metal3 s 19600 10416 20000 10472 6 proj_out[3]
port 46 nsew signal input
rlabel metal3 s 0 8064 400 8120 6 proj_out[40]
port 47 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 proj_out[41]
port 48 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 proj_out[42]
port 49 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 proj_out[43]
port 50 nsew signal input
rlabel metal3 s 0 10416 400 10472 6 proj_out[44]
port 51 nsew signal input
rlabel metal2 s 7728 19600 7784 20000 6 proj_out[45]
port 52 nsew signal input
rlabel metal3 s 0 9408 400 9464 6 proj_out[46]
port 53 nsew signal input
rlabel metal2 s 8064 19600 8120 20000 6 proj_out[47]
port 54 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 proj_out[4]
port 55 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 proj_out[5]
port 56 nsew signal input
rlabel metal2 s 10752 0 10808 400 6 proj_out[6]
port 57 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 proj_out[7]
port 58 nsew signal input
rlabel metal3 s 0 11424 400 11480 6 proj_out[8]
port 59 nsew signal input
rlabel metal2 s 9744 19600 9800 20000 6 proj_out[9]
port 60 nsew signal input
rlabel metal3 s 0 8736 400 8792 6 sel[0]
port 61 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 sel[1]
port 62 nsew signal input
rlabel metal4 s 2923 1538 3083 18454 6 vdd
port 63 nsew power bidirectional
rlabel metal4 s 7585 1538 7745 18454 6 vdd
port 63 nsew power bidirectional
rlabel metal4 s 12247 1538 12407 18454 6 vdd
port 63 nsew power bidirectional
rlabel metal4 s 16909 1538 17069 18454 6 vdd
port 63 nsew power bidirectional
rlabel metal4 s 5254 1538 5414 18454 6 vss
port 64 nsew ground bidirectional
rlabel metal4 s 9916 1538 10076 18454 6 vss
port 64 nsew ground bidirectional
rlabel metal4 s 14578 1538 14738 18454 6 vss
port 64 nsew ground bidirectional
rlabel metal4 s 19240 1538 19400 18454 6 vss
port 64 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 416262
string GDS_FILE /home/htamas/progs/gfmpw1-multi/openlane/output_mux/runs/23_12_12_04_50/results/signoff/output_mux.magic.gds
string GDS_START 74920
<< end >>

