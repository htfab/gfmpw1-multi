magic
tech gf180mcuD
magscale 1 5
timestamp 1702359423
<< obsm1 >>
rect 672 463 59304 58438
<< metal2 >>
rect 0 0 56 400
rect 12768 0 12824 400
rect 13104 0 13160 400
rect 13440 0 13496 400
rect 14112 0 14168 400
rect 14784 0 14840 400
rect 15456 0 15512 400
rect 18144 0 18200 400
rect 18480 0 18536 400
rect 20496 0 20552 400
rect 29568 0 29624 400
rect 35952 0 36008 400
rect 36288 0 36344 400
rect 36624 0 36680 400
rect 37296 0 37352 400
rect 37632 0 37688 400
rect 37968 0 38024 400
rect 38304 0 38360 400
rect 38640 0 38696 400
rect 38976 0 39032 400
rect 39312 0 39368 400
<< obsm2 >>
rect 854 430 59010 58427
rect 854 400 12738 430
rect 12854 400 13074 430
rect 13190 400 13410 430
rect 13526 400 14082 430
rect 14198 400 14754 430
rect 14870 400 15426 430
rect 15542 400 18114 430
rect 18230 400 18450 430
rect 18566 400 20466 430
rect 20582 400 29538 430
rect 29654 400 35922 430
rect 36038 400 36258 430
rect 36374 400 36594 430
rect 36710 400 37266 430
rect 37382 400 37602 430
rect 37718 400 37938 430
rect 38054 400 38274 430
rect 38390 400 38610 430
rect 38726 400 38946 430
rect 39062 400 39282 430
rect 39398 400 59010 430
<< metal3 >>
rect 59600 21504 60000 21560
rect 59600 21168 60000 21224
rect 59600 20832 60000 20888
rect 59600 20496 60000 20552
rect 59600 19488 60000 19544
rect 59600 19152 60000 19208
rect 0 18480 400 18536
rect 0 16464 400 16520
rect 0 16128 400 16184
rect 0 15792 400 15848
rect 0 15456 400 15512
rect 0 14784 400 14840
<< obsm3 >>
rect 400 21590 59600 58422
rect 400 21474 59570 21590
rect 400 21254 59600 21474
rect 400 21138 59570 21254
rect 400 20918 59600 21138
rect 400 20802 59570 20918
rect 400 20582 59600 20802
rect 400 20466 59570 20582
rect 400 19574 59600 20466
rect 400 19458 59570 19574
rect 400 19238 59600 19458
rect 400 19122 59570 19238
rect 400 18566 59600 19122
rect 430 18450 59600 18566
rect 400 16550 59600 18450
rect 430 16434 59600 16550
rect 400 16214 59600 16434
rect 430 16098 59600 16214
rect 400 15878 59600 16098
rect 430 15762 59600 15878
rect 400 15542 59600 15762
rect 430 15426 59600 15542
rect 400 14870 59600 15426
rect 430 14754 59600 14870
rect 400 1554 59600 14754
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
<< obsm4 >>
rect 17486 5665 17554 58119
rect 17774 5665 25234 58119
rect 25454 5665 32914 58119
rect 33134 5665 40594 58119
rect 40814 5665 45962 58119
<< labels >>
rlabel metal2 s 29568 0 29624 400 6 clk
port 1 nsew signal input
rlabel metal3 s 0 18480 400 18536 6 in[0]
port 2 nsew signal input
rlabel metal2 s 13440 0 13496 400 6 in[10]
port 3 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 in[11]
port 4 nsew signal input
rlabel metal2 s 36288 0 36344 400 6 in[12]
port 5 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 in[13]
port 6 nsew signal input
rlabel metal2 s 35952 0 36008 400 6 in[14]
port 7 nsew signal input
rlabel metal2 s 37296 0 37352 400 6 in[15]
port 8 nsew signal input
rlabel metal2 s 39312 0 39368 400 6 in[16]
port 9 nsew signal input
rlabel metal2 s 38976 0 39032 400 6 in[17]
port 10 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 in[18]
port 11 nsew signal input
rlabel metal3 s 0 16464 400 16520 6 in[1]
port 12 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 in[2]
port 13 nsew signal input
rlabel metal2 s 14784 0 14840 400 6 in[3]
port 14 nsew signal input
rlabel metal3 s 0 14784 400 14840 6 in[4]
port 15 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 in[5]
port 16 nsew signal input
rlabel metal3 s 0 15792 400 15848 6 in[6]
port 17 nsew signal input
rlabel metal3 s 0 16128 400 16184 6 in[7]
port 18 nsew signal input
rlabel metal3 s 0 15456 400 15512 6 in[8]
port 19 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 in[9]
port 20 nsew signal input
rlabel metal2 s 20496 0 20552 400 6 out[0]
port 21 nsew signal output
rlabel metal3 s 59600 19488 60000 19544 6 out[10]
port 22 nsew signal output
rlabel metal3 s 59600 19152 60000 19208 6 out[11]
port 23 nsew signal output
rlabel metal2 s 15456 0 15512 400 6 out[1]
port 24 nsew signal output
rlabel metal2 s 18144 0 18200 400 6 out[2]
port 25 nsew signal output
rlabel metal2 s 38640 0 38696 400 6 out[3]
port 26 nsew signal output
rlabel metal2 s 37632 0 37688 400 6 out[4]
port 27 nsew signal output
rlabel metal2 s 37968 0 38024 400 6 out[5]
port 28 nsew signal output
rlabel metal3 s 59600 21504 60000 21560 6 out[6]
port 29 nsew signal output
rlabel metal3 s 59600 21168 60000 21224 6 out[7]
port 30 nsew signal output
rlabel metal3 s 59600 20832 60000 20888 6 out[8]
port 31 nsew signal output
rlabel metal3 s 59600 20496 60000 20552 6 out[9]
port 32 nsew signal output
rlabel metal2 s 0 0 56 400 6 rst_n
port 33 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 35 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6047754
string GDS_FILE /home/htamas/test/caravel_user_project/openlane/unigate/runs/23_12_12_06_27/results/signoff/unigate.magic.gds
string GDS_START 469442
<< end >>

