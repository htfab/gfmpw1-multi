VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rotfpga2b
  CLASS BLOCK ;
  FOREIGN rotfpga2b ;
  ORIGIN 0.000 0.000 ;
  SIZE 1280.000 BY 1280.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END clk
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1186.080 4.000 1186.640 ;
    END
  END in[0]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 0.000 568.400 4.000 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 0.000 578.480 4.000 ;
    END
  END in[11]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 0.000 591.920 4.000 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 0.000 588.560 4.000 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 0.000 581.840 4.000 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 0.000 575.120 4.000 ;
    END
  END in[15]
  PIN in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 0.000 571.760 4.000 ;
    END
  END in[16]
  PIN in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END in[17]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 0.000 585.200 4.000 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 0.000 333.200 4.000 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 0.000 410.480 4.000 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1276.000 413.280 1280.000 413.840 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1276.000 588.000 1280.000 588.560 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 1276.000 780.080 1280.000 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 1276.000 763.280 1280.000 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 1276.000 518.000 1280.000 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 829.920 4.000 830.480 ;
    END
  END in[9]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1276.000 1075.200 1280.000 1075.760 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1276.000 1253.280 1280.000 1253.840 ;
    END
  END out[11]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 0.000 534.800 4.000 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1276.000 450.240 1280.000 450.800 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1276.000 608.160 1280.000 608.720 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 809.760 1276.000 810.320 1280.000 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 786.240 1276.000 786.800 1280.000 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 1276.000 534.800 1280.000 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 776.160 4.000 776.720 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 0.000 403.760 4.000 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 1276.000 904.400 1280.000 ;
    END
  END out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 0.000 7.280 4.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 1262.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1262.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1262.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1272.880 1263.210 ;
      LAYER Metal2 ;
        RECT 8.540 1275.700 517.140 1276.000 ;
        RECT 518.300 1275.700 533.940 1276.000 ;
        RECT 535.100 1275.700 762.420 1276.000 ;
        RECT 763.580 1275.700 779.220 1276.000 ;
        RECT 780.380 1275.700 785.940 1276.000 ;
        RECT 787.100 1275.700 809.460 1276.000 ;
        RECT 810.620 1275.700 903.540 1276.000 ;
        RECT 904.700 1275.700 1271.060 1276.000 ;
        RECT 8.540 4.300 1271.060 1275.700 ;
        RECT 8.540 3.450 332.340 4.300 ;
        RECT 333.500 3.450 386.100 4.300 ;
        RECT 387.260 3.450 402.900 4.300 ;
        RECT 404.060 3.450 409.620 4.300 ;
        RECT 410.780 3.450 533.940 4.300 ;
        RECT 535.100 3.450 567.540 4.300 ;
        RECT 568.700 3.450 570.900 4.300 ;
        RECT 572.060 3.450 574.260 4.300 ;
        RECT 575.420 3.450 577.620 4.300 ;
        RECT 578.780 3.450 580.980 4.300 ;
        RECT 582.140 3.450 584.340 4.300 ;
        RECT 585.500 3.450 587.700 4.300 ;
        RECT 588.860 3.450 591.060 4.300 ;
        RECT 592.220 3.450 1271.060 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1254.140 1276.000 1262.380 ;
        RECT 4.000 1252.980 1275.700 1254.140 ;
        RECT 4.000 1186.940 1276.000 1252.980 ;
        RECT 4.300 1185.780 1276.000 1186.940 ;
        RECT 4.000 1076.060 1276.000 1185.780 ;
        RECT 4.000 1074.900 1275.700 1076.060 ;
        RECT 4.000 830.780 1276.000 1074.900 ;
        RECT 4.300 829.620 1276.000 830.780 ;
        RECT 4.000 777.020 1276.000 829.620 ;
        RECT 4.300 775.860 1276.000 777.020 ;
        RECT 4.000 609.020 1276.000 775.860 ;
        RECT 4.000 607.860 1275.700 609.020 ;
        RECT 4.000 588.860 1276.000 607.860 ;
        RECT 4.000 587.700 1275.700 588.860 ;
        RECT 4.000 451.100 1276.000 587.700 ;
        RECT 4.000 449.940 1275.700 451.100 ;
        RECT 4.000 414.140 1276.000 449.940 ;
        RECT 4.000 412.980 1275.700 414.140 ;
        RECT 4.000 2.940 1276.000 412.980 ;
      LAYER Metal4 ;
        RECT 84.700 15.080 98.740 1261.030 ;
        RECT 100.940 15.080 175.540 1261.030 ;
        RECT 177.740 15.080 252.340 1261.030 ;
        RECT 254.540 15.080 329.140 1261.030 ;
        RECT 331.340 15.080 405.940 1261.030 ;
        RECT 408.140 15.080 482.740 1261.030 ;
        RECT 484.940 15.080 559.540 1261.030 ;
        RECT 561.740 15.080 636.340 1261.030 ;
        RECT 638.540 15.080 713.140 1261.030 ;
        RECT 715.340 15.080 789.940 1261.030 ;
        RECT 792.140 15.080 866.740 1261.030 ;
        RECT 868.940 15.080 943.540 1261.030 ;
        RECT 945.740 15.080 1020.340 1261.030 ;
        RECT 1022.540 15.080 1097.140 1261.030 ;
        RECT 1099.340 15.080 1173.940 1261.030 ;
        RECT 1176.140 15.080 1211.140 1261.030 ;
        RECT 84.700 2.890 1211.140 15.080 ;
  END
END rotfpga2b
END LIBRARY

