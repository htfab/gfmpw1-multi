magic
tech gf180mcuD
magscale 1 5
timestamp 1702353929
<< metal1 >>
rect 672 6285 7360 6302
rect 672 6259 2259 6285
rect 2285 6259 2311 6285
rect 2337 6259 2363 6285
rect 2389 6259 3911 6285
rect 3937 6259 3963 6285
rect 3989 6259 4015 6285
rect 4041 6259 5563 6285
rect 5589 6259 5615 6285
rect 5641 6259 5667 6285
rect 5693 6259 7215 6285
rect 7241 6259 7267 6285
rect 7293 6259 7319 6285
rect 7345 6259 7360 6285
rect 672 6242 7360 6259
rect 4047 6201 4073 6207
rect 4047 6169 4073 6175
rect 3431 6145 3457 6151
rect 3431 6113 3457 6119
rect 3711 6145 3737 6151
rect 3711 6113 3737 6119
rect 4215 6145 4241 6151
rect 4215 6113 4241 6119
rect 4383 6145 4409 6151
rect 4383 6113 4409 6119
rect 4831 6145 4857 6151
rect 5833 6119 5839 6145
rect 5865 6119 5871 6145
rect 4831 6113 4857 6119
rect 3593 6063 3599 6089
rect 3625 6063 3631 6089
rect 3929 6063 3935 6089
rect 3961 6063 3967 6089
rect 4713 6063 4719 6089
rect 4745 6063 4751 6089
rect 5217 6063 5223 6089
rect 5249 6063 5255 6089
rect 6785 6063 6791 6089
rect 6817 6063 6823 6089
rect 3207 6033 3233 6039
rect 3207 6001 3233 6007
rect 6567 6033 6593 6039
rect 6729 6007 6735 6033
rect 6761 6007 6767 6033
rect 6567 6001 6593 6007
rect 672 5893 7280 5910
rect 672 5867 1433 5893
rect 1459 5867 1485 5893
rect 1511 5867 1537 5893
rect 1563 5867 3085 5893
rect 3111 5867 3137 5893
rect 3163 5867 3189 5893
rect 3215 5867 4737 5893
rect 4763 5867 4789 5893
rect 4815 5867 4841 5893
rect 4867 5867 6389 5893
rect 6415 5867 6441 5893
rect 6467 5867 6493 5893
rect 6519 5867 7280 5893
rect 672 5850 7280 5867
rect 3543 5753 3569 5759
rect 3543 5721 3569 5727
rect 3767 5753 3793 5759
rect 6225 5727 6231 5753
rect 6257 5727 6263 5753
rect 6953 5727 6959 5753
rect 6985 5727 6991 5753
rect 3767 5721 3793 5727
rect 4321 5671 4327 5697
rect 4353 5671 4359 5697
rect 5217 5671 5223 5697
rect 5249 5671 5255 5697
rect 6785 5671 6791 5697
rect 6817 5671 6823 5697
rect 4041 5615 4047 5641
rect 4073 5615 4079 5641
rect 4881 5615 4887 5641
rect 4913 5615 4919 5641
rect 4825 5559 4831 5585
rect 4857 5559 4863 5585
rect 672 5501 7360 5518
rect 672 5475 2259 5501
rect 2285 5475 2311 5501
rect 2337 5475 2363 5501
rect 2389 5475 3911 5501
rect 3937 5475 3963 5501
rect 3989 5475 4015 5501
rect 4041 5475 5563 5501
rect 5589 5475 5615 5501
rect 5641 5475 5667 5501
rect 5693 5475 7215 5501
rect 7241 5475 7267 5501
rect 7293 5475 7319 5501
rect 7345 5475 7360 5501
rect 672 5458 7360 5475
rect 4215 5417 4241 5423
rect 4215 5385 4241 5391
rect 4775 5417 4801 5423
rect 4775 5385 4801 5391
rect 3991 5361 4017 5367
rect 3991 5329 4017 5335
rect 4327 5361 4353 5367
rect 4327 5329 4353 5335
rect 4495 5361 4521 5367
rect 4495 5329 4521 5335
rect 4943 5361 4969 5367
rect 6281 5335 6287 5361
rect 6313 5335 6319 5361
rect 4943 5329 4969 5335
rect 5273 5279 5279 5305
rect 5305 5279 5311 5305
rect 7009 5279 7015 5305
rect 7041 5279 7047 5305
rect 5615 5249 5641 5255
rect 5161 5223 5167 5249
rect 5193 5223 5199 5249
rect 5615 5217 5641 5223
rect 672 5109 7280 5126
rect 672 5083 1433 5109
rect 1459 5083 1485 5109
rect 1511 5083 1537 5109
rect 1563 5083 3085 5109
rect 3111 5083 3137 5109
rect 3163 5083 3189 5109
rect 3215 5083 4737 5109
rect 4763 5083 4789 5109
rect 4815 5083 4841 5109
rect 4867 5083 6389 5109
rect 6415 5083 6441 5109
rect 6467 5083 6493 5109
rect 6519 5083 7280 5109
rect 672 5066 7280 5083
rect 5833 4943 5839 4969
rect 5865 4943 5871 4969
rect 6953 4943 6959 4969
rect 6985 4943 6991 4969
rect 4265 4887 4271 4913
rect 4297 4887 4303 4913
rect 6281 4887 6287 4913
rect 6313 4887 6319 4913
rect 855 4857 881 4863
rect 4999 4857 5025 4863
rect 4209 4831 4215 4857
rect 4241 4831 4247 4857
rect 4881 4831 4887 4857
rect 4913 4831 4919 4857
rect 855 4825 881 4831
rect 4999 4825 5025 4831
rect 1023 4801 1049 4807
rect 1023 4769 1049 4775
rect 1247 4801 1273 4807
rect 1247 4769 1273 4775
rect 6735 4801 6761 4807
rect 6735 4769 6761 4775
rect 672 4717 7360 4734
rect 672 4691 2259 4717
rect 2285 4691 2311 4717
rect 2337 4691 2363 4717
rect 2389 4691 3911 4717
rect 3937 4691 3963 4717
rect 3989 4691 4015 4717
rect 4041 4691 5563 4717
rect 5589 4691 5615 4717
rect 5641 4691 5667 4717
rect 5693 4691 7215 4717
rect 7241 4691 7267 4717
rect 7293 4691 7319 4717
rect 7345 4691 7360 4717
rect 672 4674 7360 4691
rect 5447 4633 5473 4639
rect 5447 4601 5473 4607
rect 1023 4577 1049 4583
rect 1023 4545 1049 4551
rect 4495 4577 4521 4583
rect 4495 4545 4521 4551
rect 5615 4577 5641 4583
rect 6673 4551 6679 4577
rect 6705 4551 6711 4577
rect 5615 4545 5641 4551
rect 855 4521 881 4527
rect 4377 4495 4383 4521
rect 4409 4495 4415 4521
rect 4993 4495 4999 4521
rect 5025 4495 5031 4521
rect 5889 4495 5895 4521
rect 5921 4495 5927 4521
rect 855 4489 881 4495
rect 1247 4465 1273 4471
rect 1247 4433 1273 4439
rect 4775 4465 4801 4471
rect 5217 4439 5223 4465
rect 5249 4439 5255 4465
rect 4775 4433 4801 4439
rect 672 4325 7280 4342
rect 672 4299 1433 4325
rect 1459 4299 1485 4325
rect 1511 4299 1537 4325
rect 1563 4299 3085 4325
rect 3111 4299 3137 4325
rect 3163 4299 3189 4325
rect 3215 4299 4737 4325
rect 4763 4299 4789 4325
rect 4815 4299 4841 4325
rect 4867 4299 6389 4325
rect 6415 4299 6441 4325
rect 6467 4299 6493 4325
rect 6519 4299 7280 4325
rect 672 4282 7280 4299
rect 4999 4185 5025 4191
rect 4999 4153 5025 4159
rect 6343 4185 6369 4191
rect 6343 4153 6369 4159
rect 7015 4129 7041 4135
rect 1297 4103 1303 4129
rect 1329 4103 1335 4129
rect 4321 4103 4327 4129
rect 4353 4103 4359 4129
rect 5385 4103 5391 4129
rect 5417 4103 5423 4129
rect 6785 4103 6791 4129
rect 6817 4103 6823 4129
rect 7015 4097 7041 4103
rect 855 4073 881 4079
rect 855 4041 881 4047
rect 1807 4073 1833 4079
rect 4097 4047 4103 4073
rect 4129 4047 4135 4073
rect 4881 4047 4887 4073
rect 4913 4047 4919 4073
rect 1807 4041 1833 4047
rect 1023 4017 1049 4023
rect 1023 3985 1049 3991
rect 1191 4017 1217 4023
rect 1191 3985 1217 3991
rect 1583 4017 1609 4023
rect 1583 3985 1609 3991
rect 672 3933 7360 3950
rect 672 3907 2259 3933
rect 2285 3907 2311 3933
rect 2337 3907 2363 3933
rect 2389 3907 3911 3933
rect 3937 3907 3963 3933
rect 3989 3907 4015 3933
rect 4041 3907 5563 3933
rect 5589 3907 5615 3933
rect 5641 3907 5667 3933
rect 5693 3907 7215 3933
rect 7241 3907 7267 3933
rect 7293 3907 7319 3933
rect 7345 3907 7360 3933
rect 672 3890 7360 3907
rect 2529 3767 2535 3793
rect 2561 3767 2567 3793
rect 3313 3767 3319 3793
rect 3345 3767 3351 3793
rect 6617 3767 6623 3793
rect 6649 3767 6655 3793
rect 1185 3711 1191 3737
rect 1217 3711 1223 3737
rect 4153 3711 4159 3737
rect 4185 3711 4191 3737
rect 5161 3711 5167 3737
rect 5193 3711 5199 3737
rect 5889 3711 5895 3737
rect 5921 3711 5927 3737
rect 1527 3681 1553 3687
rect 1129 3655 1135 3681
rect 1161 3655 1167 3681
rect 1527 3649 1553 3655
rect 1751 3681 1777 3687
rect 1751 3649 1777 3655
rect 2479 3681 2505 3687
rect 2479 3649 2505 3655
rect 3487 3681 3513 3687
rect 3487 3649 3513 3655
rect 3823 3681 3849 3687
rect 5447 3681 5473 3687
rect 4265 3655 4271 3681
rect 4297 3655 4303 3681
rect 5217 3655 5223 3681
rect 5249 3655 5255 3681
rect 3823 3649 3849 3655
rect 5447 3649 5473 3655
rect 672 3541 7280 3558
rect 672 3515 1433 3541
rect 1459 3515 1485 3541
rect 1511 3515 1537 3541
rect 1563 3515 3085 3541
rect 3111 3515 3137 3541
rect 3163 3515 3189 3541
rect 3215 3515 4737 3541
rect 4763 3515 4789 3541
rect 4815 3515 4841 3541
rect 4867 3515 6389 3541
rect 6415 3515 6441 3541
rect 6467 3515 6493 3541
rect 6519 3515 7280 3541
rect 672 3498 7280 3515
rect 3319 3401 3345 3407
rect 1409 3375 1415 3401
rect 1441 3375 1447 3401
rect 2865 3375 2871 3401
rect 2897 3375 2903 3401
rect 3319 3369 3345 3375
rect 3991 3401 4017 3407
rect 6281 3375 6287 3401
rect 6313 3375 6319 3401
rect 3991 3369 4017 3375
rect 2479 3345 2505 3351
rect 905 3319 911 3345
rect 937 3319 943 3345
rect 2137 3319 2143 3345
rect 2169 3319 2175 3345
rect 2977 3319 2983 3345
rect 3009 3319 3015 3345
rect 3593 3319 3599 3345
rect 3625 3319 3631 3345
rect 5217 3319 5223 3345
rect 5249 3319 5255 3345
rect 2479 3313 2505 3319
rect 4999 3289 5025 3295
rect 1689 3263 1695 3289
rect 1721 3263 1727 3289
rect 4041 3263 4047 3289
rect 4073 3263 4079 3289
rect 4881 3263 4887 3289
rect 4913 3263 4919 3289
rect 4999 3257 5025 3263
rect 6735 3289 6761 3295
rect 6735 3257 6761 3263
rect 6903 3289 6929 3295
rect 6903 3257 6929 3263
rect 1023 3233 1049 3239
rect 1023 3201 1049 3207
rect 3711 3233 3737 3239
rect 3711 3201 3737 3207
rect 672 3149 7360 3166
rect 672 3123 2259 3149
rect 2285 3123 2311 3149
rect 2337 3123 2363 3149
rect 2389 3123 3911 3149
rect 3937 3123 3963 3149
rect 3989 3123 4015 3149
rect 4041 3123 5563 3149
rect 5589 3123 5615 3149
rect 5641 3123 5667 3149
rect 5693 3123 7215 3149
rect 7241 3123 7267 3149
rect 7293 3123 7319 3149
rect 7345 3123 7360 3149
rect 672 3106 7360 3123
rect 1801 3039 1807 3065
rect 1833 3039 1839 3065
rect 2143 3009 2169 3015
rect 5447 3009 5473 3015
rect 1073 2983 1079 3009
rect 1105 2983 1111 3009
rect 3649 2983 3655 3009
rect 3681 2983 3687 3009
rect 2143 2977 2169 2983
rect 5447 2977 5473 2983
rect 5615 3009 5641 3015
rect 6673 2983 6679 3009
rect 6705 2983 6711 3009
rect 5615 2977 5641 2983
rect 2199 2953 2225 2959
rect 4495 2953 4521 2959
rect 1633 2927 1639 2953
rect 1665 2927 1671 2953
rect 2361 2927 2367 2953
rect 2393 2927 2399 2953
rect 3817 2927 3823 2953
rect 3849 2927 3855 2953
rect 4265 2927 4271 2953
rect 4297 2927 4303 2953
rect 2199 2921 2225 2927
rect 4495 2921 4521 2927
rect 4943 2953 4969 2959
rect 4943 2921 4969 2927
rect 5223 2953 5249 2959
rect 5777 2927 5783 2953
rect 5809 2927 5815 2953
rect 5223 2921 5249 2927
rect 967 2897 993 2903
rect 967 2865 993 2871
rect 672 2757 7280 2774
rect 672 2731 1433 2757
rect 1459 2731 1485 2757
rect 1511 2731 1537 2757
rect 1563 2731 3085 2757
rect 3111 2731 3137 2757
rect 3163 2731 3189 2757
rect 3215 2731 4737 2757
rect 4763 2731 4789 2757
rect 4815 2731 4841 2757
rect 4867 2731 6389 2757
rect 6415 2731 6441 2757
rect 6467 2731 6493 2757
rect 6519 2731 7280 2757
rect 672 2714 7280 2731
rect 1807 2617 1833 2623
rect 1807 2585 1833 2591
rect 855 2561 881 2567
rect 855 2529 881 2535
rect 1191 2561 1217 2567
rect 1191 2529 1217 2535
rect 1583 2561 1609 2567
rect 1583 2529 1609 2535
rect 3655 2561 3681 2567
rect 3655 2529 3681 2535
rect 3935 2561 3961 2567
rect 3935 2529 3961 2535
rect 6455 2561 6481 2567
rect 6455 2529 6481 2535
rect 6903 2561 6929 2567
rect 6903 2529 6929 2535
rect 1023 2505 1049 2511
rect 1023 2473 1049 2479
rect 1359 2505 1385 2511
rect 1359 2473 1385 2479
rect 6287 2505 6313 2511
rect 6287 2473 6313 2479
rect 6735 2505 6761 2511
rect 6735 2473 6761 2479
rect 672 2365 7360 2382
rect 672 2339 2259 2365
rect 2285 2339 2311 2365
rect 2337 2339 2363 2365
rect 2389 2339 3911 2365
rect 3937 2339 3963 2365
rect 3989 2339 4015 2365
rect 4041 2339 5563 2365
rect 5589 2339 5615 2365
rect 5641 2339 5667 2365
rect 5693 2339 7215 2365
rect 7241 2339 7267 2365
rect 7293 2339 7319 2365
rect 7345 2339 7360 2365
rect 672 2322 7360 2339
rect 1023 2281 1049 2287
rect 1023 2249 1049 2255
rect 1359 2281 1385 2287
rect 1359 2249 1385 2255
rect 6623 2281 6649 2287
rect 6623 2249 6649 2255
rect 6903 2281 6929 2287
rect 6903 2249 6929 2255
rect 855 2225 881 2231
rect 7071 2225 7097 2231
rect 3425 2199 3431 2225
rect 3457 2199 3463 2225
rect 855 2193 881 2199
rect 7071 2193 7097 2199
rect 1191 2169 1217 2175
rect 1191 2137 1217 2143
rect 3263 2169 3289 2175
rect 4769 2143 4775 2169
rect 4801 2143 4807 2169
rect 3263 2137 3289 2143
rect 1583 2113 1609 2119
rect 1583 2081 1609 2087
rect 3095 2113 3121 2119
rect 3095 2081 3121 2087
rect 4047 2113 4073 2119
rect 4047 2081 4073 2087
rect 5279 2057 5305 2063
rect 5279 2025 5305 2031
rect 672 1973 7280 1990
rect 672 1947 1433 1973
rect 1459 1947 1485 1973
rect 1511 1947 1537 1973
rect 1563 1947 3085 1973
rect 3111 1947 3137 1973
rect 3163 1947 3189 1973
rect 3215 1947 4737 1973
rect 4763 1947 4789 1973
rect 4815 1947 4841 1973
rect 4867 1947 6389 1973
rect 6415 1947 6441 1973
rect 6467 1947 6493 1973
rect 6519 1947 7280 1973
rect 672 1930 7280 1947
rect 1247 1833 1273 1839
rect 1247 1801 1273 1807
rect 5335 1833 5361 1839
rect 5335 1801 5361 1807
rect 7127 1833 7153 1839
rect 7127 1801 7153 1807
rect 3375 1777 3401 1783
rect 3593 1751 3599 1777
rect 3625 1751 3631 1777
rect 3929 1751 3935 1777
rect 3961 1751 3967 1777
rect 4265 1751 4271 1777
rect 4297 1751 4303 1777
rect 4937 1751 4943 1777
rect 4969 1751 4975 1777
rect 3375 1745 3401 1751
rect 855 1721 881 1727
rect 855 1689 881 1695
rect 1023 1721 1049 1727
rect 1023 1689 1049 1695
rect 1471 1721 1497 1727
rect 1471 1689 1497 1695
rect 3823 1721 3849 1727
rect 3823 1689 3849 1695
rect 4159 1721 4185 1727
rect 4159 1689 4185 1695
rect 3481 1639 3487 1665
rect 3513 1639 3519 1665
rect 672 1581 7360 1598
rect 672 1555 2259 1581
rect 2285 1555 2311 1581
rect 2337 1555 2363 1581
rect 2389 1555 3911 1581
rect 3937 1555 3963 1581
rect 3989 1555 4015 1581
rect 4041 1555 5563 1581
rect 5589 1555 5615 1581
rect 5641 1555 5667 1581
rect 5693 1555 7215 1581
rect 7241 1555 7267 1581
rect 7293 1555 7319 1581
rect 7345 1555 7360 1581
rect 672 1538 7360 1555
<< via1 >>
rect 2259 6259 2285 6285
rect 2311 6259 2337 6285
rect 2363 6259 2389 6285
rect 3911 6259 3937 6285
rect 3963 6259 3989 6285
rect 4015 6259 4041 6285
rect 5563 6259 5589 6285
rect 5615 6259 5641 6285
rect 5667 6259 5693 6285
rect 7215 6259 7241 6285
rect 7267 6259 7293 6285
rect 7319 6259 7345 6285
rect 4047 6175 4073 6201
rect 3431 6119 3457 6145
rect 3711 6119 3737 6145
rect 4215 6119 4241 6145
rect 4383 6119 4409 6145
rect 4831 6119 4857 6145
rect 5839 6119 5865 6145
rect 3599 6063 3625 6089
rect 3935 6063 3961 6089
rect 4719 6063 4745 6089
rect 5223 6063 5249 6089
rect 6791 6063 6817 6089
rect 3207 6007 3233 6033
rect 6567 6007 6593 6033
rect 6735 6007 6761 6033
rect 1433 5867 1459 5893
rect 1485 5867 1511 5893
rect 1537 5867 1563 5893
rect 3085 5867 3111 5893
rect 3137 5867 3163 5893
rect 3189 5867 3215 5893
rect 4737 5867 4763 5893
rect 4789 5867 4815 5893
rect 4841 5867 4867 5893
rect 6389 5867 6415 5893
rect 6441 5867 6467 5893
rect 6493 5867 6519 5893
rect 3543 5727 3569 5753
rect 3767 5727 3793 5753
rect 6231 5727 6257 5753
rect 6959 5727 6985 5753
rect 4327 5671 4353 5697
rect 5223 5671 5249 5697
rect 6791 5671 6817 5697
rect 4047 5615 4073 5641
rect 4887 5615 4913 5641
rect 4831 5559 4857 5585
rect 2259 5475 2285 5501
rect 2311 5475 2337 5501
rect 2363 5475 2389 5501
rect 3911 5475 3937 5501
rect 3963 5475 3989 5501
rect 4015 5475 4041 5501
rect 5563 5475 5589 5501
rect 5615 5475 5641 5501
rect 5667 5475 5693 5501
rect 7215 5475 7241 5501
rect 7267 5475 7293 5501
rect 7319 5475 7345 5501
rect 4215 5391 4241 5417
rect 4775 5391 4801 5417
rect 3991 5335 4017 5361
rect 4327 5335 4353 5361
rect 4495 5335 4521 5361
rect 4943 5335 4969 5361
rect 6287 5335 6313 5361
rect 5279 5279 5305 5305
rect 7015 5279 7041 5305
rect 5167 5223 5193 5249
rect 5615 5223 5641 5249
rect 1433 5083 1459 5109
rect 1485 5083 1511 5109
rect 1537 5083 1563 5109
rect 3085 5083 3111 5109
rect 3137 5083 3163 5109
rect 3189 5083 3215 5109
rect 4737 5083 4763 5109
rect 4789 5083 4815 5109
rect 4841 5083 4867 5109
rect 6389 5083 6415 5109
rect 6441 5083 6467 5109
rect 6493 5083 6519 5109
rect 5839 4943 5865 4969
rect 6959 4943 6985 4969
rect 4271 4887 4297 4913
rect 6287 4887 6313 4913
rect 855 4831 881 4857
rect 4215 4831 4241 4857
rect 4887 4831 4913 4857
rect 4999 4831 5025 4857
rect 1023 4775 1049 4801
rect 1247 4775 1273 4801
rect 6735 4775 6761 4801
rect 2259 4691 2285 4717
rect 2311 4691 2337 4717
rect 2363 4691 2389 4717
rect 3911 4691 3937 4717
rect 3963 4691 3989 4717
rect 4015 4691 4041 4717
rect 5563 4691 5589 4717
rect 5615 4691 5641 4717
rect 5667 4691 5693 4717
rect 7215 4691 7241 4717
rect 7267 4691 7293 4717
rect 7319 4691 7345 4717
rect 5447 4607 5473 4633
rect 1023 4551 1049 4577
rect 4495 4551 4521 4577
rect 5615 4551 5641 4577
rect 6679 4551 6705 4577
rect 855 4495 881 4521
rect 4383 4495 4409 4521
rect 4999 4495 5025 4521
rect 5895 4495 5921 4521
rect 1247 4439 1273 4465
rect 4775 4439 4801 4465
rect 5223 4439 5249 4465
rect 1433 4299 1459 4325
rect 1485 4299 1511 4325
rect 1537 4299 1563 4325
rect 3085 4299 3111 4325
rect 3137 4299 3163 4325
rect 3189 4299 3215 4325
rect 4737 4299 4763 4325
rect 4789 4299 4815 4325
rect 4841 4299 4867 4325
rect 6389 4299 6415 4325
rect 6441 4299 6467 4325
rect 6493 4299 6519 4325
rect 4999 4159 5025 4185
rect 6343 4159 6369 4185
rect 1303 4103 1329 4129
rect 4327 4103 4353 4129
rect 5391 4103 5417 4129
rect 6791 4103 6817 4129
rect 7015 4103 7041 4129
rect 855 4047 881 4073
rect 1807 4047 1833 4073
rect 4103 4047 4129 4073
rect 4887 4047 4913 4073
rect 1023 3991 1049 4017
rect 1191 3991 1217 4017
rect 1583 3991 1609 4017
rect 2259 3907 2285 3933
rect 2311 3907 2337 3933
rect 2363 3907 2389 3933
rect 3911 3907 3937 3933
rect 3963 3907 3989 3933
rect 4015 3907 4041 3933
rect 5563 3907 5589 3933
rect 5615 3907 5641 3933
rect 5667 3907 5693 3933
rect 7215 3907 7241 3933
rect 7267 3907 7293 3933
rect 7319 3907 7345 3933
rect 2535 3767 2561 3793
rect 3319 3767 3345 3793
rect 6623 3767 6649 3793
rect 1191 3711 1217 3737
rect 4159 3711 4185 3737
rect 5167 3711 5193 3737
rect 5895 3711 5921 3737
rect 1135 3655 1161 3681
rect 1527 3655 1553 3681
rect 1751 3655 1777 3681
rect 2479 3655 2505 3681
rect 3487 3655 3513 3681
rect 3823 3655 3849 3681
rect 4271 3655 4297 3681
rect 5223 3655 5249 3681
rect 5447 3655 5473 3681
rect 1433 3515 1459 3541
rect 1485 3515 1511 3541
rect 1537 3515 1563 3541
rect 3085 3515 3111 3541
rect 3137 3515 3163 3541
rect 3189 3515 3215 3541
rect 4737 3515 4763 3541
rect 4789 3515 4815 3541
rect 4841 3515 4867 3541
rect 6389 3515 6415 3541
rect 6441 3515 6467 3541
rect 6493 3515 6519 3541
rect 1415 3375 1441 3401
rect 2871 3375 2897 3401
rect 3319 3375 3345 3401
rect 3991 3375 4017 3401
rect 6287 3375 6313 3401
rect 911 3319 937 3345
rect 2143 3319 2169 3345
rect 2479 3319 2505 3345
rect 2983 3319 3009 3345
rect 3599 3319 3625 3345
rect 5223 3319 5249 3345
rect 1695 3263 1721 3289
rect 4047 3263 4073 3289
rect 4887 3263 4913 3289
rect 4999 3263 5025 3289
rect 6735 3263 6761 3289
rect 6903 3263 6929 3289
rect 1023 3207 1049 3233
rect 3711 3207 3737 3233
rect 2259 3123 2285 3149
rect 2311 3123 2337 3149
rect 2363 3123 2389 3149
rect 3911 3123 3937 3149
rect 3963 3123 3989 3149
rect 4015 3123 4041 3149
rect 5563 3123 5589 3149
rect 5615 3123 5641 3149
rect 5667 3123 5693 3149
rect 7215 3123 7241 3149
rect 7267 3123 7293 3149
rect 7319 3123 7345 3149
rect 1807 3039 1833 3065
rect 1079 2983 1105 3009
rect 2143 2983 2169 3009
rect 3655 2983 3681 3009
rect 5447 2983 5473 3009
rect 5615 2983 5641 3009
rect 6679 2983 6705 3009
rect 1639 2927 1665 2953
rect 2199 2927 2225 2953
rect 2367 2927 2393 2953
rect 3823 2927 3849 2953
rect 4271 2927 4297 2953
rect 4495 2927 4521 2953
rect 4943 2927 4969 2953
rect 5223 2927 5249 2953
rect 5783 2927 5809 2953
rect 967 2871 993 2897
rect 1433 2731 1459 2757
rect 1485 2731 1511 2757
rect 1537 2731 1563 2757
rect 3085 2731 3111 2757
rect 3137 2731 3163 2757
rect 3189 2731 3215 2757
rect 4737 2731 4763 2757
rect 4789 2731 4815 2757
rect 4841 2731 4867 2757
rect 6389 2731 6415 2757
rect 6441 2731 6467 2757
rect 6493 2731 6519 2757
rect 1807 2591 1833 2617
rect 855 2535 881 2561
rect 1191 2535 1217 2561
rect 1583 2535 1609 2561
rect 3655 2535 3681 2561
rect 3935 2535 3961 2561
rect 6455 2535 6481 2561
rect 6903 2535 6929 2561
rect 1023 2479 1049 2505
rect 1359 2479 1385 2505
rect 6287 2479 6313 2505
rect 6735 2479 6761 2505
rect 2259 2339 2285 2365
rect 2311 2339 2337 2365
rect 2363 2339 2389 2365
rect 3911 2339 3937 2365
rect 3963 2339 3989 2365
rect 4015 2339 4041 2365
rect 5563 2339 5589 2365
rect 5615 2339 5641 2365
rect 5667 2339 5693 2365
rect 7215 2339 7241 2365
rect 7267 2339 7293 2365
rect 7319 2339 7345 2365
rect 1023 2255 1049 2281
rect 1359 2255 1385 2281
rect 6623 2255 6649 2281
rect 6903 2255 6929 2281
rect 855 2199 881 2225
rect 3431 2199 3457 2225
rect 7071 2199 7097 2225
rect 1191 2143 1217 2169
rect 3263 2143 3289 2169
rect 4775 2143 4801 2169
rect 1583 2087 1609 2113
rect 3095 2087 3121 2113
rect 4047 2087 4073 2113
rect 5279 2031 5305 2057
rect 1433 1947 1459 1973
rect 1485 1947 1511 1973
rect 1537 1947 1563 1973
rect 3085 1947 3111 1973
rect 3137 1947 3163 1973
rect 3189 1947 3215 1973
rect 4737 1947 4763 1973
rect 4789 1947 4815 1973
rect 4841 1947 4867 1973
rect 6389 1947 6415 1973
rect 6441 1947 6467 1973
rect 6493 1947 6519 1973
rect 1247 1807 1273 1833
rect 5335 1807 5361 1833
rect 7127 1807 7153 1833
rect 3375 1751 3401 1777
rect 3599 1751 3625 1777
rect 3935 1751 3961 1777
rect 4271 1751 4297 1777
rect 4943 1751 4969 1777
rect 855 1695 881 1721
rect 1023 1695 1049 1721
rect 1471 1695 1497 1721
rect 3823 1695 3849 1721
rect 4159 1695 4185 1721
rect 3487 1639 3513 1665
rect 2259 1555 2285 1581
rect 2311 1555 2337 1581
rect 2363 1555 2389 1581
rect 3911 1555 3937 1581
rect 3963 1555 3989 1581
rect 4015 1555 4041 1581
rect 5563 1555 5589 1581
rect 5615 1555 5641 1581
rect 5667 1555 5693 1581
rect 7215 1555 7241 1581
rect 7267 1555 7293 1581
rect 7319 1555 7345 1581
<< metal2 >>
rect 4368 7600 4424 8000
rect 4704 7600 4760 8000
rect 5712 7600 5768 8000
rect 3598 7098 3626 7103
rect 2258 6286 2390 6291
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2258 6253 2390 6258
rect 3430 6146 3458 6151
rect 3430 6099 3458 6118
rect 3598 6089 3626 7070
rect 3910 6286 4042 6291
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 3910 6253 4042 6258
rect 4046 6202 4074 6207
rect 3598 6063 3599 6089
rect 3625 6063 3626 6089
rect 3206 6033 3234 6039
rect 3206 6007 3207 6033
rect 3233 6007 3234 6033
rect 3206 5978 3234 6007
rect 3206 5945 3234 5950
rect 1432 5894 1564 5899
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1432 5861 1564 5866
rect 3084 5894 3216 5899
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3084 5861 3216 5866
rect 3542 5754 3570 5759
rect 3598 5754 3626 6063
rect 3542 5753 3626 5754
rect 3542 5727 3543 5753
rect 3569 5727 3626 5753
rect 3542 5726 3626 5727
rect 3710 6145 3738 6151
rect 3710 6119 3711 6145
rect 3737 6119 3738 6145
rect 3542 5721 3570 5726
rect 2258 5502 2390 5507
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2258 5469 2390 5474
rect 3710 5250 3738 6119
rect 3766 6090 3794 6095
rect 3766 5753 3794 6062
rect 3934 6089 3962 6095
rect 3934 6063 3935 6089
rect 3961 6063 3962 6089
rect 3934 5978 3962 6063
rect 3934 5945 3962 5950
rect 3766 5727 3767 5753
rect 3793 5727 3794 5753
rect 3766 5721 3794 5727
rect 4046 5641 4074 6174
rect 4214 6146 4242 6151
rect 4382 6146 4410 7600
rect 4214 6145 4298 6146
rect 4214 6119 4215 6145
rect 4241 6119 4298 6145
rect 4214 6118 4298 6119
rect 4214 6113 4242 6118
rect 4046 5615 4047 5641
rect 4073 5615 4074 5641
rect 4046 5609 4074 5615
rect 3910 5502 4042 5507
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 3910 5469 4042 5474
rect 4214 5418 4242 5423
rect 4214 5371 4242 5390
rect 3990 5362 4018 5367
rect 3990 5315 4018 5334
rect 3710 5217 3738 5222
rect 4046 5250 4074 5255
rect 4074 5222 4130 5250
rect 4046 5217 4074 5222
rect 1432 5110 1564 5115
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1432 5077 1564 5082
rect 3084 5110 3216 5115
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3084 5077 3216 5082
rect 854 4857 882 4863
rect 854 4831 855 4857
rect 881 4831 882 4857
rect 854 4746 882 4831
rect 1022 4802 1050 4807
rect 1022 4801 1106 4802
rect 1022 4775 1023 4801
rect 1049 4775 1106 4801
rect 1022 4774 1106 4775
rect 1022 4769 1050 4774
rect 854 4713 882 4718
rect 1022 4577 1050 4583
rect 1022 4551 1023 4577
rect 1049 4551 1050 4577
rect 854 4521 882 4527
rect 854 4495 855 4521
rect 881 4495 882 4521
rect 854 4410 882 4495
rect 854 4377 882 4382
rect 1022 4214 1050 4551
rect 966 4186 1050 4214
rect 854 4074 882 4079
rect 854 4027 882 4046
rect 910 3682 938 3687
rect 910 3402 938 3654
rect 910 3345 938 3374
rect 910 3319 911 3345
rect 937 3319 938 3345
rect 910 3313 938 3319
rect 854 3066 882 3071
rect 854 2618 882 3038
rect 966 2897 994 4186
rect 1022 4017 1050 4023
rect 1022 3991 1023 4017
rect 1049 3991 1050 4017
rect 1022 3570 1050 3991
rect 1078 3794 1106 4774
rect 1246 4801 1274 4807
rect 1246 4775 1247 4801
rect 1273 4775 1274 4801
rect 1246 4746 1274 4775
rect 1246 4713 1274 4718
rect 2258 4718 2390 4723
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2258 4685 2390 4690
rect 3910 4718 4042 4723
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 3910 4685 4042 4690
rect 1246 4465 1274 4471
rect 1246 4439 1247 4465
rect 1273 4439 1274 4465
rect 1246 4410 1274 4439
rect 1246 4377 1274 4382
rect 1432 4326 1564 4331
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1432 4293 1564 4298
rect 3084 4326 3216 4331
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3084 4293 3216 4298
rect 1302 4129 1330 4135
rect 1302 4103 1303 4129
rect 1329 4103 1330 4129
rect 1190 4018 1218 4023
rect 1078 3761 1106 3766
rect 1134 4017 1218 4018
rect 1134 3991 1191 4017
rect 1217 3991 1218 4017
rect 1134 3990 1218 3991
rect 1134 3681 1162 3990
rect 1190 3985 1218 3990
rect 1302 4018 1330 4103
rect 1806 4074 1834 4079
rect 1806 4027 1834 4046
rect 4102 4073 4130 5222
rect 4270 4913 4298 6118
rect 4382 6099 4410 6118
rect 4718 6090 4746 7600
rect 5562 6286 5694 6291
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5562 6253 5694 6258
rect 4830 6146 4858 6151
rect 4830 6145 5026 6146
rect 4830 6119 4831 6145
rect 4857 6119 5026 6145
rect 4830 6118 5026 6119
rect 4830 6113 4858 6118
rect 4718 6043 4746 6062
rect 4736 5894 4868 5899
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4736 5861 4868 5866
rect 4326 5698 4354 5703
rect 4326 5651 4354 5670
rect 4774 5698 4802 5703
rect 4494 5418 4522 5423
rect 4270 4887 4271 4913
rect 4297 4887 4298 4913
rect 4270 4881 4298 4887
rect 4326 5361 4354 5367
rect 4326 5335 4327 5361
rect 4353 5335 4354 5361
rect 4214 4858 4242 4863
rect 4214 4811 4242 4830
rect 4326 4129 4354 5335
rect 4494 5361 4522 5390
rect 4774 5417 4802 5670
rect 4886 5698 4914 5703
rect 4886 5641 4914 5670
rect 4886 5615 4887 5641
rect 4913 5615 4914 5641
rect 4886 5609 4914 5615
rect 4774 5391 4775 5417
rect 4801 5391 4802 5417
rect 4774 5385 4802 5391
rect 4830 5585 4858 5591
rect 4830 5559 4831 5585
rect 4857 5559 4858 5585
rect 4494 5335 4495 5361
rect 4521 5335 4522 5361
rect 4494 5329 4522 5335
rect 4830 5194 4858 5559
rect 4942 5362 4970 5367
rect 4942 5315 4970 5334
rect 4662 5166 4858 5194
rect 4494 4577 4522 4583
rect 4494 4551 4495 4577
rect 4521 4551 4522 4577
rect 4382 4522 4410 4527
rect 4382 4475 4410 4494
rect 4326 4103 4327 4129
rect 4353 4103 4354 4129
rect 4326 4097 4354 4103
rect 4102 4047 4103 4073
rect 4129 4047 4130 4073
rect 4102 4041 4130 4047
rect 1582 4018 1610 4023
rect 1302 4017 1610 4018
rect 1302 3991 1583 4017
rect 1609 3991 1610 4017
rect 1302 3990 1610 3991
rect 1134 3655 1135 3681
rect 1161 3655 1162 3681
rect 1134 3649 1162 3655
rect 1190 3737 1218 3743
rect 1190 3711 1191 3737
rect 1217 3711 1218 3737
rect 1022 3542 1106 3570
rect 1078 3346 1106 3542
rect 1190 3402 1218 3711
rect 1302 3738 1330 3990
rect 1582 3985 1610 3990
rect 2258 3934 2390 3939
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2258 3901 2390 3906
rect 3910 3934 4042 3939
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 3910 3901 4042 3906
rect 1302 3705 1330 3710
rect 2534 3793 2562 3799
rect 2534 3767 2535 3793
rect 2561 3767 2562 3793
rect 1526 3681 1554 3687
rect 1526 3655 1527 3681
rect 1553 3655 1554 3681
rect 1526 3626 1554 3655
rect 1750 3682 1778 3687
rect 1750 3635 1778 3654
rect 2478 3681 2506 3687
rect 2478 3655 2479 3681
rect 2505 3655 2506 3681
rect 1078 3313 1106 3318
rect 1134 3374 1218 3402
rect 1358 3598 1554 3626
rect 1358 3402 1386 3598
rect 1432 3542 1564 3547
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1432 3509 1564 3514
rect 1414 3402 1442 3407
rect 1358 3401 1442 3402
rect 1358 3375 1415 3401
rect 1441 3375 1442 3401
rect 1358 3374 1442 3375
rect 1022 3234 1050 3239
rect 1134 3234 1162 3374
rect 1414 3369 1442 3374
rect 2142 3345 2170 3351
rect 2142 3319 2143 3345
rect 2169 3319 2170 3345
rect 1694 3290 1722 3295
rect 1694 3289 1834 3290
rect 1694 3263 1695 3289
rect 1721 3263 1834 3289
rect 1694 3262 1834 3263
rect 1694 3257 1722 3262
rect 1022 3233 1162 3234
rect 1022 3207 1023 3233
rect 1049 3207 1162 3233
rect 1022 3206 1162 3207
rect 1022 3201 1050 3206
rect 1806 3065 1834 3262
rect 1806 3039 1807 3065
rect 1833 3039 1834 3065
rect 1806 3033 1834 3039
rect 1078 3009 1106 3015
rect 1078 2983 1079 3009
rect 1105 2983 1106 3009
rect 966 2871 967 2897
rect 993 2871 994 2897
rect 966 2865 994 2871
rect 1022 2954 1050 2959
rect 854 2561 882 2590
rect 854 2535 855 2561
rect 881 2535 882 2561
rect 854 2529 882 2535
rect 966 2674 994 2679
rect 854 2394 882 2399
rect 854 2225 882 2366
rect 966 2282 994 2646
rect 1022 2505 1050 2926
rect 1022 2479 1023 2505
rect 1049 2479 1050 2505
rect 1022 2473 1050 2479
rect 1022 2282 1050 2287
rect 966 2281 1050 2282
rect 966 2255 1023 2281
rect 1049 2255 1050 2281
rect 966 2254 1050 2255
rect 1022 2249 1050 2254
rect 854 2199 855 2225
rect 881 2199 882 2225
rect 854 2193 882 2199
rect 854 1722 882 1727
rect 854 1675 882 1694
rect 1022 1722 1050 1727
rect 1078 1722 1106 2983
rect 2142 3009 2170 3319
rect 2142 2983 2143 3009
rect 2169 2983 2170 3009
rect 2142 2977 2170 2983
rect 2198 3346 2226 3351
rect 1638 2954 1666 2959
rect 1358 2953 1666 2954
rect 1358 2927 1639 2953
rect 1665 2927 1666 2953
rect 1358 2926 1666 2927
rect 1190 2730 1218 2735
rect 1190 2562 1218 2702
rect 1190 2515 1218 2534
rect 1358 2505 1386 2926
rect 1638 2921 1666 2926
rect 2198 2953 2226 3318
rect 2478 3345 2506 3655
rect 2478 3319 2479 3345
rect 2505 3319 2506 3345
rect 2478 3313 2506 3319
rect 2258 3150 2390 3155
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2258 3117 2390 3122
rect 2198 2927 2199 2953
rect 2225 2927 2226 2953
rect 2198 2921 2226 2927
rect 2366 2954 2394 2959
rect 2366 2907 2394 2926
rect 1432 2758 1564 2763
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1432 2725 1564 2730
rect 1806 2618 1834 2623
rect 1806 2571 1834 2590
rect 1582 2562 1610 2567
rect 1582 2515 1610 2534
rect 1358 2479 1359 2505
rect 1385 2479 1386 2505
rect 1358 2473 1386 2479
rect 1246 2394 1274 2399
rect 1190 2169 1218 2175
rect 1190 2143 1191 2169
rect 1217 2143 1218 2169
rect 1190 2058 1218 2143
rect 1190 2025 1218 2030
rect 1246 1833 1274 2366
rect 2258 2366 2390 2371
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2258 2333 2390 2338
rect 1358 2282 1386 2287
rect 1358 2235 1386 2254
rect 2534 2282 2562 3767
rect 2870 3794 2898 3799
rect 2870 3401 2898 3766
rect 3318 3793 3346 3799
rect 3318 3767 3319 3793
rect 3345 3767 3346 3793
rect 3084 3542 3216 3547
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3084 3509 3216 3514
rect 2870 3375 2871 3401
rect 2897 3375 2898 3401
rect 2870 3369 2898 3375
rect 3318 3401 3346 3767
rect 4158 3737 4186 3743
rect 4158 3711 4159 3737
rect 4185 3711 4186 3737
rect 3318 3375 3319 3401
rect 3345 3375 3346 3401
rect 3318 3369 3346 3375
rect 3486 3681 3514 3687
rect 3822 3682 3850 3687
rect 3486 3655 3487 3681
rect 3513 3655 3514 3681
rect 2982 3345 3010 3351
rect 2982 3319 2983 3345
rect 3009 3319 3010 3345
rect 2982 2674 3010 3319
rect 3084 2758 3216 2763
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3084 2725 3216 2730
rect 2982 2641 3010 2646
rect 3486 2562 3514 3655
rect 3598 3681 3850 3682
rect 3598 3655 3823 3681
rect 3849 3655 3850 3681
rect 3598 3654 3850 3655
rect 3598 3345 3626 3654
rect 3822 3649 3850 3654
rect 3990 3402 4018 3407
rect 3990 3401 4130 3402
rect 3990 3375 3991 3401
rect 4017 3375 4130 3401
rect 3990 3374 4130 3375
rect 3990 3369 4018 3374
rect 3598 3319 3599 3345
rect 3625 3319 3626 3345
rect 3598 3313 3626 3319
rect 4046 3289 4074 3295
rect 4046 3263 4047 3289
rect 4073 3263 4074 3289
rect 3710 3233 3738 3239
rect 3710 3207 3711 3233
rect 3737 3207 3738 3233
rect 3654 3010 3682 3015
rect 3654 2963 3682 2982
rect 3710 2674 3738 3207
rect 4046 3234 4074 3263
rect 4046 3201 4074 3206
rect 3910 3150 4042 3155
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 3910 3117 4042 3122
rect 3710 2641 3738 2646
rect 3822 2953 3850 2959
rect 3822 2927 3823 2953
rect 3849 2927 3850 2953
rect 3654 2562 3682 2567
rect 3486 2561 3682 2562
rect 3486 2535 3655 2561
rect 3681 2535 3682 2561
rect 3486 2534 3682 2535
rect 3654 2529 3682 2534
rect 2534 2249 2562 2254
rect 3430 2226 3458 2231
rect 3430 2225 3626 2226
rect 3430 2199 3431 2225
rect 3457 2199 3626 2225
rect 3430 2198 3626 2199
rect 3430 2193 3458 2198
rect 3262 2169 3290 2175
rect 3262 2143 3263 2169
rect 3289 2143 3290 2169
rect 1582 2113 1610 2119
rect 1582 2087 1583 2113
rect 1609 2087 1610 2113
rect 1582 2058 1610 2087
rect 3094 2114 3122 2119
rect 3262 2114 3290 2143
rect 3094 2113 3290 2114
rect 3094 2087 3095 2113
rect 3121 2087 3290 2113
rect 3094 2086 3290 2087
rect 3094 2058 3122 2086
rect 1582 2025 1610 2030
rect 2982 2030 3122 2058
rect 1432 1974 1564 1979
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1432 1941 1564 1946
rect 1246 1807 1247 1833
rect 1273 1807 1274 1833
rect 1246 1801 1274 1807
rect 1022 1721 1106 1722
rect 1022 1695 1023 1721
rect 1049 1695 1106 1721
rect 1022 1694 1106 1695
rect 1470 1722 1498 1727
rect 1022 1689 1050 1694
rect 1470 1675 1498 1694
rect 2258 1582 2390 1587
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2258 1549 2390 1554
rect 2982 1442 3010 2030
rect 3084 1974 3216 1979
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3084 1941 3216 1946
rect 3374 1778 3402 1783
rect 3542 1778 3570 1783
rect 3374 1777 3542 1778
rect 3374 1751 3375 1777
rect 3401 1751 3542 1777
rect 3374 1750 3542 1751
rect 3374 1745 3402 1750
rect 3486 1666 3514 1671
rect 3374 1665 3514 1666
rect 3374 1639 3487 1665
rect 3513 1639 3514 1665
rect 3374 1638 3514 1639
rect 2982 1414 3066 1442
rect 3038 400 3066 1414
rect 3374 400 3402 1638
rect 3486 1633 3514 1638
rect 3542 1106 3570 1750
rect 3598 1777 3626 2198
rect 3598 1751 3599 1777
rect 3625 1751 3626 1777
rect 3598 1745 3626 1751
rect 3822 1721 3850 2927
rect 3934 2562 3962 2567
rect 3934 2515 3962 2534
rect 3910 2366 4042 2371
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 3910 2333 4042 2338
rect 4102 2282 4130 3374
rect 4102 2249 4130 2254
rect 4158 3010 4186 3711
rect 4494 3738 4522 4551
rect 4494 3705 4522 3710
rect 4046 2114 4074 2119
rect 4046 2113 4130 2114
rect 4046 2087 4047 2113
rect 4073 2087 4130 2113
rect 4046 2086 4130 2087
rect 4046 2081 4074 2086
rect 3934 1778 3962 1783
rect 3934 1731 3962 1750
rect 4102 1778 4130 2086
rect 3822 1695 3823 1721
rect 3849 1695 3850 1721
rect 3822 1689 3850 1695
rect 3910 1582 4042 1587
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 3910 1549 4042 1554
rect 4102 1498 4130 1750
rect 4158 1721 4186 2982
rect 4270 3681 4298 3687
rect 4270 3655 4271 3681
rect 4297 3655 4298 3681
rect 4270 2953 4298 3655
rect 4662 3178 4690 5166
rect 4736 5110 4868 5115
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4998 5082 5026 6118
rect 5222 6090 5250 6095
rect 5222 6089 5474 6090
rect 5222 6063 5223 6089
rect 5249 6063 5474 6089
rect 5222 6062 5474 6063
rect 5222 6057 5250 6062
rect 5222 5698 5250 5703
rect 5222 5651 5250 5670
rect 5278 5305 5306 5311
rect 5278 5279 5279 5305
rect 5305 5279 5306 5305
rect 4736 5077 4868 5082
rect 4942 5054 5026 5082
rect 5166 5249 5194 5255
rect 5166 5223 5167 5249
rect 5193 5223 5194 5249
rect 4886 4857 4914 4863
rect 4886 4831 4887 4857
rect 4913 4831 4914 4857
rect 4718 4522 4746 4527
rect 4746 4494 4802 4522
rect 4718 4489 4746 4494
rect 4774 4465 4802 4494
rect 4774 4439 4775 4465
rect 4801 4439 4802 4465
rect 4774 4433 4802 4439
rect 4886 4466 4914 4831
rect 4942 4858 4970 5054
rect 4942 4522 4970 4830
rect 4998 4857 5026 4863
rect 4998 4831 4999 4857
rect 5025 4831 5026 4857
rect 4998 4802 5026 4831
rect 4998 4769 5026 4774
rect 4998 4522 5026 4527
rect 4942 4521 5026 4522
rect 4942 4495 4999 4521
rect 5025 4495 5026 4521
rect 4942 4494 5026 4495
rect 4998 4489 5026 4494
rect 4886 4433 4914 4438
rect 4736 4326 4868 4331
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4736 4293 4868 4298
rect 4886 4242 4914 4247
rect 4886 4073 4914 4214
rect 5166 4242 5194 5223
rect 5278 5250 5306 5279
rect 5278 5217 5306 5222
rect 5446 4633 5474 6062
rect 5562 5502 5694 5507
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5562 5469 5694 5474
rect 5726 5362 5754 7600
rect 5838 6762 5866 6767
rect 5838 6145 5866 6734
rect 6342 6426 6370 6431
rect 5838 6119 5839 6145
rect 5865 6119 5866 6145
rect 5838 6113 5866 6119
rect 6286 6398 6342 6426
rect 6230 6090 6258 6095
rect 6230 5753 6258 6062
rect 6230 5727 6231 5753
rect 6257 5727 6258 5753
rect 6230 5721 6258 5727
rect 5726 5329 5754 5334
rect 6286 5361 6314 6398
rect 6342 6393 6370 6398
rect 7214 6286 7346 6291
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7214 6253 7346 6258
rect 6790 6202 6818 6207
rect 6790 6089 6818 6174
rect 6790 6063 6791 6089
rect 6817 6063 6818 6089
rect 6790 6057 6818 6063
rect 6566 6033 6594 6039
rect 6566 6007 6567 6033
rect 6593 6007 6594 6033
rect 6388 5894 6520 5899
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6388 5861 6520 5866
rect 6286 5335 6287 5361
rect 6313 5335 6314 5361
rect 6286 5329 6314 5335
rect 5614 5249 5642 5255
rect 5782 5250 5810 5255
rect 5614 5223 5615 5249
rect 5641 5223 5642 5249
rect 5614 5194 5642 5223
rect 5614 5161 5642 5166
rect 5726 5222 5782 5250
rect 5562 4718 5694 4723
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5562 4685 5694 4690
rect 5446 4607 5447 4633
rect 5473 4607 5474 4633
rect 5446 4601 5474 4607
rect 5614 4578 5642 4583
rect 5726 4578 5754 5222
rect 5782 5217 5810 5222
rect 6566 5250 6594 6007
rect 6734 6033 6762 6039
rect 6734 6007 6735 6033
rect 6761 6007 6762 6033
rect 6734 5698 6762 6007
rect 6958 5753 6986 5759
rect 6958 5727 6959 5753
rect 6985 5727 6986 5753
rect 6734 5665 6762 5670
rect 6790 5697 6818 5703
rect 6790 5671 6791 5697
rect 6817 5671 6818 5697
rect 6566 5217 6594 5222
rect 6388 5110 6520 5115
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6388 5077 6520 5082
rect 6678 5026 6706 5031
rect 6790 5026 6818 5671
rect 6958 5698 6986 5727
rect 6958 5665 6986 5670
rect 7214 5502 7346 5507
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7214 5469 7346 5474
rect 7014 5305 7042 5311
rect 7014 5279 7015 5305
rect 7041 5279 7042 5305
rect 6846 5194 6874 5199
rect 6874 5166 6930 5194
rect 6846 5161 6874 5166
rect 6790 4998 6874 5026
rect 5838 4969 5866 4975
rect 5838 4943 5839 4969
rect 5865 4943 5866 4969
rect 5838 4634 5866 4943
rect 5838 4601 5866 4606
rect 6286 4913 6314 4919
rect 6286 4887 6287 4913
rect 6313 4887 6314 4913
rect 5614 4577 5754 4578
rect 5614 4551 5615 4577
rect 5641 4551 5754 4577
rect 5614 4550 5754 4551
rect 5614 4545 5642 4550
rect 5894 4522 5922 4527
rect 5166 4209 5194 4214
rect 5222 4466 5250 4471
rect 4998 4186 5026 4191
rect 4998 4139 5026 4158
rect 5222 4130 5250 4438
rect 5894 4242 5922 4494
rect 5894 4209 5922 4214
rect 5390 4130 5418 4135
rect 5222 4102 5390 4130
rect 5390 4083 5418 4102
rect 4886 4047 4887 4073
rect 4913 4047 4914 4073
rect 4886 4041 4914 4047
rect 5562 3934 5694 3939
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5562 3901 5694 3906
rect 5166 3737 5194 3743
rect 5166 3711 5167 3737
rect 5193 3711 5194 3737
rect 4736 3542 4868 3547
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4736 3509 4868 3514
rect 4886 3346 4914 3351
rect 4886 3289 4914 3318
rect 4886 3263 4887 3289
rect 4913 3263 4914 3289
rect 4886 3257 4914 3263
rect 4998 3290 5026 3295
rect 4998 3243 5026 3262
rect 4662 3145 4690 3150
rect 5166 3234 5194 3711
rect 5894 3738 5922 3743
rect 5894 3691 5922 3710
rect 4270 2927 4271 2953
rect 4297 2927 4298 2953
rect 4270 2562 4298 2927
rect 4494 2954 4522 2959
rect 4942 2954 4970 2959
rect 4494 2953 4970 2954
rect 4494 2927 4495 2953
rect 4521 2927 4943 2953
rect 4969 2927 4970 2953
rect 4494 2926 4970 2927
rect 4494 2921 4522 2926
rect 4942 2921 4970 2926
rect 5166 2842 5194 3206
rect 5222 3681 5250 3687
rect 5222 3655 5223 3681
rect 5249 3655 5250 3681
rect 5222 3346 5250 3655
rect 5222 2953 5250 3318
rect 5446 3681 5474 3687
rect 5446 3655 5447 3681
rect 5473 3655 5474 3681
rect 5446 3009 5474 3655
rect 6286 3682 6314 4887
rect 6678 4577 6706 4998
rect 6734 4802 6762 4807
rect 6734 4755 6762 4774
rect 6678 4551 6679 4577
rect 6705 4551 6706 4577
rect 6678 4545 6706 4551
rect 6622 4410 6650 4415
rect 6388 4326 6520 4331
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6388 4293 6520 4298
rect 6342 4185 6370 4191
rect 6342 4159 6343 4185
rect 6369 4159 6370 4185
rect 6342 4074 6370 4159
rect 6342 4041 6370 4046
rect 6622 3793 6650 4382
rect 6846 4186 6874 4998
rect 6846 4153 6874 4158
rect 6790 4129 6818 4135
rect 6790 4103 6791 4129
rect 6817 4103 6818 4129
rect 6790 4074 6818 4103
rect 6790 4046 6874 4074
rect 6790 3850 6818 3855
rect 6622 3767 6623 3793
rect 6649 3767 6650 3793
rect 6622 3761 6650 3767
rect 6734 3822 6790 3850
rect 6286 3649 6314 3654
rect 6678 3738 6706 3743
rect 6388 3542 6520 3547
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6388 3509 6520 3514
rect 6286 3402 6314 3407
rect 6286 3355 6314 3374
rect 5562 3150 5694 3155
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5562 3117 5694 3122
rect 5446 2983 5447 3009
rect 5473 2983 5474 3009
rect 5446 2977 5474 2983
rect 5614 3009 5642 3015
rect 5614 2983 5615 3009
rect 5641 2983 5642 3009
rect 5222 2927 5223 2953
rect 5249 2927 5250 2953
rect 5222 2921 5250 2927
rect 5614 2954 5642 2983
rect 6678 3009 6706 3710
rect 6734 3289 6762 3822
rect 6790 3817 6818 3822
rect 6734 3263 6735 3289
rect 6761 3263 6762 3289
rect 6734 3257 6762 3263
rect 6790 3682 6818 3687
rect 6790 3178 6818 3654
rect 6846 3290 6874 4046
rect 6902 3402 6930 5166
rect 6958 4969 6986 4975
rect 6958 4943 6959 4969
rect 6985 4943 6986 4969
rect 6958 4522 6986 4943
rect 6958 4489 6986 4494
rect 7014 4242 7042 5279
rect 7214 4718 7346 4723
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7214 4685 7346 4690
rect 6958 4214 7042 4242
rect 6958 3850 6986 4214
rect 7014 4130 7042 4135
rect 7014 4083 7042 4102
rect 7214 3934 7346 3939
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7214 3901 7346 3906
rect 6958 3817 6986 3822
rect 6902 3374 6986 3402
rect 6846 3257 6874 3262
rect 6902 3289 6930 3295
rect 6902 3263 6903 3289
rect 6929 3263 6930 3289
rect 6902 3234 6930 3263
rect 6902 3201 6930 3206
rect 6678 2983 6679 3009
rect 6705 2983 6706 3009
rect 6678 2977 6706 2983
rect 6734 3150 6818 3178
rect 5782 2954 5810 2959
rect 5614 2953 5810 2954
rect 5614 2927 5783 2953
rect 5809 2927 5810 2953
rect 5614 2926 5810 2927
rect 5782 2921 5810 2926
rect 5222 2842 5250 2847
rect 5166 2814 5222 2842
rect 5222 2809 5250 2814
rect 6286 2842 6314 2847
rect 4736 2758 4868 2763
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4736 2725 4868 2730
rect 4270 2529 4298 2534
rect 4774 2674 4802 2679
rect 4774 2169 4802 2646
rect 4774 2143 4775 2169
rect 4801 2143 4802 2169
rect 4774 2137 4802 2143
rect 4942 2562 4970 2567
rect 4382 2058 4410 2063
rect 4270 1778 4298 1783
rect 4270 1731 4298 1750
rect 4158 1695 4159 1721
rect 4185 1695 4186 1721
rect 4158 1689 4186 1695
rect 4046 1470 4130 1498
rect 3542 1078 3738 1106
rect 3710 400 3738 1078
rect 4046 400 4074 1470
rect 4382 400 4410 2030
rect 4736 1974 4868 1979
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4736 1941 4868 1946
rect 4718 1834 4746 1839
rect 4718 400 4746 1806
rect 4942 1777 4970 2534
rect 6286 2505 6314 2814
rect 6388 2758 6520 2763
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6388 2725 6520 2730
rect 6566 2730 6594 2735
rect 6566 2618 6594 2702
rect 6454 2590 6594 2618
rect 6454 2561 6482 2590
rect 6454 2535 6455 2561
rect 6481 2535 6482 2561
rect 6454 2529 6482 2535
rect 6286 2479 6287 2505
rect 6313 2479 6314 2505
rect 6286 2473 6314 2479
rect 5562 2366 5694 2371
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5562 2333 5694 2338
rect 6566 2282 6594 2590
rect 6734 2505 6762 3150
rect 6902 2562 6930 2567
rect 6958 2562 6986 3374
rect 7214 3150 7346 3155
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7214 3117 7346 3122
rect 6902 2561 6986 2562
rect 6902 2535 6903 2561
rect 6929 2535 6986 2561
rect 6902 2534 6986 2535
rect 7070 3066 7098 3071
rect 6902 2529 6930 2534
rect 6734 2479 6735 2505
rect 6761 2479 6762 2505
rect 6734 2473 6762 2479
rect 6622 2282 6650 2287
rect 6566 2281 6650 2282
rect 6566 2255 6623 2281
rect 6649 2255 6650 2281
rect 6566 2254 6650 2255
rect 6622 2249 6650 2254
rect 6902 2282 6930 2287
rect 6902 2235 6930 2254
rect 7070 2226 7098 3038
rect 7214 2366 7346 2371
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7214 2333 7346 2338
rect 7070 2225 7154 2226
rect 7070 2199 7071 2225
rect 7097 2199 7154 2225
rect 7070 2198 7154 2199
rect 7070 2193 7098 2198
rect 5278 2058 5306 2063
rect 5278 2011 5306 2030
rect 6388 1974 6520 1979
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6388 1941 6520 1946
rect 5334 1834 5362 1839
rect 5334 1787 5362 1806
rect 7126 1833 7154 2198
rect 7126 1807 7127 1833
rect 7153 1807 7154 1833
rect 7126 1801 7154 1807
rect 4942 1751 4943 1777
rect 4969 1751 4970 1777
rect 4942 1745 4970 1751
rect 5562 1582 5694 1587
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5562 1549 5694 1554
rect 7214 1582 7346 1587
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7214 1549 7346 1554
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
<< via2 >>
rect 3598 7070 3626 7098
rect 2258 6285 2286 6286
rect 2258 6259 2259 6285
rect 2259 6259 2285 6285
rect 2285 6259 2286 6285
rect 2258 6258 2286 6259
rect 2310 6285 2338 6286
rect 2310 6259 2311 6285
rect 2311 6259 2337 6285
rect 2337 6259 2338 6285
rect 2310 6258 2338 6259
rect 2362 6285 2390 6286
rect 2362 6259 2363 6285
rect 2363 6259 2389 6285
rect 2389 6259 2390 6285
rect 2362 6258 2390 6259
rect 3430 6145 3458 6146
rect 3430 6119 3431 6145
rect 3431 6119 3457 6145
rect 3457 6119 3458 6145
rect 3430 6118 3458 6119
rect 3910 6285 3938 6286
rect 3910 6259 3911 6285
rect 3911 6259 3937 6285
rect 3937 6259 3938 6285
rect 3910 6258 3938 6259
rect 3962 6285 3990 6286
rect 3962 6259 3963 6285
rect 3963 6259 3989 6285
rect 3989 6259 3990 6285
rect 3962 6258 3990 6259
rect 4014 6285 4042 6286
rect 4014 6259 4015 6285
rect 4015 6259 4041 6285
rect 4041 6259 4042 6285
rect 4014 6258 4042 6259
rect 4046 6201 4074 6202
rect 4046 6175 4047 6201
rect 4047 6175 4073 6201
rect 4073 6175 4074 6201
rect 4046 6174 4074 6175
rect 3206 5950 3234 5978
rect 1432 5893 1460 5894
rect 1432 5867 1433 5893
rect 1433 5867 1459 5893
rect 1459 5867 1460 5893
rect 1432 5866 1460 5867
rect 1484 5893 1512 5894
rect 1484 5867 1485 5893
rect 1485 5867 1511 5893
rect 1511 5867 1512 5893
rect 1484 5866 1512 5867
rect 1536 5893 1564 5894
rect 1536 5867 1537 5893
rect 1537 5867 1563 5893
rect 1563 5867 1564 5893
rect 1536 5866 1564 5867
rect 3084 5893 3112 5894
rect 3084 5867 3085 5893
rect 3085 5867 3111 5893
rect 3111 5867 3112 5893
rect 3084 5866 3112 5867
rect 3136 5893 3164 5894
rect 3136 5867 3137 5893
rect 3137 5867 3163 5893
rect 3163 5867 3164 5893
rect 3136 5866 3164 5867
rect 3188 5893 3216 5894
rect 3188 5867 3189 5893
rect 3189 5867 3215 5893
rect 3215 5867 3216 5893
rect 3188 5866 3216 5867
rect 2258 5501 2286 5502
rect 2258 5475 2259 5501
rect 2259 5475 2285 5501
rect 2285 5475 2286 5501
rect 2258 5474 2286 5475
rect 2310 5501 2338 5502
rect 2310 5475 2311 5501
rect 2311 5475 2337 5501
rect 2337 5475 2338 5501
rect 2310 5474 2338 5475
rect 2362 5501 2390 5502
rect 2362 5475 2363 5501
rect 2363 5475 2389 5501
rect 2389 5475 2390 5501
rect 2362 5474 2390 5475
rect 3766 6062 3794 6090
rect 3934 5950 3962 5978
rect 3910 5501 3938 5502
rect 3910 5475 3911 5501
rect 3911 5475 3937 5501
rect 3937 5475 3938 5501
rect 3910 5474 3938 5475
rect 3962 5501 3990 5502
rect 3962 5475 3963 5501
rect 3963 5475 3989 5501
rect 3989 5475 3990 5501
rect 3962 5474 3990 5475
rect 4014 5501 4042 5502
rect 4014 5475 4015 5501
rect 4015 5475 4041 5501
rect 4041 5475 4042 5501
rect 4014 5474 4042 5475
rect 4214 5417 4242 5418
rect 4214 5391 4215 5417
rect 4215 5391 4241 5417
rect 4241 5391 4242 5417
rect 4214 5390 4242 5391
rect 3990 5361 4018 5362
rect 3990 5335 3991 5361
rect 3991 5335 4017 5361
rect 4017 5335 4018 5361
rect 3990 5334 4018 5335
rect 3710 5222 3738 5250
rect 4046 5222 4074 5250
rect 1432 5109 1460 5110
rect 1432 5083 1433 5109
rect 1433 5083 1459 5109
rect 1459 5083 1460 5109
rect 1432 5082 1460 5083
rect 1484 5109 1512 5110
rect 1484 5083 1485 5109
rect 1485 5083 1511 5109
rect 1511 5083 1512 5109
rect 1484 5082 1512 5083
rect 1536 5109 1564 5110
rect 1536 5083 1537 5109
rect 1537 5083 1563 5109
rect 1563 5083 1564 5109
rect 1536 5082 1564 5083
rect 3084 5109 3112 5110
rect 3084 5083 3085 5109
rect 3085 5083 3111 5109
rect 3111 5083 3112 5109
rect 3084 5082 3112 5083
rect 3136 5109 3164 5110
rect 3136 5083 3137 5109
rect 3137 5083 3163 5109
rect 3163 5083 3164 5109
rect 3136 5082 3164 5083
rect 3188 5109 3216 5110
rect 3188 5083 3189 5109
rect 3189 5083 3215 5109
rect 3215 5083 3216 5109
rect 3188 5082 3216 5083
rect 854 4718 882 4746
rect 854 4382 882 4410
rect 854 4073 882 4074
rect 854 4047 855 4073
rect 855 4047 881 4073
rect 881 4047 882 4073
rect 854 4046 882 4047
rect 910 3654 938 3682
rect 910 3374 938 3402
rect 854 3038 882 3066
rect 1246 4718 1274 4746
rect 2258 4717 2286 4718
rect 2258 4691 2259 4717
rect 2259 4691 2285 4717
rect 2285 4691 2286 4717
rect 2258 4690 2286 4691
rect 2310 4717 2338 4718
rect 2310 4691 2311 4717
rect 2311 4691 2337 4717
rect 2337 4691 2338 4717
rect 2310 4690 2338 4691
rect 2362 4717 2390 4718
rect 2362 4691 2363 4717
rect 2363 4691 2389 4717
rect 2389 4691 2390 4717
rect 2362 4690 2390 4691
rect 3910 4717 3938 4718
rect 3910 4691 3911 4717
rect 3911 4691 3937 4717
rect 3937 4691 3938 4717
rect 3910 4690 3938 4691
rect 3962 4717 3990 4718
rect 3962 4691 3963 4717
rect 3963 4691 3989 4717
rect 3989 4691 3990 4717
rect 3962 4690 3990 4691
rect 4014 4717 4042 4718
rect 4014 4691 4015 4717
rect 4015 4691 4041 4717
rect 4041 4691 4042 4717
rect 4014 4690 4042 4691
rect 1246 4382 1274 4410
rect 1432 4325 1460 4326
rect 1432 4299 1433 4325
rect 1433 4299 1459 4325
rect 1459 4299 1460 4325
rect 1432 4298 1460 4299
rect 1484 4325 1512 4326
rect 1484 4299 1485 4325
rect 1485 4299 1511 4325
rect 1511 4299 1512 4325
rect 1484 4298 1512 4299
rect 1536 4325 1564 4326
rect 1536 4299 1537 4325
rect 1537 4299 1563 4325
rect 1563 4299 1564 4325
rect 1536 4298 1564 4299
rect 3084 4325 3112 4326
rect 3084 4299 3085 4325
rect 3085 4299 3111 4325
rect 3111 4299 3112 4325
rect 3084 4298 3112 4299
rect 3136 4325 3164 4326
rect 3136 4299 3137 4325
rect 3137 4299 3163 4325
rect 3163 4299 3164 4325
rect 3136 4298 3164 4299
rect 3188 4325 3216 4326
rect 3188 4299 3189 4325
rect 3189 4299 3215 4325
rect 3215 4299 3216 4325
rect 3188 4298 3216 4299
rect 1078 3766 1106 3794
rect 1806 4073 1834 4074
rect 1806 4047 1807 4073
rect 1807 4047 1833 4073
rect 1833 4047 1834 4073
rect 1806 4046 1834 4047
rect 4382 6145 4410 6146
rect 4382 6119 4383 6145
rect 4383 6119 4409 6145
rect 4409 6119 4410 6145
rect 4382 6118 4410 6119
rect 5562 6285 5590 6286
rect 5562 6259 5563 6285
rect 5563 6259 5589 6285
rect 5589 6259 5590 6285
rect 5562 6258 5590 6259
rect 5614 6285 5642 6286
rect 5614 6259 5615 6285
rect 5615 6259 5641 6285
rect 5641 6259 5642 6285
rect 5614 6258 5642 6259
rect 5666 6285 5694 6286
rect 5666 6259 5667 6285
rect 5667 6259 5693 6285
rect 5693 6259 5694 6285
rect 5666 6258 5694 6259
rect 4718 6089 4746 6090
rect 4718 6063 4719 6089
rect 4719 6063 4745 6089
rect 4745 6063 4746 6089
rect 4718 6062 4746 6063
rect 4736 5893 4764 5894
rect 4736 5867 4737 5893
rect 4737 5867 4763 5893
rect 4763 5867 4764 5893
rect 4736 5866 4764 5867
rect 4788 5893 4816 5894
rect 4788 5867 4789 5893
rect 4789 5867 4815 5893
rect 4815 5867 4816 5893
rect 4788 5866 4816 5867
rect 4840 5893 4868 5894
rect 4840 5867 4841 5893
rect 4841 5867 4867 5893
rect 4867 5867 4868 5893
rect 4840 5866 4868 5867
rect 4326 5697 4354 5698
rect 4326 5671 4327 5697
rect 4327 5671 4353 5697
rect 4353 5671 4354 5697
rect 4326 5670 4354 5671
rect 4774 5670 4802 5698
rect 4494 5390 4522 5418
rect 4214 4857 4242 4858
rect 4214 4831 4215 4857
rect 4215 4831 4241 4857
rect 4241 4831 4242 4857
rect 4214 4830 4242 4831
rect 4886 5670 4914 5698
rect 4942 5361 4970 5362
rect 4942 5335 4943 5361
rect 4943 5335 4969 5361
rect 4969 5335 4970 5361
rect 4942 5334 4970 5335
rect 4382 4521 4410 4522
rect 4382 4495 4383 4521
rect 4383 4495 4409 4521
rect 4409 4495 4410 4521
rect 4382 4494 4410 4495
rect 2258 3933 2286 3934
rect 2258 3907 2259 3933
rect 2259 3907 2285 3933
rect 2285 3907 2286 3933
rect 2258 3906 2286 3907
rect 2310 3933 2338 3934
rect 2310 3907 2311 3933
rect 2311 3907 2337 3933
rect 2337 3907 2338 3933
rect 2310 3906 2338 3907
rect 2362 3933 2390 3934
rect 2362 3907 2363 3933
rect 2363 3907 2389 3933
rect 2389 3907 2390 3933
rect 2362 3906 2390 3907
rect 3910 3933 3938 3934
rect 3910 3907 3911 3933
rect 3911 3907 3937 3933
rect 3937 3907 3938 3933
rect 3910 3906 3938 3907
rect 3962 3933 3990 3934
rect 3962 3907 3963 3933
rect 3963 3907 3989 3933
rect 3989 3907 3990 3933
rect 3962 3906 3990 3907
rect 4014 3933 4042 3934
rect 4014 3907 4015 3933
rect 4015 3907 4041 3933
rect 4041 3907 4042 3933
rect 4014 3906 4042 3907
rect 1302 3710 1330 3738
rect 1750 3681 1778 3682
rect 1750 3655 1751 3681
rect 1751 3655 1777 3681
rect 1777 3655 1778 3681
rect 1750 3654 1778 3655
rect 1078 3318 1106 3346
rect 1432 3541 1460 3542
rect 1432 3515 1433 3541
rect 1433 3515 1459 3541
rect 1459 3515 1460 3541
rect 1432 3514 1460 3515
rect 1484 3541 1512 3542
rect 1484 3515 1485 3541
rect 1485 3515 1511 3541
rect 1511 3515 1512 3541
rect 1484 3514 1512 3515
rect 1536 3541 1564 3542
rect 1536 3515 1537 3541
rect 1537 3515 1563 3541
rect 1563 3515 1564 3541
rect 1536 3514 1564 3515
rect 1022 2926 1050 2954
rect 854 2590 882 2618
rect 966 2646 994 2674
rect 854 2366 882 2394
rect 854 1721 882 1722
rect 854 1695 855 1721
rect 855 1695 881 1721
rect 881 1695 882 1721
rect 854 1694 882 1695
rect 2198 3318 2226 3346
rect 1190 2702 1218 2730
rect 1190 2561 1218 2562
rect 1190 2535 1191 2561
rect 1191 2535 1217 2561
rect 1217 2535 1218 2561
rect 1190 2534 1218 2535
rect 2258 3149 2286 3150
rect 2258 3123 2259 3149
rect 2259 3123 2285 3149
rect 2285 3123 2286 3149
rect 2258 3122 2286 3123
rect 2310 3149 2338 3150
rect 2310 3123 2311 3149
rect 2311 3123 2337 3149
rect 2337 3123 2338 3149
rect 2310 3122 2338 3123
rect 2362 3149 2390 3150
rect 2362 3123 2363 3149
rect 2363 3123 2389 3149
rect 2389 3123 2390 3149
rect 2362 3122 2390 3123
rect 2366 2953 2394 2954
rect 2366 2927 2367 2953
rect 2367 2927 2393 2953
rect 2393 2927 2394 2953
rect 2366 2926 2394 2927
rect 1432 2757 1460 2758
rect 1432 2731 1433 2757
rect 1433 2731 1459 2757
rect 1459 2731 1460 2757
rect 1432 2730 1460 2731
rect 1484 2757 1512 2758
rect 1484 2731 1485 2757
rect 1485 2731 1511 2757
rect 1511 2731 1512 2757
rect 1484 2730 1512 2731
rect 1536 2757 1564 2758
rect 1536 2731 1537 2757
rect 1537 2731 1563 2757
rect 1563 2731 1564 2757
rect 1536 2730 1564 2731
rect 1806 2617 1834 2618
rect 1806 2591 1807 2617
rect 1807 2591 1833 2617
rect 1833 2591 1834 2617
rect 1806 2590 1834 2591
rect 1582 2561 1610 2562
rect 1582 2535 1583 2561
rect 1583 2535 1609 2561
rect 1609 2535 1610 2561
rect 1582 2534 1610 2535
rect 1246 2366 1274 2394
rect 1190 2030 1218 2058
rect 2258 2365 2286 2366
rect 2258 2339 2259 2365
rect 2259 2339 2285 2365
rect 2285 2339 2286 2365
rect 2258 2338 2286 2339
rect 2310 2365 2338 2366
rect 2310 2339 2311 2365
rect 2311 2339 2337 2365
rect 2337 2339 2338 2365
rect 2310 2338 2338 2339
rect 2362 2365 2390 2366
rect 2362 2339 2363 2365
rect 2363 2339 2389 2365
rect 2389 2339 2390 2365
rect 2362 2338 2390 2339
rect 1358 2281 1386 2282
rect 1358 2255 1359 2281
rect 1359 2255 1385 2281
rect 1385 2255 1386 2281
rect 1358 2254 1386 2255
rect 2870 3766 2898 3794
rect 3084 3541 3112 3542
rect 3084 3515 3085 3541
rect 3085 3515 3111 3541
rect 3111 3515 3112 3541
rect 3084 3514 3112 3515
rect 3136 3541 3164 3542
rect 3136 3515 3137 3541
rect 3137 3515 3163 3541
rect 3163 3515 3164 3541
rect 3136 3514 3164 3515
rect 3188 3541 3216 3542
rect 3188 3515 3189 3541
rect 3189 3515 3215 3541
rect 3215 3515 3216 3541
rect 3188 3514 3216 3515
rect 3084 2757 3112 2758
rect 3084 2731 3085 2757
rect 3085 2731 3111 2757
rect 3111 2731 3112 2757
rect 3084 2730 3112 2731
rect 3136 2757 3164 2758
rect 3136 2731 3137 2757
rect 3137 2731 3163 2757
rect 3163 2731 3164 2757
rect 3136 2730 3164 2731
rect 3188 2757 3216 2758
rect 3188 2731 3189 2757
rect 3189 2731 3215 2757
rect 3215 2731 3216 2757
rect 3188 2730 3216 2731
rect 2982 2646 3010 2674
rect 3654 3009 3682 3010
rect 3654 2983 3655 3009
rect 3655 2983 3681 3009
rect 3681 2983 3682 3009
rect 3654 2982 3682 2983
rect 4046 3206 4074 3234
rect 3910 3149 3938 3150
rect 3910 3123 3911 3149
rect 3911 3123 3937 3149
rect 3937 3123 3938 3149
rect 3910 3122 3938 3123
rect 3962 3149 3990 3150
rect 3962 3123 3963 3149
rect 3963 3123 3989 3149
rect 3989 3123 3990 3149
rect 3962 3122 3990 3123
rect 4014 3149 4042 3150
rect 4014 3123 4015 3149
rect 4015 3123 4041 3149
rect 4041 3123 4042 3149
rect 4014 3122 4042 3123
rect 3710 2646 3738 2674
rect 2534 2254 2562 2282
rect 1582 2030 1610 2058
rect 1432 1973 1460 1974
rect 1432 1947 1433 1973
rect 1433 1947 1459 1973
rect 1459 1947 1460 1973
rect 1432 1946 1460 1947
rect 1484 1973 1512 1974
rect 1484 1947 1485 1973
rect 1485 1947 1511 1973
rect 1511 1947 1512 1973
rect 1484 1946 1512 1947
rect 1536 1973 1564 1974
rect 1536 1947 1537 1973
rect 1537 1947 1563 1973
rect 1563 1947 1564 1973
rect 1536 1946 1564 1947
rect 1470 1721 1498 1722
rect 1470 1695 1471 1721
rect 1471 1695 1497 1721
rect 1497 1695 1498 1721
rect 1470 1694 1498 1695
rect 2258 1581 2286 1582
rect 2258 1555 2259 1581
rect 2259 1555 2285 1581
rect 2285 1555 2286 1581
rect 2258 1554 2286 1555
rect 2310 1581 2338 1582
rect 2310 1555 2311 1581
rect 2311 1555 2337 1581
rect 2337 1555 2338 1581
rect 2310 1554 2338 1555
rect 2362 1581 2390 1582
rect 2362 1555 2363 1581
rect 2363 1555 2389 1581
rect 2389 1555 2390 1581
rect 2362 1554 2390 1555
rect 3084 1973 3112 1974
rect 3084 1947 3085 1973
rect 3085 1947 3111 1973
rect 3111 1947 3112 1973
rect 3084 1946 3112 1947
rect 3136 1973 3164 1974
rect 3136 1947 3137 1973
rect 3137 1947 3163 1973
rect 3163 1947 3164 1973
rect 3136 1946 3164 1947
rect 3188 1973 3216 1974
rect 3188 1947 3189 1973
rect 3189 1947 3215 1973
rect 3215 1947 3216 1973
rect 3188 1946 3216 1947
rect 3542 1750 3570 1778
rect 3934 2561 3962 2562
rect 3934 2535 3935 2561
rect 3935 2535 3961 2561
rect 3961 2535 3962 2561
rect 3934 2534 3962 2535
rect 3910 2365 3938 2366
rect 3910 2339 3911 2365
rect 3911 2339 3937 2365
rect 3937 2339 3938 2365
rect 3910 2338 3938 2339
rect 3962 2365 3990 2366
rect 3962 2339 3963 2365
rect 3963 2339 3989 2365
rect 3989 2339 3990 2365
rect 3962 2338 3990 2339
rect 4014 2365 4042 2366
rect 4014 2339 4015 2365
rect 4015 2339 4041 2365
rect 4041 2339 4042 2365
rect 4014 2338 4042 2339
rect 4102 2254 4130 2282
rect 4494 3710 4522 3738
rect 4158 2982 4186 3010
rect 3934 1777 3962 1778
rect 3934 1751 3935 1777
rect 3935 1751 3961 1777
rect 3961 1751 3962 1777
rect 3934 1750 3962 1751
rect 4102 1750 4130 1778
rect 3910 1581 3938 1582
rect 3910 1555 3911 1581
rect 3911 1555 3937 1581
rect 3937 1555 3938 1581
rect 3910 1554 3938 1555
rect 3962 1581 3990 1582
rect 3962 1555 3963 1581
rect 3963 1555 3989 1581
rect 3989 1555 3990 1581
rect 3962 1554 3990 1555
rect 4014 1581 4042 1582
rect 4014 1555 4015 1581
rect 4015 1555 4041 1581
rect 4041 1555 4042 1581
rect 4014 1554 4042 1555
rect 4736 5109 4764 5110
rect 4736 5083 4737 5109
rect 4737 5083 4763 5109
rect 4763 5083 4764 5109
rect 4736 5082 4764 5083
rect 4788 5109 4816 5110
rect 4788 5083 4789 5109
rect 4789 5083 4815 5109
rect 4815 5083 4816 5109
rect 4788 5082 4816 5083
rect 4840 5109 4868 5110
rect 4840 5083 4841 5109
rect 4841 5083 4867 5109
rect 4867 5083 4868 5109
rect 4840 5082 4868 5083
rect 5222 5697 5250 5698
rect 5222 5671 5223 5697
rect 5223 5671 5249 5697
rect 5249 5671 5250 5697
rect 5222 5670 5250 5671
rect 4718 4494 4746 4522
rect 4942 4830 4970 4858
rect 4998 4774 5026 4802
rect 4886 4438 4914 4466
rect 4736 4325 4764 4326
rect 4736 4299 4737 4325
rect 4737 4299 4763 4325
rect 4763 4299 4764 4325
rect 4736 4298 4764 4299
rect 4788 4325 4816 4326
rect 4788 4299 4789 4325
rect 4789 4299 4815 4325
rect 4815 4299 4816 4325
rect 4788 4298 4816 4299
rect 4840 4325 4868 4326
rect 4840 4299 4841 4325
rect 4841 4299 4867 4325
rect 4867 4299 4868 4325
rect 4840 4298 4868 4299
rect 4886 4214 4914 4242
rect 5278 5222 5306 5250
rect 5562 5501 5590 5502
rect 5562 5475 5563 5501
rect 5563 5475 5589 5501
rect 5589 5475 5590 5501
rect 5562 5474 5590 5475
rect 5614 5501 5642 5502
rect 5614 5475 5615 5501
rect 5615 5475 5641 5501
rect 5641 5475 5642 5501
rect 5614 5474 5642 5475
rect 5666 5501 5694 5502
rect 5666 5475 5667 5501
rect 5667 5475 5693 5501
rect 5693 5475 5694 5501
rect 5666 5474 5694 5475
rect 5838 6734 5866 6762
rect 6342 6398 6370 6426
rect 6230 6062 6258 6090
rect 5726 5334 5754 5362
rect 7214 6285 7242 6286
rect 7214 6259 7215 6285
rect 7215 6259 7241 6285
rect 7241 6259 7242 6285
rect 7214 6258 7242 6259
rect 7266 6285 7294 6286
rect 7266 6259 7267 6285
rect 7267 6259 7293 6285
rect 7293 6259 7294 6285
rect 7266 6258 7294 6259
rect 7318 6285 7346 6286
rect 7318 6259 7319 6285
rect 7319 6259 7345 6285
rect 7345 6259 7346 6285
rect 7318 6258 7346 6259
rect 6790 6174 6818 6202
rect 6388 5893 6416 5894
rect 6388 5867 6389 5893
rect 6389 5867 6415 5893
rect 6415 5867 6416 5893
rect 6388 5866 6416 5867
rect 6440 5893 6468 5894
rect 6440 5867 6441 5893
rect 6441 5867 6467 5893
rect 6467 5867 6468 5893
rect 6440 5866 6468 5867
rect 6492 5893 6520 5894
rect 6492 5867 6493 5893
rect 6493 5867 6519 5893
rect 6519 5867 6520 5893
rect 6492 5866 6520 5867
rect 5614 5166 5642 5194
rect 5782 5222 5810 5250
rect 5562 4717 5590 4718
rect 5562 4691 5563 4717
rect 5563 4691 5589 4717
rect 5589 4691 5590 4717
rect 5562 4690 5590 4691
rect 5614 4717 5642 4718
rect 5614 4691 5615 4717
rect 5615 4691 5641 4717
rect 5641 4691 5642 4717
rect 5614 4690 5642 4691
rect 5666 4717 5694 4718
rect 5666 4691 5667 4717
rect 5667 4691 5693 4717
rect 5693 4691 5694 4717
rect 5666 4690 5694 4691
rect 6734 5670 6762 5698
rect 6566 5222 6594 5250
rect 6388 5109 6416 5110
rect 6388 5083 6389 5109
rect 6389 5083 6415 5109
rect 6415 5083 6416 5109
rect 6388 5082 6416 5083
rect 6440 5109 6468 5110
rect 6440 5083 6441 5109
rect 6441 5083 6467 5109
rect 6467 5083 6468 5109
rect 6440 5082 6468 5083
rect 6492 5109 6520 5110
rect 6492 5083 6493 5109
rect 6493 5083 6519 5109
rect 6519 5083 6520 5109
rect 6492 5082 6520 5083
rect 6678 4998 6706 5026
rect 6958 5670 6986 5698
rect 7214 5501 7242 5502
rect 7214 5475 7215 5501
rect 7215 5475 7241 5501
rect 7241 5475 7242 5501
rect 7214 5474 7242 5475
rect 7266 5501 7294 5502
rect 7266 5475 7267 5501
rect 7267 5475 7293 5501
rect 7293 5475 7294 5501
rect 7266 5474 7294 5475
rect 7318 5501 7346 5502
rect 7318 5475 7319 5501
rect 7319 5475 7345 5501
rect 7345 5475 7346 5501
rect 7318 5474 7346 5475
rect 6846 5166 6874 5194
rect 5838 4606 5866 4634
rect 5894 4521 5922 4522
rect 5894 4495 5895 4521
rect 5895 4495 5921 4521
rect 5921 4495 5922 4521
rect 5894 4494 5922 4495
rect 5166 4214 5194 4242
rect 5222 4465 5250 4466
rect 5222 4439 5223 4465
rect 5223 4439 5249 4465
rect 5249 4439 5250 4465
rect 5222 4438 5250 4439
rect 4998 4185 5026 4186
rect 4998 4159 4999 4185
rect 4999 4159 5025 4185
rect 5025 4159 5026 4185
rect 4998 4158 5026 4159
rect 5894 4214 5922 4242
rect 5390 4129 5418 4130
rect 5390 4103 5391 4129
rect 5391 4103 5417 4129
rect 5417 4103 5418 4129
rect 5390 4102 5418 4103
rect 5562 3933 5590 3934
rect 5562 3907 5563 3933
rect 5563 3907 5589 3933
rect 5589 3907 5590 3933
rect 5562 3906 5590 3907
rect 5614 3933 5642 3934
rect 5614 3907 5615 3933
rect 5615 3907 5641 3933
rect 5641 3907 5642 3933
rect 5614 3906 5642 3907
rect 5666 3933 5694 3934
rect 5666 3907 5667 3933
rect 5667 3907 5693 3933
rect 5693 3907 5694 3933
rect 5666 3906 5694 3907
rect 4736 3541 4764 3542
rect 4736 3515 4737 3541
rect 4737 3515 4763 3541
rect 4763 3515 4764 3541
rect 4736 3514 4764 3515
rect 4788 3541 4816 3542
rect 4788 3515 4789 3541
rect 4789 3515 4815 3541
rect 4815 3515 4816 3541
rect 4788 3514 4816 3515
rect 4840 3541 4868 3542
rect 4840 3515 4841 3541
rect 4841 3515 4867 3541
rect 4867 3515 4868 3541
rect 4840 3514 4868 3515
rect 4886 3318 4914 3346
rect 4998 3289 5026 3290
rect 4998 3263 4999 3289
rect 4999 3263 5025 3289
rect 5025 3263 5026 3289
rect 4998 3262 5026 3263
rect 4662 3150 4690 3178
rect 5894 3737 5922 3738
rect 5894 3711 5895 3737
rect 5895 3711 5921 3737
rect 5921 3711 5922 3737
rect 5894 3710 5922 3711
rect 5166 3206 5194 3234
rect 5222 3345 5250 3346
rect 5222 3319 5223 3345
rect 5223 3319 5249 3345
rect 5249 3319 5250 3345
rect 5222 3318 5250 3319
rect 6734 4801 6762 4802
rect 6734 4775 6735 4801
rect 6735 4775 6761 4801
rect 6761 4775 6762 4801
rect 6734 4774 6762 4775
rect 6622 4382 6650 4410
rect 6388 4325 6416 4326
rect 6388 4299 6389 4325
rect 6389 4299 6415 4325
rect 6415 4299 6416 4325
rect 6388 4298 6416 4299
rect 6440 4325 6468 4326
rect 6440 4299 6441 4325
rect 6441 4299 6467 4325
rect 6467 4299 6468 4325
rect 6440 4298 6468 4299
rect 6492 4325 6520 4326
rect 6492 4299 6493 4325
rect 6493 4299 6519 4325
rect 6519 4299 6520 4325
rect 6492 4298 6520 4299
rect 6342 4046 6370 4074
rect 6846 4158 6874 4186
rect 6790 3822 6818 3850
rect 6286 3654 6314 3682
rect 6678 3710 6706 3738
rect 6388 3541 6416 3542
rect 6388 3515 6389 3541
rect 6389 3515 6415 3541
rect 6415 3515 6416 3541
rect 6388 3514 6416 3515
rect 6440 3541 6468 3542
rect 6440 3515 6441 3541
rect 6441 3515 6467 3541
rect 6467 3515 6468 3541
rect 6440 3514 6468 3515
rect 6492 3541 6520 3542
rect 6492 3515 6493 3541
rect 6493 3515 6519 3541
rect 6519 3515 6520 3541
rect 6492 3514 6520 3515
rect 6286 3401 6314 3402
rect 6286 3375 6287 3401
rect 6287 3375 6313 3401
rect 6313 3375 6314 3401
rect 6286 3374 6314 3375
rect 5562 3149 5590 3150
rect 5562 3123 5563 3149
rect 5563 3123 5589 3149
rect 5589 3123 5590 3149
rect 5562 3122 5590 3123
rect 5614 3149 5642 3150
rect 5614 3123 5615 3149
rect 5615 3123 5641 3149
rect 5641 3123 5642 3149
rect 5614 3122 5642 3123
rect 5666 3149 5694 3150
rect 5666 3123 5667 3149
rect 5667 3123 5693 3149
rect 5693 3123 5694 3149
rect 5666 3122 5694 3123
rect 6790 3654 6818 3682
rect 6958 4494 6986 4522
rect 7214 4717 7242 4718
rect 7214 4691 7215 4717
rect 7215 4691 7241 4717
rect 7241 4691 7242 4717
rect 7214 4690 7242 4691
rect 7266 4717 7294 4718
rect 7266 4691 7267 4717
rect 7267 4691 7293 4717
rect 7293 4691 7294 4717
rect 7266 4690 7294 4691
rect 7318 4717 7346 4718
rect 7318 4691 7319 4717
rect 7319 4691 7345 4717
rect 7345 4691 7346 4717
rect 7318 4690 7346 4691
rect 7014 4129 7042 4130
rect 7014 4103 7015 4129
rect 7015 4103 7041 4129
rect 7041 4103 7042 4129
rect 7014 4102 7042 4103
rect 7214 3933 7242 3934
rect 7214 3907 7215 3933
rect 7215 3907 7241 3933
rect 7241 3907 7242 3933
rect 7214 3906 7242 3907
rect 7266 3933 7294 3934
rect 7266 3907 7267 3933
rect 7267 3907 7293 3933
rect 7293 3907 7294 3933
rect 7266 3906 7294 3907
rect 7318 3933 7346 3934
rect 7318 3907 7319 3933
rect 7319 3907 7345 3933
rect 7345 3907 7346 3933
rect 7318 3906 7346 3907
rect 6958 3822 6986 3850
rect 6846 3262 6874 3290
rect 6902 3206 6930 3234
rect 5222 2814 5250 2842
rect 6286 2814 6314 2842
rect 4736 2757 4764 2758
rect 4736 2731 4737 2757
rect 4737 2731 4763 2757
rect 4763 2731 4764 2757
rect 4736 2730 4764 2731
rect 4788 2757 4816 2758
rect 4788 2731 4789 2757
rect 4789 2731 4815 2757
rect 4815 2731 4816 2757
rect 4788 2730 4816 2731
rect 4840 2757 4868 2758
rect 4840 2731 4841 2757
rect 4841 2731 4867 2757
rect 4867 2731 4868 2757
rect 4840 2730 4868 2731
rect 4270 2534 4298 2562
rect 4774 2646 4802 2674
rect 4942 2534 4970 2562
rect 4382 2030 4410 2058
rect 4270 1777 4298 1778
rect 4270 1751 4271 1777
rect 4271 1751 4297 1777
rect 4297 1751 4298 1777
rect 4270 1750 4298 1751
rect 4736 1973 4764 1974
rect 4736 1947 4737 1973
rect 4737 1947 4763 1973
rect 4763 1947 4764 1973
rect 4736 1946 4764 1947
rect 4788 1973 4816 1974
rect 4788 1947 4789 1973
rect 4789 1947 4815 1973
rect 4815 1947 4816 1973
rect 4788 1946 4816 1947
rect 4840 1973 4868 1974
rect 4840 1947 4841 1973
rect 4841 1947 4867 1973
rect 4867 1947 4868 1973
rect 4840 1946 4868 1947
rect 4718 1806 4746 1834
rect 6388 2757 6416 2758
rect 6388 2731 6389 2757
rect 6389 2731 6415 2757
rect 6415 2731 6416 2757
rect 6388 2730 6416 2731
rect 6440 2757 6468 2758
rect 6440 2731 6441 2757
rect 6441 2731 6467 2757
rect 6467 2731 6468 2757
rect 6440 2730 6468 2731
rect 6492 2757 6520 2758
rect 6492 2731 6493 2757
rect 6493 2731 6519 2757
rect 6519 2731 6520 2757
rect 6492 2730 6520 2731
rect 6566 2702 6594 2730
rect 5562 2365 5590 2366
rect 5562 2339 5563 2365
rect 5563 2339 5589 2365
rect 5589 2339 5590 2365
rect 5562 2338 5590 2339
rect 5614 2365 5642 2366
rect 5614 2339 5615 2365
rect 5615 2339 5641 2365
rect 5641 2339 5642 2365
rect 5614 2338 5642 2339
rect 5666 2365 5694 2366
rect 5666 2339 5667 2365
rect 5667 2339 5693 2365
rect 5693 2339 5694 2365
rect 5666 2338 5694 2339
rect 7214 3149 7242 3150
rect 7214 3123 7215 3149
rect 7215 3123 7241 3149
rect 7241 3123 7242 3149
rect 7214 3122 7242 3123
rect 7266 3149 7294 3150
rect 7266 3123 7267 3149
rect 7267 3123 7293 3149
rect 7293 3123 7294 3149
rect 7266 3122 7294 3123
rect 7318 3149 7346 3150
rect 7318 3123 7319 3149
rect 7319 3123 7345 3149
rect 7345 3123 7346 3149
rect 7318 3122 7346 3123
rect 7070 3038 7098 3066
rect 6902 2281 6930 2282
rect 6902 2255 6903 2281
rect 6903 2255 6929 2281
rect 6929 2255 6930 2281
rect 6902 2254 6930 2255
rect 7214 2365 7242 2366
rect 7214 2339 7215 2365
rect 7215 2339 7241 2365
rect 7241 2339 7242 2365
rect 7214 2338 7242 2339
rect 7266 2365 7294 2366
rect 7266 2339 7267 2365
rect 7267 2339 7293 2365
rect 7293 2339 7294 2365
rect 7266 2338 7294 2339
rect 7318 2365 7346 2366
rect 7318 2339 7319 2365
rect 7319 2339 7345 2365
rect 7345 2339 7346 2365
rect 7318 2338 7346 2339
rect 5278 2057 5306 2058
rect 5278 2031 5279 2057
rect 5279 2031 5305 2057
rect 5305 2031 5306 2057
rect 5278 2030 5306 2031
rect 6388 1973 6416 1974
rect 6388 1947 6389 1973
rect 6389 1947 6415 1973
rect 6415 1947 6416 1973
rect 6388 1946 6416 1947
rect 6440 1973 6468 1974
rect 6440 1947 6441 1973
rect 6441 1947 6467 1973
rect 6467 1947 6468 1973
rect 6440 1946 6468 1947
rect 6492 1973 6520 1974
rect 6492 1947 6493 1973
rect 6493 1947 6519 1973
rect 6519 1947 6520 1973
rect 6492 1946 6520 1947
rect 5334 1833 5362 1834
rect 5334 1807 5335 1833
rect 5335 1807 5361 1833
rect 5361 1807 5362 1833
rect 5334 1806 5362 1807
rect 5562 1581 5590 1582
rect 5562 1555 5563 1581
rect 5563 1555 5589 1581
rect 5589 1555 5590 1581
rect 5562 1554 5590 1555
rect 5614 1581 5642 1582
rect 5614 1555 5615 1581
rect 5615 1555 5641 1581
rect 5641 1555 5642 1581
rect 5614 1554 5642 1555
rect 5666 1581 5694 1582
rect 5666 1555 5667 1581
rect 5667 1555 5693 1581
rect 5693 1555 5694 1581
rect 5666 1554 5694 1555
rect 7214 1581 7242 1582
rect 7214 1555 7215 1581
rect 7215 1555 7241 1581
rect 7241 1555 7242 1581
rect 7214 1554 7242 1555
rect 7266 1581 7294 1582
rect 7266 1555 7267 1581
rect 7267 1555 7293 1581
rect 7293 1555 7294 1581
rect 7266 1554 7294 1555
rect 7318 1581 7346 1582
rect 7318 1555 7319 1581
rect 7319 1555 7345 1581
rect 7345 1555 7346 1581
rect 7318 1554 7346 1555
<< metal3 >>
rect 7600 7098 8000 7112
rect 3593 7070 3598 7098
rect 3626 7070 8000 7098
rect 7600 7056 8000 7070
rect 7600 6762 8000 6776
rect 5833 6734 5838 6762
rect 5866 6734 8000 6762
rect 7600 6720 8000 6734
rect 7600 6426 8000 6440
rect 6337 6398 6342 6426
rect 6370 6398 8000 6426
rect 7600 6384 8000 6398
rect 2253 6258 2258 6286
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2390 6258 2395 6286
rect 3905 6258 3910 6286
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 4042 6258 4047 6286
rect 5557 6258 5562 6286
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5694 6258 5699 6286
rect 7209 6258 7214 6286
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7346 6258 7351 6286
rect 4041 6174 4046 6202
rect 4074 6174 6790 6202
rect 6818 6174 6823 6202
rect 3425 6118 3430 6146
rect 3458 6118 4382 6146
rect 4410 6118 4415 6146
rect 7600 6090 8000 6104
rect 3761 6062 3766 6090
rect 3794 6062 4718 6090
rect 4746 6062 4751 6090
rect 6225 6062 6230 6090
rect 6258 6062 8000 6090
rect 7600 6048 8000 6062
rect 3201 5950 3206 5978
rect 3234 5950 3934 5978
rect 3962 5950 5082 5978
rect 1427 5866 1432 5894
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1564 5866 1569 5894
rect 3079 5866 3084 5894
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3216 5866 3221 5894
rect 4731 5866 4736 5894
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4868 5866 4873 5894
rect 5054 5754 5082 5950
rect 6383 5866 6388 5894
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6520 5866 6525 5894
rect 7600 5754 8000 5768
rect 5054 5726 8000 5754
rect 7600 5712 8000 5726
rect 4321 5670 4326 5698
rect 4354 5670 4774 5698
rect 4802 5670 4807 5698
rect 4881 5670 4886 5698
rect 4914 5670 5222 5698
rect 5250 5670 6734 5698
rect 6762 5670 6958 5698
rect 6986 5670 6991 5698
rect 2253 5474 2258 5502
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2390 5474 2395 5502
rect 3905 5474 3910 5502
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 4042 5474 4047 5502
rect 5557 5474 5562 5502
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5694 5474 5699 5502
rect 7209 5474 7214 5502
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7346 5474 7351 5502
rect 7600 5418 8000 5432
rect 4209 5390 4214 5418
rect 4242 5390 4494 5418
rect 4522 5390 8000 5418
rect 7600 5376 8000 5390
rect 3985 5334 3990 5362
rect 4018 5334 4942 5362
rect 4970 5334 5726 5362
rect 5754 5334 5759 5362
rect 3705 5222 3710 5250
rect 3738 5222 4046 5250
rect 4074 5222 5278 5250
rect 5306 5222 5311 5250
rect 5777 5222 5782 5250
rect 5810 5222 6566 5250
rect 6594 5222 6599 5250
rect 5609 5166 5614 5194
rect 5642 5166 6846 5194
rect 6874 5166 6879 5194
rect 1427 5082 1432 5110
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1564 5082 1569 5110
rect 3079 5082 3084 5110
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3216 5082 3221 5110
rect 4731 5082 4736 5110
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4868 5082 4873 5110
rect 6383 5082 6388 5110
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6520 5082 6525 5110
rect 7600 5082 8000 5096
rect 6678 5054 8000 5082
rect 6678 5026 6706 5054
rect 7600 5040 8000 5054
rect 6673 4998 6678 5026
rect 6706 4998 6711 5026
rect 4209 4830 4214 4858
rect 4242 4830 4942 4858
rect 4970 4830 4975 4858
rect 4993 4774 4998 4802
rect 5026 4774 6734 4802
rect 6762 4774 6767 4802
rect 0 4746 400 4760
rect 7600 4746 8000 4760
rect 0 4718 854 4746
rect 882 4718 1246 4746
rect 1274 4718 1279 4746
rect 0 4704 400 4718
rect 2253 4690 2258 4718
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2390 4690 2395 4718
rect 3905 4690 3910 4718
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 4042 4690 4047 4718
rect 5557 4690 5562 4718
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5694 4690 5699 4718
rect 7209 4690 7214 4718
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7346 4690 7351 4718
rect 7574 4704 8000 4746
rect 7574 4634 7602 4704
rect 5833 4606 5838 4634
rect 5866 4606 7602 4634
rect 4377 4494 4382 4522
rect 4410 4494 4718 4522
rect 4746 4494 4751 4522
rect 5889 4494 5894 4522
rect 5922 4494 6958 4522
rect 6986 4494 6991 4522
rect 4881 4438 4886 4466
rect 4914 4438 5222 4466
rect 5250 4438 5255 4466
rect 0 4410 400 4424
rect 7600 4410 8000 4424
rect 0 4382 854 4410
rect 882 4382 1246 4410
rect 1274 4382 1279 4410
rect 6617 4382 6622 4410
rect 6650 4382 8000 4410
rect 0 4368 400 4382
rect 7600 4368 8000 4382
rect 1427 4298 1432 4326
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1564 4298 1569 4326
rect 3079 4298 3084 4326
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3216 4298 3221 4326
rect 4731 4298 4736 4326
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4868 4298 4873 4326
rect 6383 4298 6388 4326
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6520 4298 6525 4326
rect 4881 4214 4886 4242
rect 4914 4214 5166 4242
rect 5194 4214 5894 4242
rect 5922 4214 5927 4242
rect 4993 4158 4998 4186
rect 5026 4158 6846 4186
rect 6874 4158 6879 4186
rect 5385 4102 5390 4130
rect 5418 4102 7014 4130
rect 7042 4102 7047 4130
rect 0 4074 400 4088
rect 7600 4074 8000 4088
rect 0 4046 854 4074
rect 882 4046 1806 4074
rect 1834 4046 1839 4074
rect 6337 4046 6342 4074
rect 6370 4046 8000 4074
rect 0 4032 400 4046
rect 7600 4032 8000 4046
rect 2253 3906 2258 3934
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2390 3906 2395 3934
rect 3905 3906 3910 3934
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 4042 3906 4047 3934
rect 5557 3906 5562 3934
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5694 3906 5699 3934
rect 7209 3906 7214 3934
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7346 3906 7351 3934
rect 6785 3822 6790 3850
rect 6818 3822 6958 3850
rect 6986 3822 6991 3850
rect 1073 3766 1078 3794
rect 1106 3766 2870 3794
rect 2898 3766 2903 3794
rect 0 3738 400 3752
rect 7600 3738 8000 3752
rect 0 3710 1302 3738
rect 1330 3710 1335 3738
rect 4489 3710 4494 3738
rect 4522 3710 5894 3738
rect 5922 3710 5927 3738
rect 6673 3710 6678 3738
rect 6706 3710 8000 3738
rect 0 3696 400 3710
rect 7600 3696 8000 3710
rect 905 3654 910 3682
rect 938 3654 1750 3682
rect 1778 3654 1783 3682
rect 6281 3654 6286 3682
rect 6314 3654 6790 3682
rect 6818 3654 6823 3682
rect 1427 3514 1432 3542
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1564 3514 1569 3542
rect 3079 3514 3084 3542
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3216 3514 3221 3542
rect 4731 3514 4736 3542
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4868 3514 4873 3542
rect 6383 3514 6388 3542
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6520 3514 6525 3542
rect 0 3402 400 3416
rect 7600 3402 8000 3416
rect 0 3374 910 3402
rect 938 3374 943 3402
rect 6281 3374 6286 3402
rect 6314 3374 8000 3402
rect 0 3360 400 3374
rect 7600 3360 8000 3374
rect 1073 3318 1078 3346
rect 1106 3318 2198 3346
rect 2226 3318 2231 3346
rect 4881 3318 4886 3346
rect 4914 3318 5222 3346
rect 5250 3318 5255 3346
rect 4993 3262 4998 3290
rect 5026 3262 6846 3290
rect 6874 3262 6879 3290
rect 4041 3206 4046 3234
rect 4074 3206 5166 3234
rect 5194 3206 5199 3234
rect 5278 3206 6902 3234
rect 6930 3206 6935 3234
rect 5278 3178 5306 3206
rect 4657 3150 4662 3178
rect 4690 3150 5306 3178
rect 2253 3122 2258 3150
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2390 3122 2395 3150
rect 3905 3122 3910 3150
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 4042 3122 4047 3150
rect 5557 3122 5562 3150
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5694 3122 5699 3150
rect 7209 3122 7214 3150
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7346 3122 7351 3150
rect 0 3066 400 3080
rect 7600 3066 8000 3080
rect 0 3038 854 3066
rect 882 3038 887 3066
rect 7065 3038 7070 3066
rect 7098 3038 8000 3066
rect 0 3024 400 3038
rect 7600 3024 8000 3038
rect 3649 2982 3654 3010
rect 3682 2982 4158 3010
rect 4186 2982 4191 3010
rect 1017 2926 1022 2954
rect 1050 2926 2366 2954
rect 2394 2926 2399 2954
rect 5217 2814 5222 2842
rect 5250 2814 6286 2842
rect 6314 2814 6319 2842
rect 0 2730 400 2744
rect 1427 2730 1432 2758
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1564 2730 1569 2758
rect 3079 2730 3084 2758
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3216 2730 3221 2758
rect 4731 2730 4736 2758
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4868 2730 4873 2758
rect 6383 2730 6388 2758
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6520 2730 6525 2758
rect 7600 2730 8000 2744
rect 0 2702 1190 2730
rect 1218 2702 1223 2730
rect 6561 2702 6566 2730
rect 6594 2702 8000 2730
rect 0 2688 400 2702
rect 7600 2688 8000 2702
rect 961 2646 966 2674
rect 994 2646 2982 2674
rect 3010 2646 3015 2674
rect 3705 2646 3710 2674
rect 3738 2646 4774 2674
rect 4802 2646 4807 2674
rect 849 2590 854 2618
rect 882 2590 1806 2618
rect 1834 2590 1839 2618
rect 1185 2534 1190 2562
rect 1218 2534 1582 2562
rect 1610 2534 1615 2562
rect 3929 2534 3934 2562
rect 3962 2534 4270 2562
rect 4298 2534 4942 2562
rect 4970 2534 4975 2562
rect 0 2394 400 2408
rect 0 2366 854 2394
rect 882 2366 1246 2394
rect 1274 2366 1279 2394
rect 0 2352 400 2366
rect 2253 2338 2258 2366
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2390 2338 2395 2366
rect 3905 2338 3910 2366
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 4042 2338 4047 2366
rect 5557 2338 5562 2366
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5694 2338 5699 2366
rect 7209 2338 7214 2366
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7346 2338 7351 2366
rect 1353 2254 1358 2282
rect 1386 2254 2534 2282
rect 2562 2254 2567 2282
rect 4097 2254 4102 2282
rect 4130 2254 6902 2282
rect 6930 2254 6935 2282
rect 0 2058 400 2072
rect 0 2030 1190 2058
rect 1218 2030 1582 2058
rect 1610 2030 1615 2058
rect 4377 2030 4382 2058
rect 4410 2030 5278 2058
rect 5306 2030 5311 2058
rect 0 2016 400 2030
rect 1427 1946 1432 1974
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1564 1946 1569 1974
rect 3079 1946 3084 1974
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3216 1946 3221 1974
rect 4731 1946 4736 1974
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4868 1946 4873 1974
rect 6383 1946 6388 1974
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6520 1946 6525 1974
rect 4713 1806 4718 1834
rect 4746 1806 5334 1834
rect 5362 1806 5367 1834
rect 3537 1750 3542 1778
rect 3570 1750 3934 1778
rect 3962 1750 3967 1778
rect 4097 1750 4102 1778
rect 4130 1750 4270 1778
rect 4298 1750 4303 1778
rect 0 1722 400 1736
rect 0 1694 854 1722
rect 882 1694 1470 1722
rect 1498 1694 1503 1722
rect 0 1680 400 1694
rect 2253 1554 2258 1582
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2390 1554 2395 1582
rect 3905 1554 3910 1582
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 4042 1554 4047 1582
rect 5557 1554 5562 1582
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5694 1554 5699 1582
rect 7209 1554 7214 1582
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7346 1554 7351 1582
<< via3 >>
rect 2258 6258 2286 6286
rect 2310 6258 2338 6286
rect 2362 6258 2390 6286
rect 3910 6258 3938 6286
rect 3962 6258 3990 6286
rect 4014 6258 4042 6286
rect 5562 6258 5590 6286
rect 5614 6258 5642 6286
rect 5666 6258 5694 6286
rect 7214 6258 7242 6286
rect 7266 6258 7294 6286
rect 7318 6258 7346 6286
rect 1432 5866 1460 5894
rect 1484 5866 1512 5894
rect 1536 5866 1564 5894
rect 3084 5866 3112 5894
rect 3136 5866 3164 5894
rect 3188 5866 3216 5894
rect 4736 5866 4764 5894
rect 4788 5866 4816 5894
rect 4840 5866 4868 5894
rect 6388 5866 6416 5894
rect 6440 5866 6468 5894
rect 6492 5866 6520 5894
rect 2258 5474 2286 5502
rect 2310 5474 2338 5502
rect 2362 5474 2390 5502
rect 3910 5474 3938 5502
rect 3962 5474 3990 5502
rect 4014 5474 4042 5502
rect 5562 5474 5590 5502
rect 5614 5474 5642 5502
rect 5666 5474 5694 5502
rect 7214 5474 7242 5502
rect 7266 5474 7294 5502
rect 7318 5474 7346 5502
rect 1432 5082 1460 5110
rect 1484 5082 1512 5110
rect 1536 5082 1564 5110
rect 3084 5082 3112 5110
rect 3136 5082 3164 5110
rect 3188 5082 3216 5110
rect 4736 5082 4764 5110
rect 4788 5082 4816 5110
rect 4840 5082 4868 5110
rect 6388 5082 6416 5110
rect 6440 5082 6468 5110
rect 6492 5082 6520 5110
rect 2258 4690 2286 4718
rect 2310 4690 2338 4718
rect 2362 4690 2390 4718
rect 3910 4690 3938 4718
rect 3962 4690 3990 4718
rect 4014 4690 4042 4718
rect 5562 4690 5590 4718
rect 5614 4690 5642 4718
rect 5666 4690 5694 4718
rect 7214 4690 7242 4718
rect 7266 4690 7294 4718
rect 7318 4690 7346 4718
rect 1432 4298 1460 4326
rect 1484 4298 1512 4326
rect 1536 4298 1564 4326
rect 3084 4298 3112 4326
rect 3136 4298 3164 4326
rect 3188 4298 3216 4326
rect 4736 4298 4764 4326
rect 4788 4298 4816 4326
rect 4840 4298 4868 4326
rect 6388 4298 6416 4326
rect 6440 4298 6468 4326
rect 6492 4298 6520 4326
rect 2258 3906 2286 3934
rect 2310 3906 2338 3934
rect 2362 3906 2390 3934
rect 3910 3906 3938 3934
rect 3962 3906 3990 3934
rect 4014 3906 4042 3934
rect 5562 3906 5590 3934
rect 5614 3906 5642 3934
rect 5666 3906 5694 3934
rect 7214 3906 7242 3934
rect 7266 3906 7294 3934
rect 7318 3906 7346 3934
rect 1432 3514 1460 3542
rect 1484 3514 1512 3542
rect 1536 3514 1564 3542
rect 3084 3514 3112 3542
rect 3136 3514 3164 3542
rect 3188 3514 3216 3542
rect 4736 3514 4764 3542
rect 4788 3514 4816 3542
rect 4840 3514 4868 3542
rect 6388 3514 6416 3542
rect 6440 3514 6468 3542
rect 6492 3514 6520 3542
rect 2258 3122 2286 3150
rect 2310 3122 2338 3150
rect 2362 3122 2390 3150
rect 3910 3122 3938 3150
rect 3962 3122 3990 3150
rect 4014 3122 4042 3150
rect 5562 3122 5590 3150
rect 5614 3122 5642 3150
rect 5666 3122 5694 3150
rect 7214 3122 7242 3150
rect 7266 3122 7294 3150
rect 7318 3122 7346 3150
rect 1432 2730 1460 2758
rect 1484 2730 1512 2758
rect 1536 2730 1564 2758
rect 3084 2730 3112 2758
rect 3136 2730 3164 2758
rect 3188 2730 3216 2758
rect 4736 2730 4764 2758
rect 4788 2730 4816 2758
rect 4840 2730 4868 2758
rect 6388 2730 6416 2758
rect 6440 2730 6468 2758
rect 6492 2730 6520 2758
rect 2258 2338 2286 2366
rect 2310 2338 2338 2366
rect 2362 2338 2390 2366
rect 3910 2338 3938 2366
rect 3962 2338 3990 2366
rect 4014 2338 4042 2366
rect 5562 2338 5590 2366
rect 5614 2338 5642 2366
rect 5666 2338 5694 2366
rect 7214 2338 7242 2366
rect 7266 2338 7294 2366
rect 7318 2338 7346 2366
rect 1432 1946 1460 1974
rect 1484 1946 1512 1974
rect 1536 1946 1564 1974
rect 3084 1946 3112 1974
rect 3136 1946 3164 1974
rect 3188 1946 3216 1974
rect 4736 1946 4764 1974
rect 4788 1946 4816 1974
rect 4840 1946 4868 1974
rect 6388 1946 6416 1974
rect 6440 1946 6468 1974
rect 6492 1946 6520 1974
rect 2258 1554 2286 1582
rect 2310 1554 2338 1582
rect 2362 1554 2390 1582
rect 3910 1554 3938 1582
rect 3962 1554 3990 1582
rect 4014 1554 4042 1582
rect 5562 1554 5590 1582
rect 5614 1554 5642 1582
rect 5666 1554 5694 1582
rect 7214 1554 7242 1582
rect 7266 1554 7294 1582
rect 7318 1554 7346 1582
<< metal4 >>
rect 1418 5894 1578 6302
rect 1418 5866 1432 5894
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1564 5866 1578 5894
rect 1418 5110 1578 5866
rect 1418 5082 1432 5110
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1564 5082 1578 5110
rect 1418 4326 1578 5082
rect 1418 4298 1432 4326
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1564 4298 1578 4326
rect 1418 3542 1578 4298
rect 1418 3514 1432 3542
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1564 3514 1578 3542
rect 1418 2758 1578 3514
rect 1418 2730 1432 2758
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1564 2730 1578 2758
rect 1418 1974 1578 2730
rect 1418 1946 1432 1974
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1564 1946 1578 1974
rect 1418 1538 1578 1946
rect 2244 6286 2404 6302
rect 2244 6258 2258 6286
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2390 6258 2404 6286
rect 2244 5502 2404 6258
rect 2244 5474 2258 5502
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2390 5474 2404 5502
rect 2244 4718 2404 5474
rect 2244 4690 2258 4718
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2390 4690 2404 4718
rect 2244 3934 2404 4690
rect 2244 3906 2258 3934
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2390 3906 2404 3934
rect 2244 3150 2404 3906
rect 2244 3122 2258 3150
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2390 3122 2404 3150
rect 2244 2366 2404 3122
rect 2244 2338 2258 2366
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2390 2338 2404 2366
rect 2244 1582 2404 2338
rect 2244 1554 2258 1582
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2390 1554 2404 1582
rect 2244 1538 2404 1554
rect 3070 5894 3230 6302
rect 3070 5866 3084 5894
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3216 5866 3230 5894
rect 3070 5110 3230 5866
rect 3070 5082 3084 5110
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3216 5082 3230 5110
rect 3070 4326 3230 5082
rect 3070 4298 3084 4326
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3216 4298 3230 4326
rect 3070 3542 3230 4298
rect 3070 3514 3084 3542
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3216 3514 3230 3542
rect 3070 2758 3230 3514
rect 3070 2730 3084 2758
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3216 2730 3230 2758
rect 3070 1974 3230 2730
rect 3070 1946 3084 1974
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3216 1946 3230 1974
rect 3070 1538 3230 1946
rect 3896 6286 4056 6302
rect 3896 6258 3910 6286
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 4042 6258 4056 6286
rect 3896 5502 4056 6258
rect 3896 5474 3910 5502
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 4042 5474 4056 5502
rect 3896 4718 4056 5474
rect 3896 4690 3910 4718
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 4042 4690 4056 4718
rect 3896 3934 4056 4690
rect 3896 3906 3910 3934
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 4042 3906 4056 3934
rect 3896 3150 4056 3906
rect 3896 3122 3910 3150
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 4042 3122 4056 3150
rect 3896 2366 4056 3122
rect 3896 2338 3910 2366
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 4042 2338 4056 2366
rect 3896 1582 4056 2338
rect 3896 1554 3910 1582
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 4042 1554 4056 1582
rect 3896 1538 4056 1554
rect 4722 5894 4882 6302
rect 4722 5866 4736 5894
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4868 5866 4882 5894
rect 4722 5110 4882 5866
rect 4722 5082 4736 5110
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4868 5082 4882 5110
rect 4722 4326 4882 5082
rect 4722 4298 4736 4326
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4868 4298 4882 4326
rect 4722 3542 4882 4298
rect 4722 3514 4736 3542
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4868 3514 4882 3542
rect 4722 2758 4882 3514
rect 4722 2730 4736 2758
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4868 2730 4882 2758
rect 4722 1974 4882 2730
rect 4722 1946 4736 1974
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4868 1946 4882 1974
rect 4722 1538 4882 1946
rect 5548 6286 5708 6302
rect 5548 6258 5562 6286
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5694 6258 5708 6286
rect 5548 5502 5708 6258
rect 5548 5474 5562 5502
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5694 5474 5708 5502
rect 5548 4718 5708 5474
rect 5548 4690 5562 4718
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5694 4690 5708 4718
rect 5548 3934 5708 4690
rect 5548 3906 5562 3934
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5694 3906 5708 3934
rect 5548 3150 5708 3906
rect 5548 3122 5562 3150
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5694 3122 5708 3150
rect 5548 2366 5708 3122
rect 5548 2338 5562 2366
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5694 2338 5708 2366
rect 5548 1582 5708 2338
rect 5548 1554 5562 1582
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5694 1554 5708 1582
rect 5548 1538 5708 1554
rect 6374 5894 6534 6302
rect 6374 5866 6388 5894
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6520 5866 6534 5894
rect 6374 5110 6534 5866
rect 6374 5082 6388 5110
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6520 5082 6534 5110
rect 6374 4326 6534 5082
rect 6374 4298 6388 4326
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6520 4298 6534 4326
rect 6374 3542 6534 4298
rect 6374 3514 6388 3542
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6520 3514 6534 3542
rect 6374 2758 6534 3514
rect 6374 2730 6388 2758
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6520 2730 6534 2758
rect 6374 1974 6534 2730
rect 6374 1946 6388 1974
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6520 1946 6534 1974
rect 6374 1538 6534 1946
rect 7200 6286 7360 6302
rect 7200 6258 7214 6286
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7346 6258 7360 6286
rect 7200 5502 7360 6258
rect 7200 5474 7214 5502
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7346 5474 7360 5502
rect 7200 4718 7360 5474
rect 7200 4690 7214 4718
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7346 4690 7360 4718
rect 7200 3934 7360 4690
rect 7200 3906 7214 3934
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7346 3906 7360 3934
rect 7200 3150 7360 3906
rect 7200 3122 7214 3150
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7346 3122 7360 3150
rect 7200 2366 7360 3122
rect 7200 2338 7214 2366
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7346 2338 7360 2366
rect 7200 1582 7360 2338
rect 7200 1554 7214 1582
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7346 1554 7360 1582
rect 7200 1538 7360 1554
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _16_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 784 0 -1 3136
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _17_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 952 0 -1 3920
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _18_
timestamp 1698431365
transform -1 0 2744 0 -1 3136
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _19_
timestamp 1698431365
transform 1 0 1288 0 1 3136
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _20_
timestamp 1698431365
transform 1 0 2744 0 1 3136
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _21_
timestamp 1698431365
transform 1 0 2296 0 -1 3920
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _22_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3584 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _23_
timestamp 1698431365
transform -1 0 4424 0 -1 3920
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _24_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3472 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _25_
timestamp 1698431365
transform 1 0 3304 0 -1 3136
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _26_
timestamp 1698431365
transform 1 0 4872 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _27_
timestamp 1698431365
transform 1 0 4872 0 -1 3920
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _28_
timestamp 1698431365
transform 1 0 5376 0 -1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _29_
timestamp 1698431365
transform 1 0 3808 0 1 3136
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _30_
timestamp 1698431365
transform 1 0 6664 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _31_
timestamp 1698431365
transform -1 0 5376 0 -1 4704
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _32_
timestamp 1698431365
transform 1 0 4256 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _33_
timestamp 1698431365
transform 1 0 3808 0 1 4704
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _34_
timestamp 1698431365
transform 1 0 6664 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _35_
timestamp 1698431365
transform 1 0 5040 0 -1 5488
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _36_
timestamp 1698431365
transform -1 0 7000 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _37_
timestamp 1698431365
transform 1 0 3808 0 1 3920
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _38_
timestamp 1698431365
transform 1 0 6664 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _39_
timestamp 1698431365
transform -1 0 7168 0 -1 6272
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _40_
timestamp 1698431365
transform -1 0 5712 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _41_
timestamp 1698431365
transform 1 0 3808 0 1 5488
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _42_
timestamp 1698431365
transform -1 0 7000 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _43_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3192 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__43__I test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3080 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 1736 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 3416 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 6664 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 7168 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 3808 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 3472 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 3584 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 4256 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 3248 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 4032 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 1456 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 1232 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 1232 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 1792 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 1232 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 1792 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 1568 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 1568 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 4088 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 1568 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_8 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1120 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_12
timestamp 1698431365
transform 1 0 1344 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_16 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_32
timestamp 1698431365
transform 1 0 2464 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_36 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_44
timestamp 1698431365
transform 1 0 3136 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_46 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3248 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 4424 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_72
timestamp 1698431365
transform 1 0 4704 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_99
timestamp 1698431365
transform 1 0 6216 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 6328 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_104
timestamp 1698431365
transform 1 0 6496 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_112
timestamp 1698431365
transform 1 0 6944 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_14
timestamp 1698431365
transform 1 0 1456 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_18
timestamp 1698431365
transform 1 0 1680 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_34
timestamp 1698431365
transform 1 0 2576 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_42
timestamp 1698431365
transform 1 0 3024 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_51
timestamp 1698431365
transform 1 0 3528 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_61
timestamp 1698431365
transform 1 0 4088 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 4536 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_98 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6160 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_102
timestamp 1698431365
transform 1 0 6384 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_104
timestamp 1698431365
transform 1 0 6496 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_107
timestamp 1698431365
transform 1 0 6664 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_109
timestamp 1698431365
transform 1 0 6776 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_14
timestamp 1698431365
transform 1 0 1456 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_18
timestamp 1698431365
transform 1 0 1680 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_22
timestamp 1698431365
transform 1 0 1904 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_30
timestamp 1698431365
transform 1 0 2352 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_37
timestamp 1698431365
transform 1 0 2744 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_45
timestamp 1698431365
transform 1 0 3192 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_49
timestamp 1698431365
transform 1 0 3416 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_51
timestamp 1698431365
transform 1 0 3528 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_60 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4032 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_92
timestamp 1698431365
transform 1 0 5824 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_96
timestamp 1698431365
transform 1 0 6048 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_98
timestamp 1698431365
transform 1 0 6160 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_113
timestamp 1698431365
transform 1 0 7000 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_115
timestamp 1698431365
transform 1 0 7112 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_37
timestamp 1698431365
transform 1 0 2744 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_45
timestamp 1698431365
transform 1 0 3192 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 4704 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_74
timestamp 1698431365
transform 1 0 4816 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_83
timestamp 1698431365
transform 1 0 5320 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_8
timestamp 1698431365
transform 1 0 1120 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_10
timestamp 1698431365
transform 1 0 1232 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_49
timestamp 1698431365
transform 1 0 3416 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_113
timestamp 1698431365
transform 1 0 7000 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_115
timestamp 1698431365
transform 1 0 7112 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698431365
transform 1 0 784 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_4
timestamp 1698431365
transform 1 0 896 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_17
timestamp 1698431365
transform 1 0 1624 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_21
timestamp 1698431365
transform 1 0 1848 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_52
timestamp 1698431365
transform 1 0 3584 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_54
timestamp 1698431365
transform 1 0 3696 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_67
timestamp 1698431365
transform 1 0 4424 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 4536 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 4704 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_74
timestamp 1698431365
transform 1 0 4816 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_87
timestamp 1698431365
transform 1 0 5544 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_89
timestamp 1698431365
transform 1 0 5656 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_14
timestamp 1698431365
transform 1 0 1456 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_18
timestamp 1698431365
transform 1 0 1680 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_22
timestamp 1698431365
transform 1 0 1904 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_30
timestamp 1698431365
transform 1 0 2352 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_37
timestamp 1698431365
transform 1 0 2744 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_53
timestamp 1698431365
transform 1 0 3640 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_55
timestamp 1698431365
transform 1 0 3752 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_115
timestamp 1698431365
transform 1 0 7112 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_8
timestamp 1698431365
transform 1 0 1120 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_12
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_44
timestamp 1698431365
transform 1 0 3136 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_60
timestamp 1698431365
transform 1 0 4032 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1698431365
transform 1 0 1120 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_12
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 2744 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_53
timestamp 1698431365
transform 1 0 3640 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_55
timestamp 1698431365
transform 1 0 3752 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_115
timestamp 1698431365
transform 1 0 7112 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 784 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_34
timestamp 1698431365
transform 1 0 2576 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_50
timestamp 1698431365
transform 1 0 3472 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_60
timestamp 1698431365
transform 1 0 4032 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_37
timestamp 1698431365
transform 1 0 2744 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_45
timestamp 1698431365
transform 1 0 3192 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_49
timestamp 1698431365
transform 1 0 3416 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_52
timestamp 1698431365
transform 1 0 3584 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_115
timestamp 1698431365
transform 1 0 7112 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_2
timestamp 1698431365
transform 1 0 784 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_36
timestamp 1698431365
transform 1 0 2688 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_46
timestamp 1698431365
transform 1 0 3248 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 784 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 4088 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 6552 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 7168 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 4592 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 4480 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 3472 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 4592 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 3808 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 5040 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 784 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 784 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 784 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 784 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 784 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 784 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 1120 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 1120 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 4424 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 1456 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output21
timestamp 1698431365
transform -1 0 3752 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4928 0 -1 6272
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform -1 0 7168 0 -1 5488
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698431365
transform 1 0 4760 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698431365
transform 1 0 4704 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698431365
transform 1 0 5096 0 1 3136
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1698431365
transform 1 0 5712 0 -1 3136
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698431365
transform 1 0 5096 0 1 3920
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output29
timestamp 1698431365
transform 1 0 5712 0 -1 3920
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output30
timestamp 1698431365
transform 1 0 5712 0 -1 4704
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output31
timestamp 1698431365
transform -1 0 6552 0 1 4704
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output32
timestamp 1698431365
transform 1 0 5096 0 1 5488
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_12 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 7280 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_13
timestamp 1698431365
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 7280 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_14
timestamp 1698431365
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 7280 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_15
timestamp 1698431365
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 7280 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_16
timestamp 1698431365
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 7280 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_17
timestamp 1698431365
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 7280 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_18
timestamp 1698431365
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 7280 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_19
timestamp 1698431365
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 7280 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_20
timestamp 1698431365
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 7280 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_21
timestamp 1698431365
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 7280 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_22
timestamp 1698431365
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 7280 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_23
timestamp 1698431365
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 7280 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_24 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_25
timestamp 1698431365
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_26
timestamp 1698431365
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_27
timestamp 1698431365
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_28
timestamp 1698431365
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_29
timestamp 1698431365
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_30
timestamp 1698431365
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_31
timestamp 1698431365
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_32
timestamp 1698431365
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_33
timestamp 1698431365
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_34
timestamp 1698431365
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_35
timestamp 1698431365
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_36
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_37
timestamp 1698431365
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_38
timestamp 1698431365
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_39
timestamp 1698431365
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_40
timestamp 1698431365
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_41
timestamp 1698431365
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_42
timestamp 1698431365
transform 1 0 2576 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_43
timestamp 1698431365
transform 1 0 4480 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_44
timestamp 1698431365
transform 1 0 6384 0 -1 6272
box -43 -43 155 435
<< labels >>
flabel metal2 s 3024 0 3080 400 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 3360 400 3416 0 FreeSans 224 0 0 0 in[0]
port 1 nsew signal input
flabel metal2 s 3696 0 3752 400 0 FreeSans 224 90 0 0 in[10]
port 2 nsew signal input
flabel metal3 s 7600 2688 8000 2744 0 FreeSans 224 0 0 0 in[11]
port 3 nsew signal input
flabel metal3 s 7600 3024 8000 3080 0 FreeSans 224 0 0 0 in[12]
port 4 nsew signal input
flabel metal2 s 4704 7600 4760 8000 0 FreeSans 224 90 0 0 in[13]
port 5 nsew signal input
flabel metal2 s 4368 7600 4424 8000 0 FreeSans 224 90 0 0 in[14]
port 6 nsew signal input
flabel metal3 s 7600 7056 8000 7112 0 FreeSans 224 0 0 0 in[15]
port 7 nsew signal input
flabel metal3 s 7600 5376 8000 5432 0 FreeSans 224 0 0 0 in[16]
port 8 nsew signal input
flabel metal3 s 7600 5712 8000 5768 0 FreeSans 224 0 0 0 in[17]
port 9 nsew signal input
flabel metal2 s 5712 7600 5768 8000 0 FreeSans 224 90 0 0 in[18]
port 10 nsew signal input
flabel metal3 s 0 1680 400 1736 0 FreeSans 224 0 0 0 in[1]
port 11 nsew signal input
flabel metal3 s 0 4368 400 4424 0 FreeSans 224 0 0 0 in[2]
port 12 nsew signal input
flabel metal3 s 0 2352 400 2408 0 FreeSans 224 0 0 0 in[3]
port 13 nsew signal input
flabel metal3 s 0 3024 400 3080 0 FreeSans 224 0 0 0 in[4]
port 14 nsew signal input
flabel metal3 s 0 4704 400 4760 0 FreeSans 224 0 0 0 in[5]
port 15 nsew signal input
flabel metal3 s 0 4032 400 4088 0 FreeSans 224 0 0 0 in[6]
port 16 nsew signal input
flabel metal3 s 0 2016 400 2072 0 FreeSans 224 0 0 0 in[7]
port 17 nsew signal input
flabel metal3 s 0 2688 400 2744 0 FreeSans 224 0 0 0 in[8]
port 18 nsew signal input
flabel metal2 s 4032 0 4088 400 0 FreeSans 224 90 0 0 in[9]
port 19 nsew signal input
flabel metal2 s 3360 0 3416 400 0 FreeSans 224 90 0 0 out[0]
port 20 nsew signal tristate
flabel metal3 s 7600 6720 8000 6776 0 FreeSans 224 0 0 0 out[10]
port 21 nsew signal tristate
flabel metal3 s 7600 6384 8000 6440 0 FreeSans 224 0 0 0 out[11]
port 22 nsew signal tristate
flabel metal2 s 4704 0 4760 400 0 FreeSans 224 90 0 0 out[1]
port 23 nsew signal tristate
flabel metal2 s 4368 0 4424 400 0 FreeSans 224 90 0 0 out[2]
port 24 nsew signal tristate
flabel metal3 s 7600 3360 8000 3416 0 FreeSans 224 0 0 0 out[3]
port 25 nsew signal tristate
flabel metal3 s 7600 3696 8000 3752 0 FreeSans 224 0 0 0 out[4]
port 26 nsew signal tristate
flabel metal3 s 7600 4032 8000 4088 0 FreeSans 224 0 0 0 out[5]
port 27 nsew signal tristate
flabel metal3 s 7600 4368 8000 4424 0 FreeSans 224 0 0 0 out[6]
port 28 nsew signal tristate
flabel metal3 s 7600 5040 8000 5096 0 FreeSans 224 0 0 0 out[7]
port 29 nsew signal tristate
flabel metal3 s 7600 4704 8000 4760 0 FreeSans 224 0 0 0 out[8]
port 30 nsew signal tristate
flabel metal3 s 7600 6048 8000 6104 0 FreeSans 224 0 0 0 out[9]
port 31 nsew signal tristate
flabel metal3 s 0 3696 400 3752 0 FreeSans 224 0 0 0 rst_n
port 32 nsew signal input
flabel metal4 s 1418 1538 1578 6302 0 FreeSans 640 90 0 0 vdd
port 33 nsew power bidirectional
flabel metal4 s 3070 1538 3230 6302 0 FreeSans 640 90 0 0 vdd
port 33 nsew power bidirectional
flabel metal4 s 4722 1538 4882 6302 0 FreeSans 640 90 0 0 vdd
port 33 nsew power bidirectional
flabel metal4 s 6374 1538 6534 6302 0 FreeSans 640 90 0 0 vdd
port 33 nsew power bidirectional
flabel metal4 s 2244 1538 2404 6302 0 FreeSans 640 90 0 0 vss
port 34 nsew ground bidirectional
flabel metal4 s 3896 1538 4056 6302 0 FreeSans 640 90 0 0 vss
port 34 nsew ground bidirectional
flabel metal4 s 5548 1538 5708 6302 0 FreeSans 640 90 0 0 vss
port 34 nsew ground bidirectional
flabel metal4 s 7200 1538 7360 6302 0 FreeSans 640 90 0 0 vss
port 34 nsew ground bidirectional
rlabel metal1 3976 5880 3976 5880 0 vdd
rlabel via1 4016 6272 4016 6272 0 vss
rlabel metal2 1820 3164 1820 3164 0 _00_
rlabel metal2 1540 3640 1540 3640 0 _01_
rlabel metal2 2156 3164 2156 3164 0 _02_
rlabel metal2 2492 3500 2492 3500 0 _03_
rlabel metal2 3332 3584 3332 3584 0 _04_
rlabel metal2 3584 2548 3584 2548 0 _05_
rlabel metal2 3612 3500 3612 3500 0 _06_
rlabel metal2 4732 2940 4732 2940 0 _07_
rlabel metal2 5460 3332 5460 3332 0 _08_
rlabel metal3 5936 3276 5936 3276 0 _09_
rlabel metal2 4788 4480 4788 4480 0 _10_
rlabel metal2 5012 4816 5012 4816 0 _11_
rlabel metal2 6944 2548 6944 2548 0 _12_
rlabel metal3 5936 4172 5936 4172 0 _13_
rlabel metal2 5684 4564 5684 4564 0 _14_
rlabel metal2 4844 5376 4844 5376 0 _15_
rlabel metal2 3024 1428 3024 1428 0 clk
rlabel metal2 924 3500 924 3500 0 in[0]
rlabel metal2 3640 1092 3640 1092 0 in[10]
rlabel metal2 6468 2576 6468 2576 0 in[11]
rlabel metal2 7084 2632 7084 2632 0 in[12]
rlabel metal2 4732 6853 4732 6853 0 in[13]
rlabel metal2 4396 6881 4396 6881 0 in[14]
rlabel metal2 3612 6580 3612 6580 0 in[15]
rlabel metal2 4508 5376 4508 5376 0 in[16]
rlabel metal2 3948 6020 3948 6020 0 in[17]
rlabel metal3 5348 5348 5348 5348 0 in[18]
rlabel metal3 623 1708 623 1708 0 in[1]
rlabel metal2 868 4452 868 4452 0 in[2]
rlabel metal2 868 2296 868 2296 0 in[3]
rlabel metal2 868 2800 868 2800 0 in[4]
rlabel metal2 868 4788 868 4788 0 in[5]
rlabel metal3 623 4060 623 4060 0 in[6]
rlabel metal2 1204 2100 1204 2100 0 in[7]
rlabel metal2 1204 2632 1204 2632 0 in[8]
rlabel metal2 4088 1484 4088 1484 0 in[9]
rlabel metal2 1092 3220 1092 3220 0 net1
rlabel metal2 4788 5544 4788 5544 0 net10
rlabel metal2 1064 1708 1064 1708 0 net11
rlabel metal2 980 3542 980 3542 0 net12
rlabel metal2 1008 2268 1008 2268 0 net13
rlabel metal2 1036 2716 1036 2716 0 net14
rlabel metal2 1064 4788 1064 4788 0 net15
rlabel metal2 1092 3444 1092 3444 0 net16
rlabel metal2 2548 3024 2548 3024 0 net17
rlabel metal2 1372 2716 1372 2716 0 net18
rlabel metal3 3920 2996 3920 2996 0 net19
rlabel metal2 3836 2324 3836 2324 0 net2
rlabel metal2 1176 4004 1176 4004 0 net20
rlabel metal2 3612 1988 3612 1988 0 net21
rlabel metal2 5460 5348 5460 5348 0 net22
rlabel metal2 6748 3556 6748 3556 0 net23
rlabel metal3 4452 2548 4452 2548 0 net24
rlabel metal2 3724 2940 3724 2940 0 net25
rlabel metal2 5236 3500 5236 3500 0 net26
rlabel metal2 5628 2968 5628 2968 0 net27
rlabel metal3 6216 4116 6216 4116 0 net28
rlabel metal2 4508 4144 4508 4144 0 net29
rlabel metal2 5180 3276 5180 3276 0 net3
rlabel metal2 5908 4368 5908 4368 0 net30
rlabel metal2 6748 2828 6748 2828 0 net31
rlabel metal3 5068 5684 5068 5684 0 net32
rlabel metal3 5516 2268 5516 2268 0 net4
rlabel metal2 4984 4508 4984 4508 0 net5
rlabel metal2 4256 6132 4256 6132 0 net6
rlabel metal2 4116 4648 4116 4648 0 net7
rlabel metal2 4340 4732 4340 4732 0 net8
rlabel metal3 5432 6188 5432 6188 0 net9
rlabel metal2 3388 1015 3388 1015 0 out[0]
rlabel metal2 5852 6440 5852 6440 0 out[10]
rlabel metal2 6300 5880 6300 5880 0 out[11]
rlabel metal3 5040 1820 5040 1820 0 out[1]
rlabel metal3 4844 2044 4844 2044 0 out[2]
rlabel metal3 6965 3388 6965 3388 0 out[3]
rlabel metal2 6692 3360 6692 3360 0 out[4]
rlabel metal2 6356 4116 6356 4116 0 out[5]
rlabel metal2 6636 4088 6636 4088 0 out[6]
rlabel metal2 6692 4788 6692 4788 0 out[7]
rlabel metal3 7609 4732 7609 4732 0 out[8]
rlabel metal2 6244 5908 6244 5908 0 out[9]
rlabel metal2 1316 3920 1316 3920 0 rst_n
<< properties >>
string FIXED_BBOX 0 0 8000 8000
<< end >>
