VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO output_mux
  CLASS BLOCK ;
  FOREIGN output_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 70.560 200.000 71.120 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 4.000 98.000 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 196.000 74.480 200.000 ;
    END
  END out[11]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 77.280 200.000 77.840 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 120.960 200.000 121.520 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 107.520 200.000 108.080 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 0.000 121.520 4.000 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 196.000 84.560 200.000 ;
    END
  END out[9]
  PIN proj_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 94.080 200.000 94.640 ;
    END
  END proj_out[0]
  PIN proj_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END proj_out[10]
  PIN proj_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 196.000 94.640 200.000 ;
    END
  END proj_out[11]
  PIN proj_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 100.800 200.000 101.360 ;
    END
  END proj_out[12]
  PIN proj_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 87.360 200.000 87.920 ;
    END
  END proj_out[13]
  PIN proj_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 110.880 200.000 111.440 ;
    END
  END proj_out[14]
  PIN proj_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 117.600 200.000 118.160 ;
    END
  END proj_out[15]
  PIN proj_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END proj_out[16]
  PIN proj_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END proj_out[17]
  PIN proj_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END proj_out[18]
  PIN proj_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END proj_out[19]
  PIN proj_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 84.000 200.000 84.560 ;
    END
  END proj_out[1]
  PIN proj_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END proj_out[20]
  PIN proj_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 196.000 91.280 200.000 ;
    END
  END proj_out[21]
  PIN proj_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END proj_out[22]
  PIN proj_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 196.000 87.920 200.000 ;
    END
  END proj_out[23]
  PIN proj_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 97.440 200.000 98.000 ;
    END
  END proj_out[24]
  PIN proj_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 90.720 200.000 91.280 ;
    END
  END proj_out[25]
  PIN proj_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 196.000 104.720 200.000 ;
    END
  END proj_out[26]
  PIN proj_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 196.000 101.360 200.000 ;
    END
  END proj_out[27]
  PIN proj_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 4.000 77.840 ;
    END
  END proj_out[28]
  PIN proj_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END proj_out[29]
  PIN proj_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 114.240 200.000 114.800 ;
    END
  END proj_out[2]
  PIN proj_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END proj_out[30]
  PIN proj_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END proj_out[31]
  PIN proj_out[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END proj_out[32]
  PIN proj_out[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END proj_out[33]
  PIN proj_out[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END proj_out[34]
  PIN proj_out[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END proj_out[35]
  PIN proj_out[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 73.920 200.000 74.480 ;
    END
  END proj_out[36]
  PIN proj_out[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 80.640 200.000 81.200 ;
    END
  END proj_out[37]
  PIN proj_out[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 196.000 111.440 200.000 ;
    END
  END proj_out[38]
  PIN proj_out[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 196.000 108.080 200.000 ;
    END
  END proj_out[39]
  PIN proj_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 104.160 200.000 104.720 ;
    END
  END proj_out[3]
  PIN proj_out[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.640 4.000 81.200 ;
    END
  END proj_out[40]
  PIN proj_out[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END proj_out[41]
  PIN proj_out[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END proj_out[42]
  PIN proj_out[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END proj_out[43]
  PIN proj_out[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END proj_out[44]
  PIN proj_out[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 196.000 77.840 200.000 ;
    END
  END proj_out[45]
  PIN proj_out[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END proj_out[46]
  PIN proj_out[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 196.000 81.200 200.000 ;
    END
  END proj_out[47]
  PIN proj_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END proj_out[4]
  PIN proj_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END proj_out[5]
  PIN proj_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END proj_out[6]
  PIN proj_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 0.000 67.760 4.000 ;
    END
  END proj_out[7]
  PIN proj_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END proj_out[8]
  PIN proj_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 196.000 98.000 200.000 ;
    END
  END proj_out[9]
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END sel[1]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 29.230 15.380 30.830 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 75.850 15.380 77.450 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.470 15.380 124.070 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.090 15.380 170.690 184.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 52.540 15.380 54.140 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.160 15.380 100.760 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 145.780 15.380 147.380 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 192.400 15.380 194.000 184.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 194.000 184.540 ;
      LAYER Metal2 ;
        RECT 8.540 195.700 73.620 196.000 ;
        RECT 74.780 195.700 76.980 196.000 ;
        RECT 78.140 195.700 80.340 196.000 ;
        RECT 81.500 195.700 83.700 196.000 ;
        RECT 84.860 195.700 87.060 196.000 ;
        RECT 88.220 195.700 90.420 196.000 ;
        RECT 91.580 195.700 93.780 196.000 ;
        RECT 94.940 195.700 97.140 196.000 ;
        RECT 98.300 195.700 100.500 196.000 ;
        RECT 101.660 195.700 103.860 196.000 ;
        RECT 105.020 195.700 107.220 196.000 ;
        RECT 108.380 195.700 110.580 196.000 ;
        RECT 111.740 195.700 193.860 196.000 ;
        RECT 8.540 4.300 193.860 195.700 ;
        RECT 8.540 4.000 63.540 4.300 ;
        RECT 64.700 4.000 66.900 4.300 ;
        RECT 68.060 4.000 70.260 4.300 ;
        RECT 71.420 4.000 73.620 4.300 ;
        RECT 74.780 4.000 76.980 4.300 ;
        RECT 78.140 4.000 80.340 4.300 ;
        RECT 81.500 4.000 83.700 4.300 ;
        RECT 84.860 4.000 87.060 4.300 ;
        RECT 88.220 4.000 90.420 4.300 ;
        RECT 91.580 4.000 93.780 4.300 ;
        RECT 94.940 4.000 97.140 4.300 ;
        RECT 98.300 4.000 100.500 4.300 ;
        RECT 101.660 4.000 103.860 4.300 ;
        RECT 105.020 4.000 107.220 4.300 ;
        RECT 108.380 4.000 110.580 4.300 ;
        RECT 111.740 4.000 113.940 4.300 ;
        RECT 115.100 4.000 117.300 4.300 ;
        RECT 118.460 4.000 120.660 4.300 ;
        RECT 121.820 4.000 193.860 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 128.540 196.000 184.380 ;
        RECT 4.300 127.380 196.000 128.540 ;
        RECT 4.000 125.180 196.000 127.380 ;
        RECT 4.300 124.020 196.000 125.180 ;
        RECT 4.000 121.820 196.000 124.020 ;
        RECT 4.300 120.660 195.700 121.820 ;
        RECT 4.000 118.460 196.000 120.660 ;
        RECT 4.300 117.300 195.700 118.460 ;
        RECT 4.000 115.100 196.000 117.300 ;
        RECT 4.300 113.940 195.700 115.100 ;
        RECT 4.000 111.740 196.000 113.940 ;
        RECT 4.300 110.580 195.700 111.740 ;
        RECT 4.000 108.380 196.000 110.580 ;
        RECT 4.300 107.220 195.700 108.380 ;
        RECT 4.000 105.020 196.000 107.220 ;
        RECT 4.300 103.860 195.700 105.020 ;
        RECT 4.000 101.660 196.000 103.860 ;
        RECT 4.300 100.500 195.700 101.660 ;
        RECT 4.000 98.300 196.000 100.500 ;
        RECT 4.300 97.140 195.700 98.300 ;
        RECT 4.000 94.940 196.000 97.140 ;
        RECT 4.300 93.780 195.700 94.940 ;
        RECT 4.000 91.580 196.000 93.780 ;
        RECT 4.300 90.420 195.700 91.580 ;
        RECT 4.000 88.220 196.000 90.420 ;
        RECT 4.300 87.060 195.700 88.220 ;
        RECT 4.000 84.860 196.000 87.060 ;
        RECT 4.300 83.700 195.700 84.860 ;
        RECT 4.000 81.500 196.000 83.700 ;
        RECT 4.300 80.340 195.700 81.500 ;
        RECT 4.000 78.140 196.000 80.340 ;
        RECT 4.300 76.980 195.700 78.140 ;
        RECT 4.000 74.780 196.000 76.980 ;
        RECT 4.000 73.620 195.700 74.780 ;
        RECT 4.000 71.420 196.000 73.620 ;
        RECT 4.000 70.260 195.700 71.420 ;
        RECT 4.000 15.540 196.000 70.260 ;
  END
END output_mux
END LIBRARY

