magic
tech gf180mcuD
magscale 1 5
timestamp 1702441055
<< obsm1 >>
rect 672 463 39312 38625
<< metal2 >>
rect 0 39600 56 40000
rect 336 39600 392 40000
rect 672 39600 728 40000
rect 1008 39600 1064 40000
rect 1344 39600 1400 40000
rect 1680 39600 1736 40000
rect 2016 39600 2072 40000
rect 2352 39600 2408 40000
rect 2688 39600 2744 40000
rect 3024 39600 3080 40000
rect 3360 39600 3416 40000
rect 3696 39600 3752 40000
rect 4032 39600 4088 40000
rect 4368 39600 4424 40000
rect 4704 39600 4760 40000
rect 5040 39600 5096 40000
rect 5376 39600 5432 40000
rect 5712 39600 5768 40000
rect 6048 39600 6104 40000
rect 6384 39600 6440 40000
rect 6720 39600 6776 40000
rect 7056 39600 7112 40000
rect 7392 39600 7448 40000
rect 7728 39600 7784 40000
rect 8064 39600 8120 40000
rect 8400 39600 8456 40000
rect 8736 39600 8792 40000
rect 9072 39600 9128 40000
rect 9408 39600 9464 40000
rect 9744 39600 9800 40000
rect 10080 39600 10136 40000
rect 10416 39600 10472 40000
rect 10752 39600 10808 40000
rect 11088 39600 11144 40000
rect 11424 39600 11480 40000
rect 11760 39600 11816 40000
rect 12096 39600 12152 40000
rect 12432 39600 12488 40000
rect 12768 39600 12824 40000
rect 13104 39600 13160 40000
rect 13440 39600 13496 40000
rect 13776 39600 13832 40000
rect 14112 39600 14168 40000
rect 14448 39600 14504 40000
rect 14784 39600 14840 40000
rect 15120 39600 15176 40000
rect 15456 39600 15512 40000
rect 15792 39600 15848 40000
rect 16128 39600 16184 40000
rect 16464 39600 16520 40000
rect 16800 39600 16856 40000
rect 17136 39600 17192 40000
rect 17472 39600 17528 40000
rect 17808 39600 17864 40000
rect 18144 39600 18200 40000
rect 18480 39600 18536 40000
rect 18816 39600 18872 40000
rect 19152 39600 19208 40000
rect 19488 39600 19544 40000
rect 19824 39600 19880 40000
rect 20160 39600 20216 40000
rect 20496 39600 20552 40000
rect 20832 39600 20888 40000
rect 21168 39600 21224 40000
rect 21504 39600 21560 40000
rect 21840 39600 21896 40000
rect 22176 39600 22232 40000
rect 22512 39600 22568 40000
rect 22848 39600 22904 40000
rect 23184 39600 23240 40000
rect 23520 39600 23576 40000
rect 23856 39600 23912 40000
rect 24192 39600 24248 40000
rect 24528 39600 24584 40000
rect 24864 39600 24920 40000
rect 25200 39600 25256 40000
rect 25536 39600 25592 40000
rect 25872 39600 25928 40000
rect 26208 39600 26264 40000
rect 26544 39600 26600 40000
rect 26880 39600 26936 40000
rect 27216 39600 27272 40000
rect 27552 39600 27608 40000
rect 27888 39600 27944 40000
rect 28224 39600 28280 40000
rect 28560 39600 28616 40000
rect 28896 39600 28952 40000
rect 29232 39600 29288 40000
rect 29568 39600 29624 40000
rect 29904 39600 29960 40000
rect 30240 39600 30296 40000
rect 30576 39600 30632 40000
rect 30912 39600 30968 40000
rect 31248 39600 31304 40000
rect 31584 39600 31640 40000
rect 31920 39600 31976 40000
rect 32256 39600 32312 40000
rect 32592 39600 32648 40000
rect 32928 39600 32984 40000
rect 33264 39600 33320 40000
rect 33600 39600 33656 40000
rect 33936 39600 33992 40000
rect 34272 39600 34328 40000
rect 34608 39600 34664 40000
rect 34944 39600 35000 40000
rect 35280 39600 35336 40000
rect 35616 39600 35672 40000
rect 35952 39600 36008 40000
rect 36288 39600 36344 40000
rect 36624 39600 36680 40000
rect 36960 39600 37016 40000
rect 37296 39600 37352 40000
rect 37632 39600 37688 40000
rect 37968 39600 38024 40000
rect 38304 39600 38360 40000
rect 38640 39600 38696 40000
rect 38976 39600 39032 40000
rect 39312 39600 39368 40000
rect 39648 39600 39704 40000
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
rect 5040 0 5096 400
rect 5376 0 5432 400
rect 5712 0 5768 400
rect 6048 0 6104 400
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12096 0 12152 400
rect 12432 0 12488 400
rect 12768 0 12824 400
rect 13104 0 13160 400
rect 13440 0 13496 400
rect 13776 0 13832 400
rect 14112 0 14168 400
rect 14448 0 14504 400
rect 14784 0 14840 400
rect 15120 0 15176 400
rect 15456 0 15512 400
rect 15792 0 15848 400
rect 16128 0 16184 400
rect 16464 0 16520 400
rect 16800 0 16856 400
rect 17136 0 17192 400
rect 17472 0 17528 400
rect 17808 0 17864 400
rect 18144 0 18200 400
rect 18480 0 18536 400
rect 18816 0 18872 400
rect 19152 0 19208 400
rect 19488 0 19544 400
rect 19824 0 19880 400
rect 20160 0 20216 400
rect 20496 0 20552 400
rect 20832 0 20888 400
rect 21168 0 21224 400
rect 21504 0 21560 400
rect 21840 0 21896 400
rect 22176 0 22232 400
rect 22512 0 22568 400
rect 22848 0 22904 400
rect 23184 0 23240 400
rect 23520 0 23576 400
rect 23856 0 23912 400
rect 24192 0 24248 400
rect 24528 0 24584 400
rect 24864 0 24920 400
rect 25200 0 25256 400
rect 25536 0 25592 400
rect 25872 0 25928 400
rect 26208 0 26264 400
rect 26544 0 26600 400
rect 26880 0 26936 400
rect 27216 0 27272 400
rect 27552 0 27608 400
rect 27888 0 27944 400
rect 28224 0 28280 400
rect 28560 0 28616 400
rect 28896 0 28952 400
rect 29232 0 29288 400
rect 29568 0 29624 400
rect 29904 0 29960 400
rect 30240 0 30296 400
rect 30576 0 30632 400
rect 30912 0 30968 400
rect 31248 0 31304 400
rect 31584 0 31640 400
rect 31920 0 31976 400
rect 32256 0 32312 400
rect 32592 0 32648 400
rect 32928 0 32984 400
rect 33264 0 33320 400
rect 33600 0 33656 400
rect 33936 0 33992 400
rect 34272 0 34328 400
rect 34608 0 34664 400
rect 34944 0 35000 400
rect 35280 0 35336 400
rect 35616 0 35672 400
rect 35952 0 36008 400
rect 36288 0 36344 400
rect 36624 0 36680 400
rect 36960 0 37016 400
rect 37296 0 37352 400
rect 37632 0 37688 400
rect 37968 0 38024 400
rect 38304 0 38360 400
rect 38640 0 38696 400
rect 38976 0 39032 400
rect 39312 0 39368 400
rect 39648 0 39704 400
<< obsm2 >>
rect 854 39570 978 39600
rect 1094 39570 1314 39600
rect 1430 39570 1650 39600
rect 1766 39570 1986 39600
rect 2102 39570 2322 39600
rect 2438 39570 2658 39600
rect 2774 39570 2994 39600
rect 3110 39570 3330 39600
rect 3446 39570 3666 39600
rect 3782 39570 4002 39600
rect 4118 39570 4338 39600
rect 4454 39570 4674 39600
rect 4790 39570 5010 39600
rect 5126 39570 5346 39600
rect 5462 39570 5682 39600
rect 5798 39570 6018 39600
rect 6134 39570 6354 39600
rect 6470 39570 6690 39600
rect 6806 39570 7026 39600
rect 7142 39570 7362 39600
rect 7478 39570 7698 39600
rect 7814 39570 8034 39600
rect 8150 39570 8370 39600
rect 8486 39570 8706 39600
rect 8822 39570 9042 39600
rect 9158 39570 9378 39600
rect 9494 39570 9714 39600
rect 9830 39570 10050 39600
rect 10166 39570 10386 39600
rect 10502 39570 10722 39600
rect 10838 39570 11058 39600
rect 11174 39570 11394 39600
rect 11510 39570 11730 39600
rect 11846 39570 12066 39600
rect 12182 39570 12402 39600
rect 12518 39570 12738 39600
rect 12854 39570 13074 39600
rect 13190 39570 13410 39600
rect 13526 39570 13746 39600
rect 13862 39570 14082 39600
rect 14198 39570 14418 39600
rect 14534 39570 14754 39600
rect 14870 39570 15090 39600
rect 15206 39570 15426 39600
rect 15542 39570 15762 39600
rect 15878 39570 16098 39600
rect 16214 39570 16434 39600
rect 16550 39570 16770 39600
rect 16886 39570 17106 39600
rect 17222 39570 17442 39600
rect 17558 39570 17778 39600
rect 17894 39570 18114 39600
rect 18230 39570 18450 39600
rect 18566 39570 18786 39600
rect 18902 39570 19122 39600
rect 19238 39570 19458 39600
rect 19574 39570 19794 39600
rect 19910 39570 20130 39600
rect 20246 39570 20466 39600
rect 20582 39570 20802 39600
rect 20918 39570 21138 39600
rect 21254 39570 21474 39600
rect 21590 39570 21810 39600
rect 21926 39570 22146 39600
rect 22262 39570 22482 39600
rect 22598 39570 22818 39600
rect 22934 39570 23154 39600
rect 23270 39570 23490 39600
rect 23606 39570 23826 39600
rect 23942 39570 24162 39600
rect 24278 39570 24498 39600
rect 24614 39570 24834 39600
rect 24950 39570 25170 39600
rect 25286 39570 25506 39600
rect 25622 39570 25842 39600
rect 25958 39570 26178 39600
rect 26294 39570 26514 39600
rect 26630 39570 26850 39600
rect 26966 39570 27186 39600
rect 27302 39570 27522 39600
rect 27638 39570 27858 39600
rect 27974 39570 28194 39600
rect 28310 39570 28530 39600
rect 28646 39570 28866 39600
rect 28982 39570 29202 39600
rect 29318 39570 29538 39600
rect 29654 39570 29874 39600
rect 29990 39570 30210 39600
rect 30326 39570 30546 39600
rect 30662 39570 30882 39600
rect 30998 39570 31218 39600
rect 31334 39570 31554 39600
rect 31670 39570 31890 39600
rect 32006 39570 32226 39600
rect 32342 39570 32562 39600
rect 32678 39570 32898 39600
rect 33014 39570 33234 39600
rect 33350 39570 33570 39600
rect 33686 39570 33906 39600
rect 34022 39570 34242 39600
rect 34358 39570 34578 39600
rect 34694 39570 34914 39600
rect 35030 39570 35250 39600
rect 35366 39570 35586 39600
rect 35702 39570 35922 39600
rect 36038 39570 36258 39600
rect 36374 39570 36594 39600
rect 36710 39570 36930 39600
rect 37046 39570 37266 39600
rect 37382 39570 37602 39600
rect 37718 39570 37938 39600
rect 38054 39570 38274 39600
rect 38390 39570 38610 39600
rect 38726 39570 38946 39600
rect 39062 39570 39242 39600
rect 854 430 39242 39570
rect 854 400 978 430
rect 1094 400 1314 430
rect 1430 400 1650 430
rect 1766 400 1986 430
rect 2102 400 2322 430
rect 2438 400 2658 430
rect 2774 400 2994 430
rect 3110 400 3330 430
rect 3446 400 3666 430
rect 3782 400 4002 430
rect 4118 400 4338 430
rect 4454 400 4674 430
rect 4790 400 5010 430
rect 5126 400 5346 430
rect 5462 400 5682 430
rect 5798 400 6018 430
rect 6134 400 6354 430
rect 6470 400 6690 430
rect 6806 400 7026 430
rect 7142 400 7362 430
rect 7478 400 7698 430
rect 7814 400 8034 430
rect 8150 400 8370 430
rect 8486 400 8706 430
rect 8822 400 9042 430
rect 9158 400 9378 430
rect 9494 400 9714 430
rect 9830 400 10050 430
rect 10166 400 10386 430
rect 10502 400 10722 430
rect 10838 400 11058 430
rect 11174 400 11394 430
rect 11510 400 11730 430
rect 11846 400 12066 430
rect 12182 400 12402 430
rect 12518 400 12738 430
rect 12854 400 13074 430
rect 13190 400 13410 430
rect 13526 400 13746 430
rect 13862 400 14082 430
rect 14198 400 14418 430
rect 14534 400 14754 430
rect 14870 400 15090 430
rect 15206 400 15426 430
rect 15542 400 15762 430
rect 15878 400 16098 430
rect 16214 400 16434 430
rect 16550 400 16770 430
rect 16886 400 17106 430
rect 17222 400 17442 430
rect 17558 400 17778 430
rect 17894 400 18114 430
rect 18230 400 18450 430
rect 18566 400 18786 430
rect 18902 400 19122 430
rect 19238 400 19458 430
rect 19574 400 19794 430
rect 19910 400 20130 430
rect 20246 400 20466 430
rect 20582 400 20802 430
rect 20918 400 21138 430
rect 21254 400 21474 430
rect 21590 400 21810 430
rect 21926 400 22146 430
rect 22262 400 22482 430
rect 22598 400 22818 430
rect 22934 400 23154 430
rect 23270 400 23490 430
rect 23606 400 23826 430
rect 23942 400 24162 430
rect 24278 400 24498 430
rect 24614 400 24834 430
rect 24950 400 25170 430
rect 25286 400 25506 430
rect 25622 400 25842 430
rect 25958 400 26178 430
rect 26294 400 26514 430
rect 26630 400 26850 430
rect 26966 400 27186 430
rect 27302 400 27522 430
rect 27638 400 27858 430
rect 27974 400 28194 430
rect 28310 400 28530 430
rect 28646 400 28866 430
rect 28982 400 29202 430
rect 29318 400 29538 430
rect 29654 400 29874 430
rect 29990 400 30210 430
rect 30326 400 30546 430
rect 30662 400 30882 430
rect 30998 400 31218 430
rect 31334 400 31554 430
rect 31670 400 31890 430
rect 32006 400 32226 430
rect 32342 400 32562 430
rect 32678 400 32898 430
rect 33014 400 33234 430
rect 33350 400 33570 430
rect 33686 400 33906 430
rect 34022 400 34242 430
rect 34358 400 34578 430
rect 34694 400 34914 430
rect 35030 400 35250 430
rect 35366 400 35586 430
rect 35702 400 35922 430
rect 36038 400 36258 430
rect 36374 400 36594 430
rect 36710 400 36930 430
rect 37046 400 37266 430
rect 37382 400 37602 430
rect 37718 400 37938 430
rect 38054 400 38274 430
rect 38390 400 38610 430
rect 38726 400 38946 430
rect 39062 400 39242 430
<< metal3 >>
rect 0 39648 400 39704
rect 39600 39648 40000 39704
rect 0 39312 400 39368
rect 39600 39312 40000 39368
rect 0 38976 400 39032
rect 39600 38976 40000 39032
rect 0 38640 400 38696
rect 39600 38640 40000 38696
rect 0 38304 400 38360
rect 39600 38304 40000 38360
rect 0 37968 400 38024
rect 39600 37968 40000 38024
rect 0 37632 400 37688
rect 39600 37632 40000 37688
rect 0 37296 400 37352
rect 39600 37296 40000 37352
rect 0 36960 400 37016
rect 39600 36960 40000 37016
rect 0 36624 400 36680
rect 39600 36624 40000 36680
rect 0 36288 400 36344
rect 39600 36288 40000 36344
rect 39600 35952 40000 36008
rect 39600 35616 40000 35672
rect 39600 35280 40000 35336
rect 39600 34944 40000 35000
rect 39600 34608 40000 34664
rect 39600 34272 40000 34328
rect 39600 33936 40000 33992
rect 0 33600 400 33656
rect 39600 33600 40000 33656
rect 0 33264 400 33320
rect 39600 33264 40000 33320
rect 0 32928 400 32984
rect 39600 32928 40000 32984
rect 0 32592 400 32648
rect 39600 32592 40000 32648
rect 0 32256 400 32312
rect 39600 32256 40000 32312
rect 0 31920 400 31976
rect 39600 31920 40000 31976
rect 0 31584 400 31640
rect 39600 31584 40000 31640
rect 0 31248 400 31304
rect 39600 31248 40000 31304
rect 0 30912 400 30968
rect 39600 30912 40000 30968
rect 0 30576 400 30632
rect 39600 30576 40000 30632
rect 0 30240 400 30296
rect 39600 30240 40000 30296
rect 0 29904 400 29960
rect 39600 29904 40000 29960
rect 0 29568 400 29624
rect 39600 29568 40000 29624
rect 0 29232 400 29288
rect 39600 29232 40000 29288
rect 0 28896 400 28952
rect 39600 28896 40000 28952
rect 0 28560 400 28616
rect 39600 28560 40000 28616
rect 0 28224 400 28280
rect 39600 28224 40000 28280
rect 0 27888 400 27944
rect 39600 27888 40000 27944
rect 0 27552 400 27608
rect 39600 27552 40000 27608
rect 0 27216 400 27272
rect 39600 27216 40000 27272
rect 0 26880 400 26936
rect 39600 26880 40000 26936
rect 0 26544 400 26600
rect 39600 26544 40000 26600
rect 0 26208 400 26264
rect 39600 26208 40000 26264
rect 0 25872 400 25928
rect 39600 25872 40000 25928
rect 0 25536 400 25592
rect 39600 25536 40000 25592
rect 0 25200 400 25256
rect 39600 25200 40000 25256
rect 0 24864 400 24920
rect 39600 24864 40000 24920
rect 0 24528 400 24584
rect 39600 24528 40000 24584
rect 0 24192 400 24248
rect 39600 24192 40000 24248
rect 0 23856 400 23912
rect 39600 23856 40000 23912
rect 0 23520 400 23576
rect 39600 23520 40000 23576
rect 0 23184 400 23240
rect 39600 23184 40000 23240
rect 0 22848 400 22904
rect 39600 22848 40000 22904
rect 0 22512 400 22568
rect 39600 22512 40000 22568
rect 0 22176 400 22232
rect 39600 22176 40000 22232
rect 0 21840 400 21896
rect 39600 21840 40000 21896
rect 0 21504 400 21560
rect 39600 21504 40000 21560
rect 0 21168 400 21224
rect 39600 21168 40000 21224
rect 0 20832 400 20888
rect 39600 20832 40000 20888
rect 0 20496 400 20552
rect 39600 20496 40000 20552
rect 0 20160 400 20216
rect 39600 20160 40000 20216
rect 0 19824 400 19880
rect 39600 19824 40000 19880
rect 0 19488 400 19544
rect 39600 19488 40000 19544
rect 0 19152 400 19208
rect 39600 19152 40000 19208
rect 0 18816 400 18872
rect 39600 18816 40000 18872
rect 0 18480 400 18536
rect 39600 18480 40000 18536
rect 0 18144 400 18200
rect 39600 18144 40000 18200
rect 0 17808 400 17864
rect 39600 17808 40000 17864
rect 0 17472 400 17528
rect 39600 17472 40000 17528
rect 0 17136 400 17192
rect 39600 17136 40000 17192
rect 0 16800 400 16856
rect 39600 16800 40000 16856
rect 0 16464 400 16520
rect 39600 16464 40000 16520
rect 0 16128 400 16184
rect 39600 16128 40000 16184
rect 0 15792 400 15848
rect 39600 15792 40000 15848
rect 0 15456 400 15512
rect 39600 15456 40000 15512
rect 0 15120 400 15176
rect 39600 15120 40000 15176
rect 0 14784 400 14840
rect 39600 14784 40000 14840
rect 0 14448 400 14504
rect 39600 14448 40000 14504
rect 0 14112 400 14168
rect 39600 14112 40000 14168
rect 0 13776 400 13832
rect 39600 13776 40000 13832
rect 0 13440 400 13496
rect 39600 13440 40000 13496
rect 0 13104 400 13160
rect 39600 13104 40000 13160
rect 0 12768 400 12824
rect 39600 12768 40000 12824
rect 0 12432 400 12488
rect 39600 12432 40000 12488
rect 0 12096 400 12152
rect 39600 12096 40000 12152
rect 0 11760 400 11816
rect 39600 11760 40000 11816
rect 0 11424 400 11480
rect 39600 11424 40000 11480
rect 0 11088 400 11144
rect 39600 11088 40000 11144
rect 0 10752 400 10808
rect 39600 10752 40000 10808
rect 0 10416 400 10472
rect 39600 10416 40000 10472
rect 0 10080 400 10136
rect 39600 10080 40000 10136
rect 0 9744 400 9800
rect 39600 9744 40000 9800
rect 0 9408 400 9464
rect 39600 9408 40000 9464
rect 0 9072 400 9128
rect 39600 9072 40000 9128
rect 0 8736 400 8792
rect 39600 8736 40000 8792
rect 0 8400 400 8456
rect 39600 8400 40000 8456
rect 0 8064 400 8120
rect 39600 8064 40000 8120
rect 0 7728 400 7784
rect 39600 7728 40000 7784
rect 0 7392 400 7448
rect 39600 7392 40000 7448
rect 0 7056 400 7112
rect 39600 7056 40000 7112
rect 0 6720 400 6776
rect 39600 6720 40000 6776
rect 0 6384 400 6440
rect 39600 6384 40000 6440
rect 0 6048 400 6104
rect 39600 6048 40000 6104
rect 39600 5712 40000 5768
rect 39600 5376 40000 5432
rect 39600 5040 40000 5096
rect 39600 4704 40000 4760
rect 39600 4368 40000 4424
rect 39600 4032 40000 4088
rect 39600 3696 40000 3752
rect 39600 3360 40000 3416
rect 39600 3024 40000 3080
rect 39600 2688 40000 2744
rect 39600 2352 40000 2408
rect 39600 2016 40000 2072
rect 39600 1680 40000 1736
rect 39600 1344 40000 1400
rect 39600 1008 40000 1064
rect 39600 672 40000 728
rect 39600 336 40000 392
rect 39600 0 40000 56
<< obsm3 >>
rect 430 38610 39570 38626
rect 400 38390 39600 38610
rect 430 38274 39570 38390
rect 400 38054 39600 38274
rect 430 37938 39570 38054
rect 400 37718 39600 37938
rect 430 37602 39570 37718
rect 400 37382 39600 37602
rect 430 37266 39570 37382
rect 400 37046 39600 37266
rect 430 36930 39570 37046
rect 400 36710 39600 36930
rect 430 36594 39570 36710
rect 400 36374 39600 36594
rect 430 36258 39570 36374
rect 400 36038 39600 36258
rect 400 35922 39570 36038
rect 400 35702 39600 35922
rect 400 35586 39570 35702
rect 400 35366 39600 35586
rect 400 35250 39570 35366
rect 400 35030 39600 35250
rect 400 34914 39570 35030
rect 400 34694 39600 34914
rect 400 34578 39570 34694
rect 400 34358 39600 34578
rect 400 34242 39570 34358
rect 400 34022 39600 34242
rect 400 33906 39570 34022
rect 400 33686 39600 33906
rect 430 33570 39570 33686
rect 400 33350 39600 33570
rect 430 33234 39570 33350
rect 400 33014 39600 33234
rect 430 32898 39570 33014
rect 400 32678 39600 32898
rect 430 32562 39570 32678
rect 400 32342 39600 32562
rect 430 32226 39570 32342
rect 400 32006 39600 32226
rect 430 31890 39570 32006
rect 400 31670 39600 31890
rect 430 31554 39570 31670
rect 400 31334 39600 31554
rect 430 31218 39570 31334
rect 400 30998 39600 31218
rect 430 30882 39570 30998
rect 400 30662 39600 30882
rect 430 30546 39570 30662
rect 400 30326 39600 30546
rect 430 30210 39570 30326
rect 400 29990 39600 30210
rect 430 29874 39570 29990
rect 400 29654 39600 29874
rect 430 29538 39570 29654
rect 400 29318 39600 29538
rect 430 29202 39570 29318
rect 400 28982 39600 29202
rect 430 28866 39570 28982
rect 400 28646 39600 28866
rect 430 28530 39570 28646
rect 400 28310 39600 28530
rect 430 28194 39570 28310
rect 400 27974 39600 28194
rect 430 27858 39570 27974
rect 400 27638 39600 27858
rect 430 27522 39570 27638
rect 400 27302 39600 27522
rect 430 27186 39570 27302
rect 400 26966 39600 27186
rect 430 26850 39570 26966
rect 400 26630 39600 26850
rect 430 26514 39570 26630
rect 400 26294 39600 26514
rect 430 26178 39570 26294
rect 400 25958 39600 26178
rect 430 25842 39570 25958
rect 400 25622 39600 25842
rect 430 25506 39570 25622
rect 400 25286 39600 25506
rect 430 25170 39570 25286
rect 400 24950 39600 25170
rect 430 24834 39570 24950
rect 400 24614 39600 24834
rect 430 24498 39570 24614
rect 400 24278 39600 24498
rect 430 24162 39570 24278
rect 400 23942 39600 24162
rect 430 23826 39570 23942
rect 400 23606 39600 23826
rect 430 23490 39570 23606
rect 400 23270 39600 23490
rect 430 23154 39570 23270
rect 400 22934 39600 23154
rect 430 22818 39570 22934
rect 400 22598 39600 22818
rect 430 22482 39570 22598
rect 400 22262 39600 22482
rect 430 22146 39570 22262
rect 400 21926 39600 22146
rect 430 21810 39570 21926
rect 400 21590 39600 21810
rect 430 21474 39570 21590
rect 400 21254 39600 21474
rect 430 21138 39570 21254
rect 400 20918 39600 21138
rect 430 20802 39570 20918
rect 400 20582 39600 20802
rect 430 20466 39570 20582
rect 400 20246 39600 20466
rect 430 20130 39570 20246
rect 400 19910 39600 20130
rect 430 19794 39570 19910
rect 400 19574 39600 19794
rect 430 19458 39570 19574
rect 400 19238 39600 19458
rect 430 19122 39570 19238
rect 400 18902 39600 19122
rect 430 18786 39570 18902
rect 400 18566 39600 18786
rect 430 18450 39570 18566
rect 400 18230 39600 18450
rect 430 18114 39570 18230
rect 400 17894 39600 18114
rect 430 17778 39570 17894
rect 400 17558 39600 17778
rect 430 17442 39570 17558
rect 400 17222 39600 17442
rect 430 17106 39570 17222
rect 400 16886 39600 17106
rect 430 16770 39570 16886
rect 400 16550 39600 16770
rect 430 16434 39570 16550
rect 400 16214 39600 16434
rect 430 16098 39570 16214
rect 400 15878 39600 16098
rect 430 15762 39570 15878
rect 400 15542 39600 15762
rect 430 15426 39570 15542
rect 400 15206 39600 15426
rect 430 15090 39570 15206
rect 400 14870 39600 15090
rect 430 14754 39570 14870
rect 400 14534 39600 14754
rect 430 14418 39570 14534
rect 400 14198 39600 14418
rect 430 14082 39570 14198
rect 400 13862 39600 14082
rect 430 13746 39570 13862
rect 400 13526 39600 13746
rect 430 13410 39570 13526
rect 400 13190 39600 13410
rect 430 13074 39570 13190
rect 400 12854 39600 13074
rect 430 12738 39570 12854
rect 400 12518 39600 12738
rect 430 12402 39570 12518
rect 400 12182 39600 12402
rect 430 12066 39570 12182
rect 400 11846 39600 12066
rect 430 11730 39570 11846
rect 400 11510 39600 11730
rect 430 11394 39570 11510
rect 400 11174 39600 11394
rect 430 11058 39570 11174
rect 400 10838 39600 11058
rect 430 10722 39570 10838
rect 400 10502 39600 10722
rect 430 10386 39570 10502
rect 400 10166 39600 10386
rect 430 10050 39570 10166
rect 400 9830 39600 10050
rect 430 9714 39570 9830
rect 400 9494 39600 9714
rect 430 9378 39570 9494
rect 400 9158 39600 9378
rect 430 9042 39570 9158
rect 400 8822 39600 9042
rect 430 8706 39570 8822
rect 400 8486 39600 8706
rect 430 8370 39570 8486
rect 400 8150 39600 8370
rect 430 8034 39570 8150
rect 400 7814 39600 8034
rect 430 7698 39570 7814
rect 400 7478 39600 7698
rect 430 7362 39570 7478
rect 400 7142 39600 7362
rect 430 7026 39570 7142
rect 400 6806 39600 7026
rect 430 6690 39570 6806
rect 400 6470 39600 6690
rect 430 6354 39570 6470
rect 400 6134 39600 6354
rect 430 6018 39570 6134
rect 400 5798 39600 6018
rect 400 5682 39570 5798
rect 400 5462 39600 5682
rect 400 5346 39570 5462
rect 400 5126 39600 5346
rect 400 5010 39570 5126
rect 400 4790 39600 5010
rect 400 4674 39570 4790
rect 400 4454 39600 4674
rect 400 4338 39570 4454
rect 400 4118 39600 4338
rect 400 4002 39570 4118
rect 400 3782 39600 4002
rect 400 3666 39570 3782
rect 400 3446 39600 3666
rect 400 3330 39570 3446
rect 400 3110 39600 3330
rect 400 2994 39570 3110
rect 400 2774 39600 2994
rect 400 2658 39570 2774
rect 400 2438 39600 2658
rect 400 2322 39570 2438
rect 400 2102 39600 2322
rect 400 1986 39570 2102
rect 400 1766 39600 1986
rect 400 1650 39570 1766
rect 400 1554 39600 1650
<< metal4 >>
rect 2224 1538 2384 38446
rect 9904 1538 10064 38446
rect 17584 1538 17744 38446
rect 25264 1538 25424 38446
rect 32944 1538 33104 38446
<< labels >>
rlabel metal3 s 39600 29232 40000 29288 6 clk
port 1 nsew signal output
rlabel metal3 s 39600 10080 40000 10136 6 in[0]
port 2 nsew signal output
rlabel metal3 s 39600 28896 40000 28952 6 in[10]
port 3 nsew signal output
rlabel metal3 s 0 33600 400 33656 6 in[11]
port 4 nsew signal output
rlabel metal2 s 25872 0 25928 400 6 in[12]
port 5 nsew signal output
rlabel metal2 s 11088 39600 11144 40000 6 in[13]
port 6 nsew signal output
rlabel metal3 s 0 6048 400 6104 6 in[14]
port 7 nsew signal output
rlabel metal2 s 25200 0 25256 400 6 in[15]
port 8 nsew signal output
rlabel metal2 s 13440 0 13496 400 6 in[16]
port 9 nsew signal output
rlabel metal2 s 29232 39600 29288 40000 6 in[17]
port 10 nsew signal output
rlabel metal2 s 25872 39600 25928 40000 6 in[1]
port 11 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 in[2]
port 12 nsew signal output
rlabel metal2 s 21504 0 21560 400 6 in[3]
port 13 nsew signal output
rlabel metal3 s 39600 12432 40000 12488 6 in[4]
port 14 nsew signal output
rlabel metal2 s 19152 39600 19208 40000 6 in[5]
port 15 nsew signal output
rlabel metal2 s 20160 39600 20216 40000 6 in[6]
port 16 nsew signal output
rlabel metal3 s 39600 10752 40000 10808 6 in[7]
port 17 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 in[8]
port 18 nsew signal output
rlabel metal3 s 0 14784 400 14840 6 in[9]
port 19 nsew signal output
rlabel metal2 s 2352 0 2408 400 6 io_in[0]
port 20 nsew signal input
rlabel metal2 s 20832 0 20888 400 6 io_in[10]
port 21 nsew signal input
rlabel metal2 s 20496 0 20552 400 6 io_in[11]
port 22 nsew signal input
rlabel metal3 s 39600 13104 40000 13160 6 io_in[12]
port 23 nsew signal input
rlabel metal2 s 18480 39600 18536 40000 6 io_in[13]
port 24 nsew signal input
rlabel metal2 s 17808 39600 17864 40000 6 io_in[14]
port 25 nsew signal input
rlabel metal3 s 39600 10416 40000 10472 6 io_in[15]
port 26 nsew signal input
rlabel metal3 s 0 18144 400 18200 6 io_in[16]
port 27 nsew signal input
rlabel metal3 s 0 16128 400 16184 6 io_in[17]
port 28 nsew signal input
rlabel metal3 s 39600 25536 40000 25592 6 io_in[18]
port 29 nsew signal input
rlabel metal3 s 0 32256 400 32312 6 io_in[19]
port 30 nsew signal input
rlabel metal2 s 32592 0 32648 400 6 io_in[1]
port 31 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 io_in[20]
port 32 nsew signal input
rlabel metal2 s 14112 39600 14168 40000 6 io_in[21]
port 33 nsew signal input
rlabel metal3 s 0 17136 400 17192 6 io_in[22]
port 34 nsew signal input
rlabel metal2 s 22176 0 22232 400 6 io_in[23]
port 35 nsew signal input
rlabel metal2 s 13776 0 13832 400 6 io_in[24]
port 36 nsew signal input
rlabel metal2 s 24192 39600 24248 40000 6 io_in[25]
port 37 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 io_in[26]
port 38 nsew signal input
rlabel metal2 s 33600 0 33656 400 6 io_in[27]
port 39 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 io_in[28]
port 40 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 io_in[29]
port 41 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 io_in[2]
port 42 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 io_in[30]
port 43 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 io_in[31]
port 44 nsew signal input
rlabel metal2 s 28224 0 28280 400 6 io_in[32]
port 45 nsew signal input
rlabel metal2 s 5376 0 5432 400 6 io_in[33]
port 46 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 io_in[34]
port 47 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 io_in[35]
port 48 nsew signal input
rlabel metal2 s 29232 0 29288 400 6 io_in[36]
port 49 nsew signal input
rlabel metal2 s 29904 0 29960 400 6 io_in[37]
port 50 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 io_in[3]
port 51 nsew signal input
rlabel metal2 s 38640 0 38696 400 6 io_in[4]
port 52 nsew signal input
rlabel metal2 s 14448 39600 14504 40000 6 io_in[5]
port 53 nsew signal input
rlabel metal3 s 39600 28224 40000 28280 6 io_in[6]
port 54 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 io_in[7]
port 55 nsew signal input
rlabel metal3 s 39600 16800 40000 16856 6 io_in[8]
port 56 nsew signal input
rlabel metal2 s 27216 39600 27272 40000 6 io_in[9]
port 57 nsew signal input
rlabel metal2 s 23184 39600 23240 40000 6 io_oeb[0]
port 58 nsew signal output
rlabel metal2 s 15792 39600 15848 40000 6 io_oeb[10]
port 59 nsew signal output
rlabel metal3 s 39600 28560 40000 28616 6 io_oeb[11]
port 60 nsew signal output
rlabel metal3 s 39600 26544 40000 26600 6 io_oeb[12]
port 61 nsew signal output
rlabel metal3 s 0 15120 400 15176 6 io_oeb[13]
port 62 nsew signal output
rlabel metal2 s 14448 0 14504 400 6 io_oeb[14]
port 63 nsew signal output
rlabel metal3 s 0 16464 400 16520 6 io_oeb[15]
port 64 nsew signal output
rlabel metal2 s 19824 0 19880 400 6 io_oeb[16]
port 65 nsew signal output
rlabel metal3 s 39600 17472 40000 17528 6 io_oeb[17]
port 66 nsew signal output
rlabel metal3 s 39600 19488 40000 19544 6 io_oeb[18]
port 67 nsew signal output
rlabel metal2 s 15120 0 15176 400 6 io_oeb[19]
port 68 nsew signal output
rlabel metal3 s 0 31920 400 31976 6 io_oeb[1]
port 69 nsew signal output
rlabel metal3 s 0 6720 400 6776 6 io_oeb[20]
port 70 nsew signal output
rlabel metal2 s 15792 0 15848 400 6 io_oeb[21]
port 71 nsew signal output
rlabel metal3 s 0 14448 400 14504 6 io_oeb[22]
port 72 nsew signal output
rlabel metal3 s 39600 15456 40000 15512 6 io_oeb[23]
port 73 nsew signal output
rlabel metal3 s 0 27216 400 27272 6 io_oeb[24]
port 74 nsew signal output
rlabel metal3 s 39600 17808 40000 17864 6 io_oeb[25]
port 75 nsew signal output
rlabel metal3 s 39600 20496 40000 20552 6 io_oeb[26]
port 76 nsew signal output
rlabel metal3 s 39600 16128 40000 16184 6 io_oeb[27]
port 77 nsew signal output
rlabel metal2 s 26544 39600 26600 40000 6 io_oeb[28]
port 78 nsew signal output
rlabel metal2 s 12432 39600 12488 40000 6 io_oeb[29]
port 79 nsew signal output
rlabel metal2 s 19488 39600 19544 40000 6 io_oeb[2]
port 80 nsew signal output
rlabel metal3 s 39600 22848 40000 22904 6 io_oeb[30]
port 81 nsew signal output
rlabel metal2 s 16464 0 16520 400 6 io_oeb[31]
port 82 nsew signal output
rlabel metal3 s 39600 12096 40000 12152 6 io_oeb[32]
port 83 nsew signal output
rlabel metal3 s 39600 21840 40000 21896 6 io_oeb[33]
port 84 nsew signal output
rlabel metal3 s 39600 21504 40000 21560 6 io_oeb[34]
port 85 nsew signal output
rlabel metal2 s 16128 39600 16184 40000 6 io_oeb[35]
port 86 nsew signal output
rlabel metal2 s 15456 39600 15512 40000 6 io_oeb[36]
port 87 nsew signal output
rlabel metal3 s 0 30912 400 30968 6 io_oeb[37]
port 88 nsew signal output
rlabel metal2 s 15120 39600 15176 40000 6 io_oeb[3]
port 89 nsew signal output
rlabel metal3 s 39600 19152 40000 19208 6 io_oeb[4]
port 90 nsew signal output
rlabel metal3 s 0 19824 400 19880 6 io_oeb[5]
port 91 nsew signal output
rlabel metal2 s 14784 0 14840 400 6 io_oeb[6]
port 92 nsew signal output
rlabel metal2 s 17136 39600 17192 40000 6 io_oeb[7]
port 93 nsew signal output
rlabel metal3 s 39600 26208 40000 26264 6 io_oeb[8]
port 94 nsew signal output
rlabel metal2 s 24528 39600 24584 40000 6 io_oeb[9]
port 95 nsew signal output
rlabel metal3 s 39600 18480 40000 18536 6 io_out[0]
port 96 nsew signal output
rlabel metal3 s 0 20160 400 20216 6 io_out[10]
port 97 nsew signal output
rlabel metal3 s 0 22512 400 22568 6 io_out[11]
port 98 nsew signal output
rlabel metal3 s 0 31248 400 31304 6 io_out[12]
port 99 nsew signal output
rlabel metal3 s 39600 24528 40000 24584 6 io_out[13]
port 100 nsew signal output
rlabel metal2 s 20160 0 20216 400 6 io_out[14]
port 101 nsew signal output
rlabel metal3 s 0 19488 400 19544 6 io_out[15]
port 102 nsew signal output
rlabel metal2 s 19152 0 19208 400 6 io_out[16]
port 103 nsew signal output
rlabel metal3 s 39600 18144 40000 18200 6 io_out[17]
port 104 nsew signal output
rlabel metal2 s 27552 39600 27608 40000 6 io_out[18]
port 105 nsew signal output
rlabel metal3 s 0 21168 400 21224 6 io_out[19]
port 106 nsew signal output
rlabel metal3 s 39600 18816 40000 18872 6 io_out[1]
port 107 nsew signal output
rlabel metal2 s 12768 39600 12824 40000 6 io_out[20]
port 108 nsew signal output
rlabel metal2 s 11424 39600 11480 40000 6 io_out[21]
port 109 nsew signal output
rlabel metal2 s 13440 39600 13496 40000 6 io_out[22]
port 110 nsew signal output
rlabel metal2 s 15456 0 15512 400 6 io_out[23]
port 111 nsew signal output
rlabel metal3 s 39600 16464 40000 16520 6 io_out[24]
port 112 nsew signal output
rlabel metal2 s 23184 0 23240 400 6 io_out[25]
port 113 nsew signal output
rlabel metal3 s 39600 15120 40000 15176 6 io_out[26]
port 114 nsew signal output
rlabel metal3 s 0 20832 400 20888 6 io_out[27]
port 115 nsew signal output
rlabel metal3 s 39600 26880 40000 26936 6 io_out[28]
port 116 nsew signal output
rlabel metal3 s 0 15456 400 15512 6 io_out[29]
port 117 nsew signal output
rlabel metal3 s 39600 20160 40000 20216 6 io_out[2]
port 118 nsew signal output
rlabel metal2 s 20496 39600 20552 40000 6 io_out[30]
port 119 nsew signal output
rlabel metal3 s 39600 23520 40000 23576 6 io_out[31]
port 120 nsew signal output
rlabel metal2 s 16800 0 16856 400 6 io_out[32]
port 121 nsew signal output
rlabel metal2 s 13776 39600 13832 40000 6 io_out[33]
port 122 nsew signal output
rlabel metal3 s 39600 12768 40000 12824 6 io_out[34]
port 123 nsew signal output
rlabel metal3 s 39600 11424 40000 11480 6 io_out[35]
port 124 nsew signal output
rlabel metal2 s 24864 39600 24920 40000 6 io_out[36]
port 125 nsew signal output
rlabel metal3 s 0 22176 400 22232 6 io_out[37]
port 126 nsew signal output
rlabel metal3 s 39600 27888 40000 27944 6 io_out[3]
port 127 nsew signal output
rlabel metal3 s 39600 27552 40000 27608 6 io_out[4]
port 128 nsew signal output
rlabel metal3 s 39600 22176 40000 22232 6 io_out[5]
port 129 nsew signal output
rlabel metal2 s 25536 0 25592 400 6 io_out[6]
port 130 nsew signal output
rlabel metal3 s 39600 24864 40000 24920 6 io_out[7]
port 131 nsew signal output
rlabel metal2 s 22848 39600 22904 40000 6 io_out[8]
port 132 nsew signal output
rlabel metal3 s 39600 19824 40000 19880 6 io_out[9]
port 133 nsew signal output
rlabel metal2 s 9744 0 9800 400 6 la_data_in[0]
port 134 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 la_data_in[10]
port 135 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 la_data_in[11]
port 136 nsew signal input
rlabel metal2 s 27552 0 27608 400 6 la_data_in[12]
port 137 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 la_data_in[13]
port 138 nsew signal input
rlabel metal2 s 33936 0 33992 400 6 la_data_in[14]
port 139 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 la_data_in[15]
port 140 nsew signal input
rlabel metal2 s 37296 0 37352 400 6 la_data_in[16]
port 141 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 la_data_in[17]
port 142 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 la_data_in[18]
port 143 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 la_data_in[19]
port 144 nsew signal input
rlabel metal2 s 39312 0 39368 400 6 la_data_in[1]
port 145 nsew signal input
rlabel metal2 s 336 0 392 400 6 la_data_in[20]
port 146 nsew signal input
rlabel metal2 s 672 0 728 400 6 la_data_in[21]
port 147 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 la_data_in[22]
port 148 nsew signal input
rlabel metal2 s 10752 0 10808 400 6 la_data_in[23]
port 149 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 la_data_in[24]
port 150 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 la_data_in[25]
port 151 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 la_data_in[26]
port 152 nsew signal input
rlabel metal2 s 39648 0 39704 400 6 la_data_in[27]
port 153 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 la_data_in[28]
port 154 nsew signal input
rlabel metal2 s 12432 0 12488 400 6 la_data_in[29]
port 155 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 la_data_in[2]
port 156 nsew signal input
rlabel metal2 s 0 0 56 400 6 la_data_in[30]
port 157 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 la_data_in[31]
port 158 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 la_data_in[32]
port 159 nsew signal input
rlabel metal2 s 26880 0 26936 400 6 la_data_in[33]
port 160 nsew signal input
rlabel metal2 s 35952 0 36008 400 6 la_data_in[34]
port 161 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 la_data_in[35]
port 162 nsew signal input
rlabel metal2 s 28896 0 28952 400 6 la_data_in[36]
port 163 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 la_data_in[37]
port 164 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 la_data_in[38]
port 165 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 la_data_in[39]
port 166 nsew signal input
rlabel metal2 s 32256 0 32312 400 6 la_data_in[3]
port 167 nsew signal input
rlabel metal2 s 12096 0 12152 400 6 la_data_in[40]
port 168 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 la_data_in[41]
port 169 nsew signal input
rlabel metal2 s 36288 0 36344 400 6 la_data_in[42]
port 170 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 la_data_in[43]
port 171 nsew signal input
rlabel metal2 s 5712 0 5768 400 6 la_data_in[44]
port 172 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 la_data_in[45]
port 173 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 la_data_in[46]
port 174 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 la_data_in[47]
port 175 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 la_data_in[48]
port 176 nsew signal input
rlabel metal2 s 31584 0 31640 400 6 la_data_in[49]
port 177 nsew signal input
rlabel metal2 s 34944 0 35000 400 6 la_data_in[4]
port 178 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 la_data_in[50]
port 179 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 la_data_in[51]
port 180 nsew signal input
rlabel metal2 s 36960 0 37016 400 6 la_data_in[52]
port 181 nsew signal input
rlabel metal2 s 37632 0 37688 400 6 la_data_in[53]
port 182 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 la_data_in[54]
port 183 nsew signal input
rlabel metal2 s 26544 0 26600 400 6 la_data_in[55]
port 184 nsew signal input
rlabel metal2 s 35616 0 35672 400 6 la_data_in[56]
port 185 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 la_data_in[57]
port 186 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 la_data_in[58]
port 187 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 la_data_in[59]
port 188 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 la_data_in[5]
port 189 nsew signal input
rlabel metal2 s 37968 0 38024 400 6 la_data_in[60]
port 190 nsew signal input
rlabel metal2 s 30912 0 30968 400 6 la_data_in[61]
port 191 nsew signal input
rlabel metal2 s 35280 0 35336 400 6 la_data_in[62]
port 192 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 la_data_in[63]
port 193 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 la_data_in[6]
port 194 nsew signal input
rlabel metal2 s 34608 0 34664 400 6 la_data_in[7]
port 195 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 la_data_in[8]
port 196 nsew signal input
rlabel metal2 s 38976 0 39032 400 6 la_data_in[9]
port 197 nsew signal input
rlabel metal3 s 39600 23184 40000 23240 6 la_data_out[0]
port 198 nsew signal output
rlabel metal3 s 39600 11760 40000 11816 6 la_data_out[10]
port 199 nsew signal output
rlabel metal3 s 0 26880 400 26936 6 la_data_out[11]
port 200 nsew signal output
rlabel metal2 s 28560 39600 28616 40000 6 la_data_out[12]
port 201 nsew signal output
rlabel metal3 s 39600 13776 40000 13832 6 la_data_out[13]
port 202 nsew signal output
rlabel metal3 s 39600 14784 40000 14840 6 la_data_out[14]
port 203 nsew signal output
rlabel metal2 s 19824 39600 19880 40000 6 la_data_out[15]
port 204 nsew signal output
rlabel metal3 s 39600 27216 40000 27272 6 la_data_out[16]
port 205 nsew signal output
rlabel metal2 s 24864 0 24920 400 6 la_data_out[17]
port 206 nsew signal output
rlabel metal2 s 16128 0 16184 400 6 la_data_out[18]
port 207 nsew signal output
rlabel metal2 s 23856 0 23912 400 6 la_data_out[19]
port 208 nsew signal output
rlabel metal2 s 23856 39600 23912 40000 6 la_data_out[1]
port 209 nsew signal output
rlabel metal2 s 22512 39600 22568 40000 6 la_data_out[20]
port 210 nsew signal output
rlabel metal3 s 0 29904 400 29960 6 la_data_out[21]
port 211 nsew signal output
rlabel metal2 s 14784 39600 14840 40000 6 la_data_out[22]
port 212 nsew signal output
rlabel metal3 s 0 6384 400 6440 6 la_data_out[23]
port 213 nsew signal output
rlabel metal2 s 24528 0 24584 400 6 la_data_out[24]
port 214 nsew signal output
rlabel metal2 s 18816 0 18872 400 6 la_data_out[25]
port 215 nsew signal output
rlabel metal3 s 39600 11088 40000 11144 6 la_data_out[26]
port 216 nsew signal output
rlabel metal3 s 39600 17136 40000 17192 6 la_data_out[27]
port 217 nsew signal output
rlabel metal3 s 0 21504 400 21560 6 la_data_out[28]
port 218 nsew signal output
rlabel metal2 s 21168 39600 21224 40000 6 la_data_out[29]
port 219 nsew signal output
rlabel metal3 s 0 28224 400 28280 6 la_data_out[2]
port 220 nsew signal output
rlabel metal3 s 0 17472 400 17528 6 la_data_out[30]
port 221 nsew signal output
rlabel metal2 s 19488 0 19544 400 6 la_data_out[31]
port 222 nsew signal output
rlabel metal2 s 24192 0 24248 400 6 la_data_out[32]
port 223 nsew signal output
rlabel metal2 s 17472 0 17528 400 6 la_data_out[33]
port 224 nsew signal output
rlabel metal2 s 16464 39600 16520 40000 6 la_data_out[34]
port 225 nsew signal output
rlabel metal2 s 18144 0 18200 400 6 la_data_out[35]
port 226 nsew signal output
rlabel metal3 s 39600 25872 40000 25928 6 la_data_out[36]
port 227 nsew signal output
rlabel metal2 s 22512 0 22568 400 6 la_data_out[37]
port 228 nsew signal output
rlabel metal2 s 27888 39600 27944 40000 6 la_data_out[38]
port 229 nsew signal output
rlabel metal2 s 18480 0 18536 400 6 la_data_out[39]
port 230 nsew signal output
rlabel metal2 s 20832 39600 20888 40000 6 la_data_out[3]
port 231 nsew signal output
rlabel metal3 s 39600 23856 40000 23912 6 la_data_out[40]
port 232 nsew signal output
rlabel metal3 s 0 32928 400 32984 6 la_data_out[41]
port 233 nsew signal output
rlabel metal2 s 17808 0 17864 400 6 la_data_out[42]
port 234 nsew signal output
rlabel metal3 s 39600 13440 40000 13496 6 la_data_out[43]
port 235 nsew signal output
rlabel metal3 s 39600 14112 40000 14168 6 la_data_out[44]
port 236 nsew signal output
rlabel metal2 s 12096 39600 12152 40000 6 la_data_out[45]
port 237 nsew signal output
rlabel metal2 s 26208 39600 26264 40000 6 la_data_out[46]
port 238 nsew signal output
rlabel metal3 s 39600 20832 40000 20888 6 la_data_out[47]
port 239 nsew signal output
rlabel metal2 s 22848 0 22904 400 6 la_data_out[48]
port 240 nsew signal output
rlabel metal2 s 23520 0 23576 400 6 la_data_out[49]
port 241 nsew signal output
rlabel metal3 s 39600 25200 40000 25256 6 la_data_out[4]
port 242 nsew signal output
rlabel metal2 s 17136 0 17192 400 6 la_data_out[50]
port 243 nsew signal output
rlabel metal2 s 13104 39600 13160 40000 6 la_data_out[51]
port 244 nsew signal output
rlabel metal2 s 22176 39600 22232 40000 6 la_data_out[52]
port 245 nsew signal output
rlabel metal3 s 0 13440 400 13496 6 la_data_out[53]
port 246 nsew signal output
rlabel metal3 s 39600 22512 40000 22568 6 la_data_out[54]
port 247 nsew signal output
rlabel metal2 s 18816 39600 18872 40000 6 la_data_out[55]
port 248 nsew signal output
rlabel metal3 s 0 28560 400 28616 6 la_data_out[56]
port 249 nsew signal output
rlabel metal3 s 0 32592 400 32648 6 la_data_out[57]
port 250 nsew signal output
rlabel metal2 s 21840 39600 21896 40000 6 la_data_out[58]
port 251 nsew signal output
rlabel metal3 s 39600 21168 40000 21224 6 la_data_out[59]
port 252 nsew signal output
rlabel metal3 s 0 7728 400 7784 6 la_data_out[5]
port 253 nsew signal output
rlabel metal3 s 0 7056 400 7112 6 la_data_out[60]
port 254 nsew signal output
rlabel metal2 s 28896 39600 28952 40000 6 la_data_out[61]
port 255 nsew signal output
rlabel metal3 s 39600 14448 40000 14504 6 la_data_out[62]
port 256 nsew signal output
rlabel metal2 s 17472 39600 17528 40000 6 la_data_out[63]
port 257 nsew signal output
rlabel metal3 s 39600 15792 40000 15848 6 la_data_out[6]
port 258 nsew signal output
rlabel metal3 s 0 16800 400 16856 6 la_data_out[7]
port 259 nsew signal output
rlabel metal3 s 39600 24192 40000 24248 6 la_data_out[8]
port 260 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 la_data_out[9]
port 261 nsew signal output
rlabel metal3 s 39600 1680 40000 1736 6 la_oenb[0]
port 262 nsew signal input
rlabel metal3 s 39600 36960 40000 37016 6 la_oenb[10]
port 263 nsew signal input
rlabel metal3 s 39600 30576 40000 30632 6 la_oenb[11]
port 264 nsew signal input
rlabel metal3 s 39600 8064 40000 8120 6 la_oenb[12]
port 265 nsew signal input
rlabel metal3 s 39600 4704 40000 4760 6 la_oenb[13]
port 266 nsew signal input
rlabel metal3 s 39600 31584 40000 31640 6 la_oenb[14]
port 267 nsew signal input
rlabel metal3 s 39600 8736 40000 8792 6 la_oenb[15]
port 268 nsew signal input
rlabel metal3 s 39600 5040 40000 5096 6 la_oenb[16]
port 269 nsew signal input
rlabel metal3 s 39600 34608 40000 34664 6 la_oenb[17]
port 270 nsew signal input
rlabel metal3 s 39600 6048 40000 6104 6 la_oenb[18]
port 271 nsew signal input
rlabel metal3 s 39600 4032 40000 4088 6 la_oenb[19]
port 272 nsew signal input
rlabel metal3 s 39600 3360 40000 3416 6 la_oenb[1]
port 273 nsew signal input
rlabel metal3 s 39600 38976 40000 39032 6 la_oenb[20]
port 274 nsew signal input
rlabel metal3 s 39600 7392 40000 7448 6 la_oenb[21]
port 275 nsew signal input
rlabel metal3 s 39600 5712 40000 5768 6 la_oenb[22]
port 276 nsew signal input
rlabel metal3 s 39600 3696 40000 3752 6 la_oenb[23]
port 277 nsew signal input
rlabel metal3 s 39600 672 40000 728 6 la_oenb[24]
port 278 nsew signal input
rlabel metal3 s 39600 37632 40000 37688 6 la_oenb[25]
port 279 nsew signal input
rlabel metal3 s 39600 0 40000 56 6 la_oenb[26]
port 280 nsew signal input
rlabel metal3 s 39600 39648 40000 39704 6 la_oenb[27]
port 281 nsew signal input
rlabel metal3 s 39600 9072 40000 9128 6 la_oenb[28]
port 282 nsew signal input
rlabel metal3 s 39600 2688 40000 2744 6 la_oenb[29]
port 283 nsew signal input
rlabel metal3 s 39600 36624 40000 36680 6 la_oenb[2]
port 284 nsew signal input
rlabel metal3 s 39600 9744 40000 9800 6 la_oenb[30]
port 285 nsew signal input
rlabel metal3 s 39600 37968 40000 38024 6 la_oenb[31]
port 286 nsew signal input
rlabel metal3 s 39600 1008 40000 1064 6 la_oenb[32]
port 287 nsew signal input
rlabel metal3 s 39600 9408 40000 9464 6 la_oenb[33]
port 288 nsew signal input
rlabel metal3 s 39600 3024 40000 3080 6 la_oenb[34]
port 289 nsew signal input
rlabel metal3 s 39600 29904 40000 29960 6 la_oenb[35]
port 290 nsew signal input
rlabel metal3 s 39600 38640 40000 38696 6 la_oenb[36]
port 291 nsew signal input
rlabel metal3 s 39600 38304 40000 38360 6 la_oenb[37]
port 292 nsew signal input
rlabel metal3 s 39600 36288 40000 36344 6 la_oenb[38]
port 293 nsew signal input
rlabel metal3 s 39600 1344 40000 1400 6 la_oenb[39]
port 294 nsew signal input
rlabel metal3 s 39600 32928 40000 32984 6 la_oenb[3]
port 295 nsew signal input
rlabel metal3 s 39600 35952 40000 36008 6 la_oenb[40]
port 296 nsew signal input
rlabel metal3 s 39600 33264 40000 33320 6 la_oenb[41]
port 297 nsew signal input
rlabel metal3 s 39600 7728 40000 7784 6 la_oenb[42]
port 298 nsew signal input
rlabel metal3 s 39600 30912 40000 30968 6 la_oenb[43]
port 299 nsew signal input
rlabel metal3 s 39600 33936 40000 33992 6 la_oenb[44]
port 300 nsew signal input
rlabel metal3 s 39600 39312 40000 39368 6 la_oenb[45]
port 301 nsew signal input
rlabel metal3 s 39600 2016 40000 2072 6 la_oenb[46]
port 302 nsew signal input
rlabel metal3 s 39600 31920 40000 31976 6 la_oenb[47]
port 303 nsew signal input
rlabel metal3 s 39600 32256 40000 32312 6 la_oenb[48]
port 304 nsew signal input
rlabel metal3 s 39600 5376 40000 5432 6 la_oenb[49]
port 305 nsew signal input
rlabel metal3 s 39600 30240 40000 30296 6 la_oenb[4]
port 306 nsew signal input
rlabel metal3 s 39600 35280 40000 35336 6 la_oenb[50]
port 307 nsew signal input
rlabel metal3 s 39600 2352 40000 2408 6 la_oenb[51]
port 308 nsew signal input
rlabel metal3 s 39600 8400 40000 8456 6 la_oenb[52]
port 309 nsew signal input
rlabel metal3 s 39600 34944 40000 35000 6 la_oenb[53]
port 310 nsew signal input
rlabel metal3 s 39600 31248 40000 31304 6 la_oenb[54]
port 311 nsew signal input
rlabel metal3 s 39600 37296 40000 37352 6 la_oenb[55]
port 312 nsew signal input
rlabel metal3 s 39600 6384 40000 6440 6 la_oenb[56]
port 313 nsew signal input
rlabel metal3 s 39600 7056 40000 7112 6 la_oenb[57]
port 314 nsew signal input
rlabel metal3 s 39600 29568 40000 29624 6 la_oenb[58]
port 315 nsew signal input
rlabel metal3 s 39600 6720 40000 6776 6 la_oenb[59]
port 316 nsew signal input
rlabel metal3 s 39600 34272 40000 34328 6 la_oenb[5]
port 317 nsew signal input
rlabel metal3 s 39600 4368 40000 4424 6 la_oenb[60]
port 318 nsew signal input
rlabel metal3 s 39600 35616 40000 35672 6 la_oenb[61]
port 319 nsew signal input
rlabel metal3 s 39600 32592 40000 32648 6 la_oenb[62]
port 320 nsew signal input
rlabel metal3 s 39600 336 40000 392 6 la_oenb[63]
port 321 nsew signal input
rlabel metal3 s 39600 33600 40000 33656 6 la_oenb[6]
port 322 nsew signal input
rlabel metal2 s 36624 39600 36680 40000 6 la_oenb[7]
port 323 nsew signal input
rlabel metal2 s 36960 39600 37016 40000 6 la_oenb[8]
port 324 nsew signal input
rlabel metal2 s 5040 39600 5096 40000 6 la_oenb[9]
port 325 nsew signal input
rlabel metal3 s 0 8736 400 8792 6 out[0]
port 326 nsew signal input
rlabel metal2 s 21504 39600 21560 40000 6 out[10]
port 327 nsew signal input
rlabel metal3 s 0 26544 400 26600 6 out[11]
port 328 nsew signal input
rlabel metal3 s 0 30240 400 30296 6 out[1]
port 329 nsew signal input
rlabel metal2 s 26880 39600 26936 40000 6 out[2]
port 330 nsew signal input
rlabel metal3 s 0 15792 400 15848 6 out[3]
port 331 nsew signal input
rlabel metal2 s 28224 39600 28280 40000 6 out[4]
port 332 nsew signal input
rlabel metal2 s 25200 39600 25256 40000 6 out[5]
port 333 nsew signal input
rlabel metal3 s 0 9744 400 9800 6 out[6]
port 334 nsew signal input
rlabel metal2 s 11760 39600 11816 40000 6 out[7]
port 335 nsew signal input
rlabel metal3 s 0 18480 400 18536 6 out[8]
port 336 nsew signal input
rlabel metal3 s 0 19152 400 19208 6 out[9]
port 337 nsew signal input
rlabel metal3 s 0 10752 400 10808 6 rst_n
port 338 nsew signal output
rlabel metal2 s 16800 39600 16856 40000 6 sel[0]
port 339 nsew signal output
rlabel metal2 s 25536 39600 25592 40000 6 sel[1]
port 340 nsew signal output
rlabel metal3 s 0 14112 400 14168 6 sel[2]
port 341 nsew signal output
rlabel metal2 s 32256 39600 32312 40000 6 user_clock2
port 342 nsew signal input
rlabel metal3 s 0 12432 400 12488 6 user_irq[0]
port 343 nsew signal output
rlabel metal3 s 0 33264 400 33320 6 user_irq[1]
port 344 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 user_irq[2]
port 345 nsew signal output
rlabel metal4 s 2224 1538 2384 38446 6 vdd
port 346 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 38446 6 vdd
port 346 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 38446 6 vdd
port 346 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 38446 6 vss
port 347 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 38446 6 vss
port 347 nsew ground bidirectional
rlabel metal2 s 23520 39600 23576 40000 6 wb_clk_i
port 348 nsew signal input
rlabel metal3 s 0 11088 400 11144 6 wb_rst_i
port 349 nsew signal input
rlabel metal2 s 18144 39600 18200 40000 6 wbs_ack_o
port 350 nsew signal output
rlabel metal2 s 36288 39600 36344 40000 6 wbs_adr_i[0]
port 351 nsew signal input
rlabel metal2 s 7392 39600 7448 40000 6 wbs_adr_i[10]
port 352 nsew signal input
rlabel metal2 s 8400 39600 8456 40000 6 wbs_adr_i[11]
port 353 nsew signal input
rlabel metal2 s 4368 39600 4424 40000 6 wbs_adr_i[12]
port 354 nsew signal input
rlabel metal2 s 33936 39600 33992 40000 6 wbs_adr_i[13]
port 355 nsew signal input
rlabel metal2 s 6384 39600 6440 40000 6 wbs_adr_i[14]
port 356 nsew signal input
rlabel metal2 s 29568 39600 29624 40000 6 wbs_adr_i[15]
port 357 nsew signal input
rlabel metal2 s 30912 39600 30968 40000 6 wbs_adr_i[16]
port 358 nsew signal input
rlabel metal2 s 39648 39600 39704 40000 6 wbs_adr_i[17]
port 359 nsew signal input
rlabel metal2 s 672 39600 728 40000 6 wbs_adr_i[18]
port 360 nsew signal input
rlabel metal2 s 38304 39600 38360 40000 6 wbs_adr_i[19]
port 361 nsew signal input
rlabel metal2 s 30240 39600 30296 40000 6 wbs_adr_i[1]
port 362 nsew signal input
rlabel metal2 s 31920 39600 31976 40000 6 wbs_adr_i[20]
port 363 nsew signal input
rlabel metal2 s 32592 39600 32648 40000 6 wbs_adr_i[21]
port 364 nsew signal input
rlabel metal2 s 33264 39600 33320 40000 6 wbs_adr_i[22]
port 365 nsew signal input
rlabel metal2 s 32928 39600 32984 40000 6 wbs_adr_i[23]
port 366 nsew signal input
rlabel metal2 s 9072 39600 9128 40000 6 wbs_adr_i[24]
port 367 nsew signal input
rlabel metal2 s 39312 39600 39368 40000 6 wbs_adr_i[25]
port 368 nsew signal input
rlabel metal2 s 29904 39600 29960 40000 6 wbs_adr_i[26]
port 369 nsew signal input
rlabel metal2 s 31584 39600 31640 40000 6 wbs_adr_i[27]
port 370 nsew signal input
rlabel metal2 s 31248 39600 31304 40000 6 wbs_adr_i[28]
port 371 nsew signal input
rlabel metal2 s 37296 39600 37352 40000 6 wbs_adr_i[29]
port 372 nsew signal input
rlabel metal2 s 30576 39600 30632 40000 6 wbs_adr_i[2]
port 373 nsew signal input
rlabel metal2 s 10752 39600 10808 40000 6 wbs_adr_i[30]
port 374 nsew signal input
rlabel metal2 s 37632 39600 37688 40000 6 wbs_adr_i[31]
port 375 nsew signal input
rlabel metal2 s 33600 39600 33656 40000 6 wbs_adr_i[3]
port 376 nsew signal input
rlabel metal2 s 9408 39600 9464 40000 6 wbs_adr_i[4]
port 377 nsew signal input
rlabel metal2 s 38976 39600 39032 40000 6 wbs_adr_i[5]
port 378 nsew signal input
rlabel metal2 s 38640 39600 38696 40000 6 wbs_adr_i[6]
port 379 nsew signal input
rlabel metal2 s 35952 39600 36008 40000 6 wbs_adr_i[7]
port 380 nsew signal input
rlabel metal2 s 2352 39600 2408 40000 6 wbs_adr_i[8]
port 381 nsew signal input
rlabel metal2 s 35280 39600 35336 40000 6 wbs_adr_i[9]
port 382 nsew signal input
rlabel metal2 s 1680 39600 1736 40000 6 wbs_cyc_i
port 383 nsew signal input
rlabel metal2 s 10080 39600 10136 40000 6 wbs_dat_i[0]
port 384 nsew signal input
rlabel metal2 s 1008 39600 1064 40000 6 wbs_dat_i[10]
port 385 nsew signal input
rlabel metal2 s 336 39600 392 40000 6 wbs_dat_i[11]
port 386 nsew signal input
rlabel metal2 s 34272 39600 34328 40000 6 wbs_dat_i[12]
port 387 nsew signal input
rlabel metal2 s 3696 39600 3752 40000 6 wbs_dat_i[13]
port 388 nsew signal input
rlabel metal2 s 1344 39600 1400 40000 6 wbs_dat_i[14]
port 389 nsew signal input
rlabel metal2 s 5376 39600 5432 40000 6 wbs_dat_i[15]
port 390 nsew signal input
rlabel metal2 s 2016 39600 2072 40000 6 wbs_dat_i[16]
port 391 nsew signal input
rlabel metal2 s 8736 39600 8792 40000 6 wbs_dat_i[17]
port 392 nsew signal input
rlabel metal2 s 4032 39600 4088 40000 6 wbs_dat_i[18]
port 393 nsew signal input
rlabel metal2 s 7056 39600 7112 40000 6 wbs_dat_i[19]
port 394 nsew signal input
rlabel metal2 s 6720 39600 6776 40000 6 wbs_dat_i[1]
port 395 nsew signal input
rlabel metal2 s 4704 39600 4760 40000 6 wbs_dat_i[20]
port 396 nsew signal input
rlabel metal2 s 5712 39600 5768 40000 6 wbs_dat_i[21]
port 397 nsew signal input
rlabel metal2 s 0 39600 56 40000 6 wbs_dat_i[22]
port 398 nsew signal input
rlabel metal2 s 37968 39600 38024 40000 6 wbs_dat_i[23]
port 399 nsew signal input
rlabel metal2 s 8064 39600 8120 40000 6 wbs_dat_i[24]
port 400 nsew signal input
rlabel metal2 s 7728 39600 7784 40000 6 wbs_dat_i[25]
port 401 nsew signal input
rlabel metal2 s 3024 39600 3080 40000 6 wbs_dat_i[26]
port 402 nsew signal input
rlabel metal2 s 2688 39600 2744 40000 6 wbs_dat_i[27]
port 403 nsew signal input
rlabel metal2 s 35616 39600 35672 40000 6 wbs_dat_i[28]
port 404 nsew signal input
rlabel metal2 s 6048 39600 6104 40000 6 wbs_dat_i[29]
port 405 nsew signal input
rlabel metal2 s 3360 39600 3416 40000 6 wbs_dat_i[2]
port 406 nsew signal input
rlabel metal2 s 10416 39600 10472 40000 6 wbs_dat_i[30]
port 407 nsew signal input
rlabel metal2 s 9744 39600 9800 40000 6 wbs_dat_i[31]
port 408 nsew signal input
rlabel metal2 s 34608 39600 34664 40000 6 wbs_dat_i[3]
port 409 nsew signal input
rlabel metal2 s 34944 39600 35000 40000 6 wbs_dat_i[4]
port 410 nsew signal input
rlabel metal3 s 0 39648 400 39704 6 wbs_dat_i[5]
port 411 nsew signal input
rlabel metal3 s 0 39312 400 39368 6 wbs_dat_i[6]
port 412 nsew signal input
rlabel metal3 s 0 38976 400 39032 6 wbs_dat_i[7]
port 413 nsew signal input
rlabel metal3 s 0 38640 400 38696 6 wbs_dat_i[8]
port 414 nsew signal input
rlabel metal3 s 0 38304 400 38360 6 wbs_dat_i[9]
port 415 nsew signal input
rlabel metal3 s 0 27552 400 27608 6 wbs_dat_o[0]
port 416 nsew signal output
rlabel metal3 s 0 28896 400 28952 6 wbs_dat_o[10]
port 417 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 wbs_dat_o[11]
port 418 nsew signal output
rlabel metal3 s 0 29232 400 29288 6 wbs_dat_o[12]
port 419 nsew signal output
rlabel metal3 s 0 13776 400 13832 6 wbs_dat_o[13]
port 420 nsew signal output
rlabel metal3 s 0 9408 400 9464 6 wbs_dat_o[14]
port 421 nsew signal output
rlabel metal3 s 0 25872 400 25928 6 wbs_dat_o[15]
port 422 nsew signal output
rlabel metal3 s 0 13104 400 13160 6 wbs_dat_o[16]
port 423 nsew signal output
rlabel metal3 s 0 7392 400 7448 6 wbs_dat_o[17]
port 424 nsew signal output
rlabel metal3 s 0 29568 400 29624 6 wbs_dat_o[18]
port 425 nsew signal output
rlabel metal3 s 0 18816 400 18872 6 wbs_dat_o[19]
port 426 nsew signal output
rlabel metal3 s 0 25536 400 25592 6 wbs_dat_o[1]
port 427 nsew signal output
rlabel metal3 s 0 25200 400 25256 6 wbs_dat_o[20]
port 428 nsew signal output
rlabel metal3 s 0 31584 400 31640 6 wbs_dat_o[21]
port 429 nsew signal output
rlabel metal3 s 0 10080 400 10136 6 wbs_dat_o[22]
port 430 nsew signal output
rlabel metal3 s 0 23856 400 23912 6 wbs_dat_o[23]
port 431 nsew signal output
rlabel metal3 s 0 24192 400 24248 6 wbs_dat_o[24]
port 432 nsew signal output
rlabel metal3 s 0 9072 400 9128 6 wbs_dat_o[25]
port 433 nsew signal output
rlabel metal3 s 0 26208 400 26264 6 wbs_dat_o[26]
port 434 nsew signal output
rlabel metal3 s 0 20496 400 20552 6 wbs_dat_o[27]
port 435 nsew signal output
rlabel metal3 s 0 23184 400 23240 6 wbs_dat_o[28]
port 436 nsew signal output
rlabel metal3 s 0 10416 400 10472 6 wbs_dat_o[29]
port 437 nsew signal output
rlabel metal3 s 0 21840 400 21896 6 wbs_dat_o[2]
port 438 nsew signal output
rlabel metal3 s 0 27888 400 27944 6 wbs_dat_o[30]
port 439 nsew signal output
rlabel metal3 s 0 22848 400 22904 6 wbs_dat_o[31]
port 440 nsew signal output
rlabel metal3 s 0 30576 400 30632 6 wbs_dat_o[3]
port 441 nsew signal output
rlabel metal3 s 0 23520 400 23576 6 wbs_dat_o[4]
port 442 nsew signal output
rlabel metal3 s 0 11760 400 11816 6 wbs_dat_o[5]
port 443 nsew signal output
rlabel metal3 s 0 24528 400 24584 6 wbs_dat_o[6]
port 444 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 wbs_dat_o[7]
port 445 nsew signal output
rlabel metal3 s 0 17808 400 17864 6 wbs_dat_o[8]
port 446 nsew signal output
rlabel metal3 s 0 24864 400 24920 6 wbs_dat_o[9]
port 447 nsew signal output
rlabel metal3 s 0 37968 400 38024 6 wbs_sel_i[0]
port 448 nsew signal input
rlabel metal3 s 0 37632 400 37688 6 wbs_sel_i[1]
port 449 nsew signal input
rlabel metal3 s 0 37296 400 37352 6 wbs_sel_i[2]
port 450 nsew signal input
rlabel metal3 s 0 36960 400 37016 6 wbs_sel_i[3]
port 451 nsew signal input
rlabel metal3 s 0 36624 400 36680 6 wbs_stb_i
port 452 nsew signal input
rlabel metal3 s 0 36288 400 36344 6 wbs_we_i
port 453 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 876954
string GDS_FILE /home/htamas/progs/gfmpw1-multi.v2/openlane/caravel_if/runs/23_12_13_05_14/results/signoff/caravel_if.magic.gds
string GDS_START 70906
<< end >>

