magic
tech gf180mcuD
magscale 1 10
timestamp 1702441052
<< metal1 >>
rect 43698 77198 43710 77250
rect 43762 77247 43774 77250
rect 44258 77247 44270 77250
rect 43762 77201 44270 77247
rect 43762 77198 43774 77201
rect 44258 77198 44270 77201
rect 44322 77198 44334 77250
rect 54450 77198 54462 77250
rect 54514 77247 54526 77250
rect 55234 77247 55246 77250
rect 54514 77201 55246 77247
rect 54514 77198 54526 77201
rect 55234 77198 55246 77201
rect 55298 77198 55310 77250
rect 27458 76974 27470 77026
rect 27522 77023 27534 77026
rect 28242 77023 28254 77026
rect 27522 76977 28254 77023
rect 27522 76974 27534 76977
rect 28242 76974 28254 76977
rect 28306 76974 28318 77026
rect 30818 76974 30830 77026
rect 30882 77023 30894 77026
rect 31714 77023 31726 77026
rect 30882 76977 31726 77023
rect 30882 76974 30894 76977
rect 31714 76974 31726 76977
rect 31778 76974 31790 77026
rect 53778 76974 53790 77026
rect 53842 77023 53854 77026
rect 54450 77023 54462 77026
rect 53842 76977 54462 77023
rect 53842 76974 53854 76977
rect 54450 76974 54462 76977
rect 54514 76974 54526 77026
rect 56466 76974 56478 77026
rect 56530 77023 56542 77026
rect 57026 77023 57038 77026
rect 56530 76977 57038 77023
rect 56530 76974 56542 76977
rect 57026 76974 57038 76977
rect 57090 76974 57102 77026
rect 1344 76858 78624 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 78624 76858
rect 1344 76772 78624 76806
rect 23102 76690 23154 76702
rect 23102 76626 23154 76638
rect 23998 76690 24050 76702
rect 23998 76626 24050 76638
rect 25230 76690 25282 76702
rect 25230 76626 25282 76638
rect 25790 76690 25842 76702
rect 25790 76626 25842 76638
rect 26462 76690 26514 76702
rect 26462 76626 26514 76638
rect 27022 76690 27074 76702
rect 27022 76626 27074 76638
rect 32510 76690 32562 76702
rect 32510 76626 32562 76638
rect 33182 76690 33234 76702
rect 33182 76626 33234 76638
rect 35198 76690 35250 76702
rect 35198 76626 35250 76638
rect 36654 76690 36706 76702
rect 36654 76626 36706 76638
rect 37886 76690 37938 76702
rect 37886 76626 37938 76638
rect 39902 76690 39954 76702
rect 39902 76626 39954 76638
rect 44270 76690 44322 76702
rect 44270 76626 44322 76638
rect 44718 76690 44770 76702
rect 44718 76626 44770 76638
rect 45278 76690 45330 76702
rect 45278 76626 45330 76638
rect 45950 76690 46002 76702
rect 45950 76626 46002 76638
rect 47966 76690 48018 76702
rect 47966 76626 48018 76638
rect 52222 76690 52274 76702
rect 52222 76626 52274 76638
rect 54462 76690 54514 76702
rect 54462 76626 54514 76638
rect 55358 76690 55410 76702
rect 55358 76626 55410 76638
rect 55694 76690 55746 76702
rect 55694 76626 55746 76638
rect 56142 76690 56194 76702
rect 56142 76626 56194 76638
rect 57038 76690 57090 76702
rect 57038 76626 57090 76638
rect 57374 76690 57426 76702
rect 57374 76626 57426 76638
rect 58046 76690 58098 76702
rect 58046 76626 58098 76638
rect 59838 76690 59890 76702
rect 59838 76626 59890 76638
rect 24894 76578 24946 76590
rect 24894 76514 24946 76526
rect 27470 76578 27522 76590
rect 27470 76514 27522 76526
rect 27806 76578 27858 76590
rect 27806 76514 27858 76526
rect 35982 76578 36034 76590
rect 35982 76514 36034 76526
rect 36318 76578 36370 76590
rect 36318 76514 36370 76526
rect 37214 76578 37266 76590
rect 37214 76514 37266 76526
rect 37550 76578 37602 76590
rect 37550 76514 37602 76526
rect 43598 76578 43650 76590
rect 43598 76514 43650 76526
rect 48638 76578 48690 76590
rect 48638 76514 48690 76526
rect 50318 76578 50370 76590
rect 54114 76526 54126 76578
rect 54178 76526 54190 76578
rect 55010 76526 55022 76578
rect 55074 76526 55086 76578
rect 56690 76526 56702 76578
rect 56754 76526 56766 76578
rect 50318 76514 50370 76526
rect 22878 76466 22930 76478
rect 22878 76402 22930 76414
rect 24558 76466 24610 76478
rect 47742 76466 47794 76478
rect 30818 76414 30830 76466
rect 30882 76414 30894 76466
rect 42578 76414 42590 76466
rect 42642 76414 42654 76466
rect 43810 76414 43822 76466
rect 43874 76414 43886 76466
rect 48850 76414 48862 76466
rect 48914 76414 48926 76466
rect 50530 76414 50542 76466
rect 50594 76414 50606 76466
rect 51202 76414 51214 76466
rect 51266 76414 51278 76466
rect 58818 76414 58830 76466
rect 58882 76414 58894 76466
rect 24558 76402 24610 76414
rect 47742 76402 47794 76414
rect 28590 76354 28642 76366
rect 28590 76290 28642 76302
rect 31614 76354 31666 76366
rect 31614 76290 31666 76302
rect 34302 76354 34354 76366
rect 34302 76290 34354 76302
rect 34526 76354 34578 76366
rect 34526 76290 34578 76302
rect 39118 76354 39170 76366
rect 46622 76354 46674 76366
rect 41010 76302 41022 76354
rect 41074 76302 41086 76354
rect 39118 76290 39170 76302
rect 46622 76290 46674 76302
rect 49310 76354 49362 76366
rect 49310 76290 49362 76302
rect 50094 76354 50146 76366
rect 50094 76290 50146 76302
rect 1344 76074 78624 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 78624 76074
rect 1344 75988 78624 76022
rect 22654 75906 22706 75918
rect 22654 75842 22706 75854
rect 30494 75906 30546 75918
rect 30494 75842 30546 75854
rect 34078 75906 34130 75918
rect 41582 75906 41634 75918
rect 38322 75854 38334 75906
rect 38386 75854 38398 75906
rect 34078 75842 34130 75854
rect 41582 75842 41634 75854
rect 28142 75794 28194 75806
rect 28142 75730 28194 75742
rect 28702 75794 28754 75806
rect 28702 75730 28754 75742
rect 37214 75794 37266 75806
rect 37214 75730 37266 75742
rect 44046 75794 44098 75806
rect 44046 75730 44098 75742
rect 50878 75794 50930 75806
rect 55694 75794 55746 75806
rect 53778 75742 53790 75794
rect 53842 75742 53854 75794
rect 50878 75730 50930 75742
rect 55694 75730 55746 75742
rect 56702 75794 56754 75806
rect 56702 75730 56754 75742
rect 25454 75682 25506 75694
rect 24994 75630 25006 75682
rect 25058 75630 25070 75682
rect 25454 75618 25506 75630
rect 29150 75682 29202 75694
rect 29150 75618 29202 75630
rect 31726 75682 31778 75694
rect 51662 75682 51714 75694
rect 58494 75682 58546 75694
rect 36418 75630 36430 75682
rect 36482 75630 36494 75682
rect 39778 75630 39790 75682
rect 39842 75630 39854 75682
rect 40562 75630 40574 75682
rect 40626 75630 40638 75682
rect 52658 75630 52670 75682
rect 52722 75630 52734 75682
rect 31726 75618 31778 75630
rect 51662 75618 51714 75630
rect 58494 75618 58546 75630
rect 29822 75570 29874 75582
rect 29822 75506 29874 75518
rect 31166 75570 31218 75582
rect 31166 75506 31218 75518
rect 43486 75570 43538 75582
rect 43486 75506 43538 75518
rect 52110 75570 52162 75582
rect 52110 75506 52162 75518
rect 56030 75570 56082 75582
rect 56030 75506 56082 75518
rect 29486 75458 29538 75470
rect 29486 75394 29538 75406
rect 1344 75290 78624 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 78624 75290
rect 1344 75204 78624 75238
rect 41918 75122 41970 75134
rect 41918 75058 41970 75070
rect 52334 75122 52386 75134
rect 52334 75058 52386 75070
rect 54350 75122 54402 75134
rect 54350 75058 54402 75070
rect 51314 74846 51326 74898
rect 51378 74846 51390 74898
rect 36654 74786 36706 74798
rect 36654 74722 36706 74734
rect 40350 74786 40402 74798
rect 40350 74722 40402 74734
rect 41022 74786 41074 74798
rect 41022 74722 41074 74734
rect 43262 74786 43314 74798
rect 43262 74722 43314 74734
rect 51102 74786 51154 74798
rect 51102 74722 51154 74734
rect 1344 74506 78624 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 78624 74506
rect 1344 74420 78624 74454
rect 1344 73722 78624 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 78624 73722
rect 1344 73636 78624 73670
rect 1344 72938 78624 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 78624 72938
rect 1344 72852 78624 72886
rect 1344 72154 78624 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 78624 72154
rect 1344 72068 78624 72102
rect 1344 71370 78624 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 78624 71370
rect 1344 71284 78624 71318
rect 1344 70586 78624 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 78624 70586
rect 1344 70500 78624 70534
rect 1344 69802 78624 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 78624 69802
rect 1344 69716 78624 69750
rect 1344 69018 78624 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 78624 69018
rect 1344 68932 78624 68966
rect 1344 68234 78624 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 78624 68234
rect 1344 68148 78624 68182
rect 1934 67954 1986 67966
rect 1934 67890 1986 67902
rect 4734 67842 4786 67854
rect 4274 67790 4286 67842
rect 4338 67790 4350 67842
rect 4734 67778 4786 67790
rect 1344 67450 78624 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 78624 67450
rect 1344 67364 78624 67398
rect 1710 67170 1762 67182
rect 1710 67106 1762 67118
rect 1344 66666 78624 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 78624 66666
rect 1344 66580 78624 66614
rect 1710 66050 1762 66062
rect 1710 65986 1762 65998
rect 1344 65882 78624 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 78624 65882
rect 1344 65796 78624 65830
rect 1710 65602 1762 65614
rect 1710 65538 1762 65550
rect 1344 65098 78624 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 78624 65098
rect 1344 65012 78624 65046
rect 2382 64818 2434 64830
rect 2382 64754 2434 64766
rect 1710 64594 1762 64606
rect 1710 64530 1762 64542
rect 2942 64594 2994 64606
rect 2942 64530 2994 64542
rect 2034 64430 2046 64482
rect 2098 64430 2110 64482
rect 1344 64314 78624 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 78624 64314
rect 1344 64228 78624 64262
rect 1710 64034 1762 64046
rect 1710 63970 1762 63982
rect 1344 63530 78624 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 78624 63530
rect 1344 63444 78624 63478
rect 1710 62914 1762 62926
rect 1710 62850 1762 62862
rect 1344 62746 78624 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 78624 62746
rect 1344 62660 78624 62694
rect 1710 62466 1762 62478
rect 1710 62402 1762 62414
rect 1344 61962 78624 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 78624 61962
rect 1344 61876 78624 61910
rect 1710 61346 1762 61358
rect 1710 61282 1762 61294
rect 1344 61178 78624 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 78624 61178
rect 1344 61092 78624 61126
rect 2034 60846 2046 60898
rect 2098 60846 2110 60898
rect 1710 60786 1762 60798
rect 1710 60722 1762 60734
rect 2494 60674 2546 60686
rect 2494 60610 2546 60622
rect 1344 60394 78624 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 78624 60394
rect 1344 60308 78624 60342
rect 2158 59890 2210 59902
rect 2158 59826 2210 59838
rect 1710 59778 1762 59790
rect 1710 59714 1762 59726
rect 1344 59610 78624 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 78624 59610
rect 1344 59524 78624 59558
rect 1710 59330 1762 59342
rect 78194 59278 78206 59330
rect 78258 59278 78270 59330
rect 1710 59266 1762 59278
rect 77970 59166 77982 59218
rect 78034 59166 78046 59218
rect 77534 59106 77586 59118
rect 77534 59042 77586 59054
rect 1344 58826 78624 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 78624 58826
rect 1344 58740 78624 58774
rect 78206 58546 78258 58558
rect 78206 58482 78258 58494
rect 1710 58210 1762 58222
rect 1710 58146 1762 58158
rect 1344 58042 78624 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 78624 58042
rect 1344 57956 78624 57990
rect 1710 57762 1762 57774
rect 1710 57698 1762 57710
rect 75618 57598 75630 57650
rect 75682 57598 75694 57650
rect 75406 57538 75458 57550
rect 77858 57486 77870 57538
rect 77922 57486 77934 57538
rect 75406 57474 75458 57486
rect 1344 57258 78624 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 78624 57258
rect 1344 57172 78624 57206
rect 1710 56642 1762 56654
rect 1710 56578 1762 56590
rect 77646 56642 77698 56654
rect 78206 56642 78258 56654
rect 77858 56590 77870 56642
rect 77922 56590 77934 56642
rect 77646 56578 77698 56590
rect 78206 56578 78258 56590
rect 1344 56474 78624 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 78624 56474
rect 1344 56388 78624 56422
rect 1710 56194 1762 56206
rect 1710 56130 1762 56142
rect 78206 56194 78258 56206
rect 78206 56130 78258 56142
rect 1344 55690 78624 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 78624 55690
rect 1344 55604 78624 55638
rect 1710 55410 1762 55422
rect 1710 55346 1762 55358
rect 2158 55186 2210 55198
rect 2158 55122 2210 55134
rect 77758 55186 77810 55198
rect 77758 55122 77810 55134
rect 78206 55074 78258 55086
rect 78206 55010 78258 55022
rect 1344 54906 78624 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 78624 54906
rect 1344 54820 78624 54854
rect 1710 54626 1762 54638
rect 1710 54562 1762 54574
rect 75618 54462 75630 54514
rect 75682 54462 75694 54514
rect 75406 54402 75458 54414
rect 77858 54350 77870 54402
rect 77922 54350 77934 54402
rect 75406 54338 75458 54350
rect 1344 54122 78624 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 78624 54122
rect 1344 54036 78624 54070
rect 78206 53842 78258 53854
rect 78206 53778 78258 53790
rect 1810 53678 1822 53730
rect 1874 53678 1886 53730
rect 2046 53506 2098 53518
rect 2046 53442 2098 53454
rect 2494 53506 2546 53518
rect 2494 53442 2546 53454
rect 1344 53338 78624 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 78624 53338
rect 1344 53252 78624 53286
rect 1710 53058 1762 53070
rect 1710 52994 1762 53006
rect 78206 52722 78258 52734
rect 78206 52658 78258 52670
rect 1344 52554 78624 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 78624 52554
rect 1344 52468 78624 52502
rect 1710 51938 1762 51950
rect 1710 51874 1762 51886
rect 78206 51938 78258 51950
rect 78206 51874 78258 51886
rect 1344 51770 78624 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 78624 51770
rect 1344 51684 78624 51718
rect 1710 51490 1762 51502
rect 1710 51426 1762 51438
rect 77870 51490 77922 51502
rect 77870 51426 77922 51438
rect 78206 51378 78258 51390
rect 78206 51314 78258 51326
rect 77646 51266 77698 51278
rect 77646 51202 77698 51214
rect 1344 50986 78624 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 78624 50986
rect 1344 50900 78624 50934
rect 1710 50370 1762 50382
rect 1710 50306 1762 50318
rect 2158 50370 2210 50382
rect 2158 50306 2210 50318
rect 77758 50370 77810 50382
rect 77758 50306 77810 50318
rect 78206 50370 78258 50382
rect 78206 50306 78258 50318
rect 1344 50202 78624 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 78624 50202
rect 1344 50116 78624 50150
rect 1710 49922 1762 49934
rect 1710 49858 1762 49870
rect 78206 49922 78258 49934
rect 78206 49858 78258 49870
rect 1344 49418 78624 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 78624 49418
rect 1344 49332 78624 49366
rect 1710 48802 1762 48814
rect 1710 48738 1762 48750
rect 78206 48802 78258 48814
rect 78206 48738 78258 48750
rect 1344 48634 78624 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 78624 48634
rect 1344 48548 78624 48582
rect 39566 48466 39618 48478
rect 39566 48402 39618 48414
rect 39790 48466 39842 48478
rect 39790 48402 39842 48414
rect 43822 48466 43874 48478
rect 43822 48402 43874 48414
rect 44382 48466 44434 48478
rect 44382 48402 44434 48414
rect 1710 48354 1762 48366
rect 1710 48290 1762 48302
rect 78206 48354 78258 48366
rect 78206 48290 78258 48302
rect 40226 48078 40238 48130
rect 40290 48078 40302 48130
rect 43362 48078 43374 48130
rect 43426 48078 43438 48130
rect 1344 47850 78624 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 78624 47850
rect 1344 47764 78624 47798
rect 36430 47570 36482 47582
rect 36430 47506 36482 47518
rect 1710 47234 1762 47246
rect 1710 47170 1762 47182
rect 35534 47234 35586 47246
rect 35534 47170 35586 47182
rect 35870 47234 35922 47246
rect 35870 47170 35922 47182
rect 78206 47234 78258 47246
rect 78206 47170 78258 47182
rect 1344 47066 78624 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 78624 47066
rect 1344 46980 78624 47014
rect 34750 46898 34802 46910
rect 34750 46834 34802 46846
rect 34974 46898 35026 46910
rect 34974 46834 35026 46846
rect 43374 46898 43426 46910
rect 43374 46834 43426 46846
rect 43934 46898 43986 46910
rect 43934 46834 43986 46846
rect 47182 46898 47234 46910
rect 47182 46834 47234 46846
rect 1710 46786 1762 46798
rect 46722 46734 46734 46786
rect 46786 46734 46798 46786
rect 1710 46722 1762 46734
rect 46498 46622 46510 46674
rect 46562 46622 46574 46674
rect 75618 46622 75630 46674
rect 75682 46622 75694 46674
rect 75406 46562 75458 46574
rect 35410 46510 35422 46562
rect 35474 46510 35486 46562
rect 42914 46510 42926 46562
rect 42978 46510 42990 46562
rect 77858 46510 77870 46562
rect 77922 46510 77934 46562
rect 75406 46498 75458 46510
rect 1344 46282 78624 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 78624 46282
rect 1344 46196 78624 46230
rect 2158 45778 2210 45790
rect 2158 45714 2210 45726
rect 77758 45778 77810 45790
rect 77758 45714 77810 45726
rect 1710 45666 1762 45678
rect 1710 45602 1762 45614
rect 78206 45666 78258 45678
rect 78206 45602 78258 45614
rect 1344 45498 78624 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 78624 45498
rect 1344 45412 78624 45446
rect 45614 45330 45666 45342
rect 45614 45266 45666 45278
rect 46174 45330 46226 45342
rect 46174 45266 46226 45278
rect 78206 45218 78258 45230
rect 78206 45154 78258 45166
rect 4846 45106 4898 45118
rect 4274 45054 4286 45106
rect 4338 45054 4350 45106
rect 4846 45042 4898 45054
rect 41470 45106 41522 45118
rect 41470 45042 41522 45054
rect 42030 45106 42082 45118
rect 42030 45042 42082 45054
rect 41010 44942 41022 44994
rect 41074 44942 41086 44994
rect 45154 44942 45166 44994
rect 45218 44942 45230 44994
rect 1934 44882 1986 44894
rect 1934 44818 1986 44830
rect 1344 44714 78624 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 78624 44714
rect 1344 44628 78624 44662
rect 34850 44382 34862 44434
rect 34914 44382 34926 44434
rect 42690 44382 42702 44434
rect 42754 44382 42766 44434
rect 44930 44382 44942 44434
rect 44994 44382 45006 44434
rect 36430 44322 36482 44334
rect 36430 44258 36482 44270
rect 34078 44210 34130 44222
rect 34078 44146 34130 44158
rect 34414 44210 34466 44222
rect 34414 44146 34466 44158
rect 43150 44210 43202 44222
rect 43150 44146 43202 44158
rect 43598 44210 43650 44222
rect 43598 44146 43650 44158
rect 1710 44098 1762 44110
rect 1710 44034 1762 44046
rect 35534 44098 35586 44110
rect 35534 44034 35586 44046
rect 35870 44098 35922 44110
rect 35870 44034 35922 44046
rect 45390 44098 45442 44110
rect 45390 44034 45442 44046
rect 45838 44098 45890 44110
rect 45838 44034 45890 44046
rect 78206 44098 78258 44110
rect 78206 44034 78258 44046
rect 1344 43930 78624 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 78624 43930
rect 1344 43844 78624 43878
rect 78206 43762 78258 43774
rect 78206 43698 78258 43710
rect 1710 43650 1762 43662
rect 1710 43586 1762 43598
rect 1344 43146 78624 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 78624 43146
rect 1344 43060 78624 43094
rect 45838 42754 45890 42766
rect 45838 42690 45890 42702
rect 1710 42530 1762 42542
rect 1710 42466 1762 42478
rect 46398 42530 46450 42542
rect 46398 42466 46450 42478
rect 46846 42530 46898 42542
rect 46846 42466 46898 42478
rect 78206 42530 78258 42542
rect 78206 42466 78258 42478
rect 1344 42362 78624 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 78624 42362
rect 1344 42276 78624 42310
rect 78206 42082 78258 42094
rect 78206 42018 78258 42030
rect 38110 41970 38162 41982
rect 4274 41918 4286 41970
rect 4338 41918 4350 41970
rect 38110 41906 38162 41918
rect 38334 41970 38386 41982
rect 38334 41906 38386 41918
rect 38894 41970 38946 41982
rect 38894 41906 38946 41918
rect 45390 41970 45442 41982
rect 45390 41906 45442 41918
rect 45950 41970 46002 41982
rect 45950 41906 46002 41918
rect 4846 41858 4898 41870
rect 44930 41806 44942 41858
rect 44994 41806 45006 41858
rect 4846 41794 4898 41806
rect 1934 41746 1986 41758
rect 1934 41682 1986 41694
rect 1344 41578 78624 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 78624 41578
rect 1344 41492 78624 41526
rect 34402 41246 34414 41298
rect 34466 41246 34478 41298
rect 1710 41074 1762 41086
rect 1710 41010 1762 41022
rect 78206 41074 78258 41086
rect 78206 41010 78258 41022
rect 2158 40962 2210 40974
rect 2158 40898 2210 40910
rect 33630 40962 33682 40974
rect 33630 40898 33682 40910
rect 33966 40962 34018 40974
rect 33966 40898 34018 40910
rect 77758 40962 77810 40974
rect 77758 40898 77810 40910
rect 1344 40794 78624 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 78624 40794
rect 1344 40708 78624 40742
rect 78206 40514 78258 40526
rect 78206 40450 78258 40462
rect 34414 40402 34466 40414
rect 34414 40338 34466 40350
rect 34638 40402 34690 40414
rect 34638 40338 34690 40350
rect 35198 40402 35250 40414
rect 35198 40338 35250 40350
rect 1710 40178 1762 40190
rect 1710 40114 1762 40126
rect 1344 40010 78624 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 78624 40010
rect 1344 39924 78624 39958
rect 78206 39730 78258 39742
rect 40338 39678 40350 39730
rect 40402 39678 40414 39730
rect 78206 39666 78258 39678
rect 41694 39618 41746 39630
rect 41694 39554 41746 39566
rect 44830 39618 44882 39630
rect 44830 39554 44882 39566
rect 1710 39394 1762 39406
rect 1710 39330 1762 39342
rect 40014 39394 40066 39406
rect 40014 39330 40066 39342
rect 40798 39394 40850 39406
rect 40798 39330 40850 39342
rect 41134 39394 41186 39406
rect 41134 39330 41186 39342
rect 45390 39394 45442 39406
rect 45390 39330 45442 39342
rect 45950 39394 46002 39406
rect 45950 39330 46002 39342
rect 1344 39226 78624 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 78624 39226
rect 1344 39140 78624 39174
rect 2046 38946 2098 38958
rect 2046 38882 2098 38894
rect 1710 38834 1762 38846
rect 1710 38770 1762 38782
rect 35310 38834 35362 38846
rect 35310 38770 35362 38782
rect 38334 38834 38386 38846
rect 38334 38770 38386 38782
rect 39230 38834 39282 38846
rect 39230 38770 39282 38782
rect 44046 38834 44098 38846
rect 44046 38770 44098 38782
rect 2494 38722 2546 38734
rect 2494 38658 2546 38670
rect 34974 38722 35026 38734
rect 34974 38658 35026 38670
rect 35870 38722 35922 38734
rect 35870 38658 35922 38670
rect 37998 38722 38050 38734
rect 39790 38722 39842 38734
rect 38770 38670 38782 38722
rect 38834 38670 38846 38722
rect 37998 38658 38050 38670
rect 39790 38658 39842 38670
rect 41022 38722 41074 38734
rect 41022 38658 41074 38670
rect 43710 38722 43762 38734
rect 43710 38658 43762 38670
rect 44606 38722 44658 38734
rect 44606 38658 44658 38670
rect 78206 38610 78258 38622
rect 78206 38546 78258 38558
rect 1344 38442 78624 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 78624 38442
rect 1344 38356 78624 38390
rect 33406 38050 33458 38062
rect 33406 37986 33458 37998
rect 1710 37826 1762 37838
rect 1710 37762 1762 37774
rect 32622 37826 32674 37838
rect 32622 37762 32674 37774
rect 32846 37826 32898 37838
rect 32846 37762 32898 37774
rect 38894 37826 38946 37838
rect 38894 37762 38946 37774
rect 78206 37826 78258 37838
rect 78206 37762 78258 37774
rect 1344 37658 78624 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 78624 37658
rect 1344 37572 78624 37606
rect 2046 37378 2098 37390
rect 2046 37314 2098 37326
rect 78206 37378 78258 37390
rect 78206 37314 78258 37326
rect 1710 37266 1762 37278
rect 1710 37202 1762 37214
rect 33854 37266 33906 37278
rect 33854 37202 33906 37214
rect 2494 37154 2546 37166
rect 2494 37090 2546 37102
rect 33518 37154 33570 37166
rect 33518 37090 33570 37102
rect 34414 37154 34466 37166
rect 34414 37090 34466 37102
rect 1344 36874 78624 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 78624 36874
rect 1344 36788 78624 36822
rect 77758 36594 77810 36606
rect 77758 36530 77810 36542
rect 34974 36482 35026 36494
rect 34974 36418 35026 36430
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 2046 36370 2098 36382
rect 2046 36306 2098 36318
rect 2942 36370 2994 36382
rect 2942 36306 2994 36318
rect 78206 36370 78258 36382
rect 78206 36306 78258 36318
rect 2382 36258 2434 36270
rect 2382 36194 2434 36206
rect 34190 36258 34242 36270
rect 34190 36194 34242 36206
rect 34414 36258 34466 36270
rect 34414 36194 34466 36206
rect 1344 36090 78624 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 78624 36090
rect 1344 36004 78624 36038
rect 1710 35810 1762 35822
rect 1710 35746 1762 35758
rect 40126 35698 40178 35710
rect 40126 35634 40178 35646
rect 43150 35698 43202 35710
rect 43150 35634 43202 35646
rect 44158 35698 44210 35710
rect 44158 35634 44210 35646
rect 33630 35586 33682 35598
rect 33630 35522 33682 35534
rect 33854 35586 33906 35598
rect 39566 35586 39618 35598
rect 34066 35534 34078 35586
rect 34130 35534 34142 35586
rect 33854 35522 33906 35534
rect 39566 35522 39618 35534
rect 41022 35586 41074 35598
rect 43586 35534 43598 35586
rect 43650 35534 43662 35586
rect 41022 35522 41074 35534
rect 78206 35474 78258 35486
rect 78206 35410 78258 35422
rect 1344 35306 78624 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 78624 35306
rect 1344 35220 78624 35254
rect 45266 34974 45278 35026
rect 45330 34974 45342 35026
rect 1810 34862 1822 34914
rect 1874 34862 1886 34914
rect 2046 34690 2098 34702
rect 2046 34626 2098 34638
rect 2494 34690 2546 34702
rect 2494 34626 2546 34638
rect 44382 34690 44434 34702
rect 44382 34626 44434 34638
rect 44830 34690 44882 34702
rect 44830 34626 44882 34638
rect 78206 34690 78258 34702
rect 78206 34626 78258 34638
rect 1344 34522 78624 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 78624 34522
rect 1344 34436 78624 34470
rect 1710 34242 1762 34254
rect 1710 34178 1762 34190
rect 77870 34242 77922 34254
rect 77870 34178 77922 34190
rect 34190 34130 34242 34142
rect 46622 34130 46674 34142
rect 34626 34078 34638 34130
rect 34690 34078 34702 34130
rect 34190 34066 34242 34078
rect 46622 34066 46674 34078
rect 78206 34130 78258 34142
rect 78206 34066 78258 34078
rect 35086 34018 35138 34030
rect 35086 33954 35138 33966
rect 46062 34018 46114 34030
rect 46062 33954 46114 33966
rect 47070 34018 47122 34030
rect 47070 33954 47122 33966
rect 77646 34018 77698 34030
rect 77646 33954 77698 33966
rect 1344 33738 78624 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 78624 33738
rect 1344 33652 78624 33686
rect 1710 33458 1762 33470
rect 1710 33394 1762 33406
rect 40462 33346 40514 33358
rect 40462 33282 40514 33294
rect 41022 33122 41074 33134
rect 41022 33058 41074 33070
rect 41582 33122 41634 33134
rect 41582 33058 41634 33070
rect 78206 33122 78258 33134
rect 78206 33058 78258 33070
rect 1344 32954 78624 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 78624 32954
rect 1344 32868 78624 32902
rect 2046 32674 2098 32686
rect 2046 32610 2098 32622
rect 78206 32674 78258 32686
rect 78206 32610 78258 32622
rect 1710 32562 1762 32574
rect 1710 32498 1762 32510
rect 44046 32562 44098 32574
rect 44046 32498 44098 32510
rect 44494 32562 44546 32574
rect 44494 32498 44546 32510
rect 2494 32450 2546 32462
rect 2494 32386 2546 32398
rect 43486 32450 43538 32462
rect 43486 32386 43538 32398
rect 1344 32170 78624 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 78624 32170
rect 1344 32084 78624 32118
rect 77758 32002 77810 32014
rect 77758 31938 77810 31950
rect 1934 31890 1986 31902
rect 1934 31826 1986 31838
rect 4846 31778 4898 31790
rect 4274 31726 4286 31778
rect 4338 31726 4350 31778
rect 4846 31714 4898 31726
rect 78206 31666 78258 31678
rect 78206 31602 78258 31614
rect 1344 31386 78624 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 78624 31386
rect 1344 31300 78624 31334
rect 2942 31218 2994 31230
rect 2942 31154 2994 31166
rect 1710 31106 1762 31118
rect 1710 31042 1762 31054
rect 2046 31106 2098 31118
rect 2046 31042 2098 31054
rect 75618 30942 75630 30994
rect 75682 30942 75694 30994
rect 75294 30882 75346 30894
rect 75294 30818 75346 30830
rect 2382 30770 2434 30782
rect 2382 30706 2434 30718
rect 77982 30770 78034 30782
rect 77982 30706 78034 30718
rect 1344 30602 78624 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 78624 30602
rect 1344 30516 78624 30550
rect 4274 30158 4286 30210
rect 4338 30158 4350 30210
rect 2482 30046 2494 30098
rect 2546 30046 2558 30098
rect 4846 29986 4898 29998
rect 4846 29922 4898 29934
rect 78206 29986 78258 29998
rect 78206 29922 78258 29934
rect 1344 29818 78624 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 78624 29818
rect 1344 29732 78624 29766
rect 78206 29538 78258 29550
rect 78206 29474 78258 29486
rect 1710 29202 1762 29214
rect 1710 29138 1762 29150
rect 1344 29034 78624 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 78624 29034
rect 1344 28948 78624 28982
rect 1934 28754 1986 28766
rect 1934 28690 1986 28702
rect 4846 28642 4898 28654
rect 4274 28590 4286 28642
rect 4338 28590 4350 28642
rect 4846 28578 4898 28590
rect 78206 28418 78258 28430
rect 78206 28354 78258 28366
rect 1344 28250 78624 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 78624 28250
rect 1344 28164 78624 28198
rect 1710 27970 1762 27982
rect 1710 27906 1762 27918
rect 78206 27970 78258 27982
rect 78206 27906 78258 27918
rect 1344 27466 78624 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 78624 27466
rect 1344 27380 78624 27414
rect 77198 27186 77250 27198
rect 77198 27122 77250 27134
rect 78206 26962 78258 26974
rect 77858 26910 77870 26962
rect 77922 26910 77934 26962
rect 78206 26898 78258 26910
rect 1710 26850 1762 26862
rect 1710 26786 1762 26798
rect 2158 26850 2210 26862
rect 2158 26786 2210 26798
rect 77534 26850 77586 26862
rect 77534 26786 77586 26798
rect 1344 26682 78624 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 78624 26682
rect 1344 26596 78624 26630
rect 1710 26402 1762 26414
rect 1710 26338 1762 26350
rect 75618 26238 75630 26290
rect 75682 26238 75694 26290
rect 75294 26178 75346 26190
rect 75294 26114 75346 26126
rect 77982 26066 78034 26078
rect 77982 26002 78034 26014
rect 1344 25898 78624 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 78624 25898
rect 1344 25812 78624 25846
rect 1710 25282 1762 25294
rect 1710 25218 1762 25230
rect 1344 25114 78624 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 78624 25114
rect 1344 25028 78624 25062
rect 1710 24834 1762 24846
rect 1710 24770 1762 24782
rect 75730 24670 75742 24722
rect 75794 24670 75806 24722
rect 75294 24610 75346 24622
rect 75294 24546 75346 24558
rect 77982 24610 78034 24622
rect 77982 24546 78034 24558
rect 1344 24330 78624 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 78624 24330
rect 1344 24244 78624 24278
rect 78206 23826 78258 23838
rect 78206 23762 78258 23774
rect 1710 23714 1762 23726
rect 1710 23650 1762 23662
rect 77758 23714 77810 23726
rect 77758 23650 77810 23662
rect 1344 23546 78624 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 78624 23546
rect 1344 23460 78624 23494
rect 1710 23266 1762 23278
rect 1710 23202 1762 23214
rect 75730 23102 75742 23154
rect 75794 23102 75806 23154
rect 75294 23042 75346 23054
rect 75294 22978 75346 22990
rect 77982 22930 78034 22942
rect 77982 22866 78034 22878
rect 1344 22762 78624 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 78624 22762
rect 1344 22676 78624 22710
rect 1934 22482 1986 22494
rect 1934 22418 1986 22430
rect 4846 22370 4898 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 4846 22306 4898 22318
rect 78206 22258 78258 22270
rect 78206 22194 78258 22206
rect 1344 21978 78624 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 78624 21978
rect 1344 21892 78624 21926
rect 1710 21810 1762 21822
rect 1710 21746 1762 21758
rect 2942 21810 2994 21822
rect 2942 21746 2994 21758
rect 2382 21698 2434 21710
rect 2034 21646 2046 21698
rect 2098 21646 2110 21698
rect 2382 21634 2434 21646
rect 75618 21534 75630 21586
rect 75682 21534 75694 21586
rect 75294 21474 75346 21486
rect 75294 21410 75346 21422
rect 77982 21474 78034 21486
rect 77982 21410 78034 21422
rect 1344 21194 78624 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 78624 21194
rect 1344 21108 78624 21142
rect 77646 20914 77698 20926
rect 77646 20850 77698 20862
rect 78206 20802 78258 20814
rect 78206 20738 78258 20750
rect 1710 20578 1762 20590
rect 77858 20526 77870 20578
rect 77922 20526 77934 20578
rect 1710 20514 1762 20526
rect 1344 20410 78624 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 78624 20410
rect 1344 20324 78624 20358
rect 2034 20078 2046 20130
rect 2098 20078 2110 20130
rect 1710 20018 1762 20030
rect 75618 19966 75630 20018
rect 75682 19966 75694 20018
rect 1710 19954 1762 19966
rect 2494 19906 2546 19918
rect 2494 19842 2546 19854
rect 75294 19906 75346 19918
rect 75294 19842 75346 19854
rect 77982 19906 78034 19918
rect 77982 19842 78034 19854
rect 1344 19626 78624 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 78624 19626
rect 1344 19540 78624 19574
rect 1710 19010 1762 19022
rect 1710 18946 1762 18958
rect 1344 18842 78624 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 78624 18842
rect 1344 18756 78624 18790
rect 1710 18562 1762 18574
rect 1710 18498 1762 18510
rect 1344 18058 78624 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 78624 18058
rect 1344 17972 78624 18006
rect 1934 17778 1986 17790
rect 1934 17714 1986 17726
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 4846 17442 4898 17454
rect 4846 17378 4898 17390
rect 1344 17274 78624 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 78624 17274
rect 1344 17188 78624 17222
rect 1710 17106 1762 17118
rect 1710 17042 1762 17054
rect 2942 17106 2994 17118
rect 2942 17042 2994 17054
rect 2382 16994 2434 17006
rect 2034 16942 2046 16994
rect 2098 16942 2110 16994
rect 2382 16930 2434 16942
rect 1344 16490 78624 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 78624 16490
rect 1344 16404 78624 16438
rect 1710 15874 1762 15886
rect 1710 15810 1762 15822
rect 1344 15706 78624 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 78624 15706
rect 1344 15620 78624 15654
rect 1710 15426 1762 15438
rect 1710 15362 1762 15374
rect 1344 14922 78624 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 78624 14922
rect 1344 14836 78624 14870
rect 1710 14306 1762 14318
rect 1710 14242 1762 14254
rect 1344 14138 78624 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 78624 14138
rect 1344 14052 78624 14086
rect 1710 13522 1762 13534
rect 1710 13458 1762 13470
rect 1344 13354 78624 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 78624 13354
rect 1344 13268 78624 13302
rect 1934 13074 1986 13086
rect 1934 13010 1986 13022
rect 4274 12910 4286 12962
rect 4338 12910 4350 12962
rect 4846 12738 4898 12750
rect 4846 12674 4898 12686
rect 1344 12570 78624 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 78624 12570
rect 1344 12484 78624 12518
rect 1710 12402 1762 12414
rect 1710 12338 1762 12350
rect 1344 11786 78624 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 78624 11786
rect 1344 11700 78624 11734
rect 1344 11002 78624 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 78624 11002
rect 1344 10916 78624 10950
rect 1344 10218 78624 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 78624 10218
rect 1344 10132 78624 10166
rect 1344 9434 78624 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 78624 9434
rect 1344 9348 78624 9382
rect 1344 8650 78624 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 78624 8650
rect 1344 8564 78624 8598
rect 1344 7866 78624 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 78624 7866
rect 1344 7780 78624 7814
rect 1344 7082 78624 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 78624 7082
rect 1344 6996 78624 7030
rect 1344 6298 78624 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 78624 6298
rect 1344 6212 78624 6246
rect 1344 5514 78624 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 78624 5514
rect 1344 5428 78624 5462
rect 43262 4898 43314 4910
rect 43262 4834 43314 4846
rect 1344 4730 78624 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 78624 4730
rect 1344 4644 78624 4678
rect 36878 4562 36930 4574
rect 36878 4498 36930 4510
rect 42478 4562 42530 4574
rect 42478 4498 42530 4510
rect 46174 4450 46226 4462
rect 46174 4386 46226 4398
rect 46622 4450 46674 4462
rect 46622 4386 46674 4398
rect 29586 4286 29598 4338
rect 29650 4286 29662 4338
rect 35970 4286 35982 4338
rect 36034 4286 36046 4338
rect 43362 4286 43374 4338
rect 43426 4286 43438 4338
rect 51986 4286 51998 4338
rect 52050 4286 52062 4338
rect 30158 4226 30210 4238
rect 30158 4162 30210 4174
rect 41134 4226 41186 4238
rect 41134 4162 41186 4174
rect 41694 4226 41746 4238
rect 41694 4162 41746 4174
rect 43038 4226 43090 4238
rect 43038 4162 43090 4174
rect 47182 4226 47234 4238
rect 47182 4162 47234 4174
rect 50878 4226 50930 4238
rect 50878 4162 50930 4174
rect 51662 4226 51714 4238
rect 51662 4162 51714 4174
rect 27358 4114 27410 4126
rect 27358 4050 27410 4062
rect 34078 4114 34130 4126
rect 44270 4114 44322 4126
rect 42802 4062 42814 4114
rect 42866 4111 42878 4114
rect 43026 4111 43038 4114
rect 42866 4065 43038 4111
rect 42866 4062 42878 4065
rect 43026 4062 43038 4065
rect 43090 4062 43102 4114
rect 34078 4050 34130 4062
rect 44270 4050 44322 4062
rect 53006 4114 53058 4126
rect 53006 4050 53058 4062
rect 1344 3946 78624 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 78624 3946
rect 1344 3860 78624 3894
rect 29150 3666 29202 3678
rect 29150 3602 29202 3614
rect 29822 3666 29874 3678
rect 29822 3602 29874 3614
rect 30494 3666 30546 3678
rect 30494 3602 30546 3614
rect 31614 3666 31666 3678
rect 31614 3602 31666 3614
rect 39902 3666 39954 3678
rect 39902 3602 39954 3614
rect 44606 3666 44658 3678
rect 44606 3602 44658 3614
rect 52222 3666 52274 3678
rect 52222 3602 52274 3614
rect 27246 3554 27298 3566
rect 27570 3502 27582 3554
rect 27634 3502 27646 3554
rect 42130 3502 42142 3554
rect 42194 3502 42206 3554
rect 42802 3502 42814 3554
rect 42866 3502 42878 3554
rect 43698 3502 43710 3554
rect 43762 3502 43774 3554
rect 46722 3502 46734 3554
rect 46786 3502 46798 3554
rect 51202 3502 51214 3554
rect 51266 3502 51278 3554
rect 27246 3490 27298 3502
rect 26798 3442 26850 3454
rect 28478 3442 28530 3454
rect 41246 3442 41298 3454
rect 27794 3390 27806 3442
rect 27858 3390 27870 3442
rect 28802 3390 28814 3442
rect 28866 3390 28878 3442
rect 26798 3378 26850 3390
rect 28478 3378 28530 3390
rect 41246 3378 41298 3390
rect 41582 3442 41634 3454
rect 41582 3378 41634 3390
rect 41918 3442 41970 3454
rect 41918 3378 41970 3390
rect 43038 3442 43090 3454
rect 43038 3378 43090 3390
rect 46510 3442 46562 3454
rect 46510 3378 46562 3390
rect 31054 3330 31106 3342
rect 31054 3266 31106 3278
rect 32510 3330 32562 3342
rect 32510 3266 32562 3278
rect 33182 3330 33234 3342
rect 33182 3266 33234 3278
rect 34526 3330 34578 3342
rect 34526 3266 34578 3278
rect 35198 3330 35250 3342
rect 35198 3266 35250 3278
rect 35982 3330 36034 3342
rect 35982 3266 36034 3278
rect 36542 3330 36594 3342
rect 36542 3266 36594 3278
rect 37214 3330 37266 3342
rect 37214 3266 37266 3278
rect 37886 3330 37938 3342
rect 37886 3266 37938 3278
rect 38558 3330 38610 3342
rect 38558 3266 38610 3278
rect 39118 3330 39170 3342
rect 39118 3266 39170 3278
rect 40574 3330 40626 3342
rect 40574 3266 40626 3278
rect 47406 3330 47458 3342
rect 47406 3266 47458 3278
rect 47854 3330 47906 3342
rect 47854 3266 47906 3278
rect 48302 3330 48354 3342
rect 48302 3266 48354 3278
rect 48750 3330 48802 3342
rect 48750 3266 48802 3278
rect 49310 3330 49362 3342
rect 49310 3266 49362 3278
rect 49982 3330 50034 3342
rect 49982 3266 50034 3278
rect 50654 3330 50706 3342
rect 50654 3266 50706 3278
rect 1344 3162 78624 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 78624 3162
rect 1344 3076 78624 3110
rect 47058 1822 47070 1874
rect 47122 1871 47134 1874
rect 47842 1871 47854 1874
rect 47122 1825 47854 1871
rect 47122 1822 47134 1825
rect 47842 1822 47854 1825
rect 47906 1822 47918 1874
rect 45826 926 45838 978
rect 45890 975 45902 978
rect 46610 975 46622 978
rect 45890 929 46622 975
rect 45890 926 45902 929
rect 46610 926 46622 929
rect 46674 926 46686 978
<< via1 >>
rect 43710 77198 43762 77250
rect 44270 77198 44322 77250
rect 54462 77198 54514 77250
rect 55246 77198 55298 77250
rect 27470 76974 27522 77026
rect 28254 76974 28306 77026
rect 30830 76974 30882 77026
rect 31726 76974 31778 77026
rect 53790 76974 53842 77026
rect 54462 76974 54514 77026
rect 56478 76974 56530 77026
rect 57038 76974 57090 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 23102 76638 23154 76690
rect 23998 76638 24050 76690
rect 25230 76638 25282 76690
rect 25790 76638 25842 76690
rect 26462 76638 26514 76690
rect 27022 76638 27074 76690
rect 32510 76638 32562 76690
rect 33182 76638 33234 76690
rect 35198 76638 35250 76690
rect 36654 76638 36706 76690
rect 37886 76638 37938 76690
rect 39902 76638 39954 76690
rect 44270 76638 44322 76690
rect 44718 76638 44770 76690
rect 45278 76638 45330 76690
rect 45950 76638 46002 76690
rect 47966 76638 48018 76690
rect 52222 76638 52274 76690
rect 54462 76638 54514 76690
rect 55358 76638 55410 76690
rect 55694 76638 55746 76690
rect 56142 76638 56194 76690
rect 57038 76638 57090 76690
rect 57374 76638 57426 76690
rect 58046 76638 58098 76690
rect 59838 76638 59890 76690
rect 24894 76526 24946 76578
rect 27470 76526 27522 76578
rect 27806 76526 27858 76578
rect 35982 76526 36034 76578
rect 36318 76526 36370 76578
rect 37214 76526 37266 76578
rect 37550 76526 37602 76578
rect 43598 76526 43650 76578
rect 48638 76526 48690 76578
rect 50318 76526 50370 76578
rect 54126 76526 54178 76578
rect 55022 76526 55074 76578
rect 56702 76526 56754 76578
rect 22878 76414 22930 76466
rect 24558 76414 24610 76466
rect 30830 76414 30882 76466
rect 42590 76414 42642 76466
rect 43822 76414 43874 76466
rect 47742 76414 47794 76466
rect 48862 76414 48914 76466
rect 50542 76414 50594 76466
rect 51214 76414 51266 76466
rect 58830 76414 58882 76466
rect 28590 76302 28642 76354
rect 31614 76302 31666 76354
rect 34302 76302 34354 76354
rect 34526 76302 34578 76354
rect 39118 76302 39170 76354
rect 41022 76302 41074 76354
rect 46622 76302 46674 76354
rect 49310 76302 49362 76354
rect 50094 76302 50146 76354
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 22654 75854 22706 75906
rect 30494 75854 30546 75906
rect 34078 75854 34130 75906
rect 38334 75854 38386 75906
rect 41582 75854 41634 75906
rect 28142 75742 28194 75794
rect 28702 75742 28754 75794
rect 37214 75742 37266 75794
rect 44046 75742 44098 75794
rect 50878 75742 50930 75794
rect 53790 75742 53842 75794
rect 55694 75742 55746 75794
rect 56702 75742 56754 75794
rect 25006 75630 25058 75682
rect 25454 75630 25506 75682
rect 29150 75630 29202 75682
rect 31726 75630 31778 75682
rect 36430 75630 36482 75682
rect 39790 75630 39842 75682
rect 40574 75630 40626 75682
rect 51662 75630 51714 75682
rect 52670 75630 52722 75682
rect 58494 75630 58546 75682
rect 29822 75518 29874 75570
rect 31166 75518 31218 75570
rect 43486 75518 43538 75570
rect 52110 75518 52162 75570
rect 56030 75518 56082 75570
rect 29486 75406 29538 75458
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 41918 75070 41970 75122
rect 52334 75070 52386 75122
rect 54350 75070 54402 75122
rect 51326 74846 51378 74898
rect 36654 74734 36706 74786
rect 40350 74734 40402 74786
rect 41022 74734 41074 74786
rect 43262 74734 43314 74786
rect 51102 74734 51154 74786
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 1934 67902 1986 67954
rect 4286 67790 4338 67842
rect 4734 67790 4786 67842
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 1710 67118 1762 67170
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 1710 65998 1762 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 1710 65550 1762 65602
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 2382 64766 2434 64818
rect 1710 64542 1762 64594
rect 2942 64542 2994 64594
rect 2046 64430 2098 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 1710 63982 1762 64034
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 1710 62862 1762 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 1710 62414 1762 62466
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 1710 61294 1762 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 2046 60846 2098 60898
rect 1710 60734 1762 60786
rect 2494 60622 2546 60674
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 2158 59838 2210 59890
rect 1710 59726 1762 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 1710 59278 1762 59330
rect 78206 59278 78258 59330
rect 77982 59166 78034 59218
rect 77534 59054 77586 59106
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 78206 58494 78258 58546
rect 1710 58158 1762 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 1710 57710 1762 57762
rect 75630 57598 75682 57650
rect 75406 57486 75458 57538
rect 77870 57486 77922 57538
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 1710 56590 1762 56642
rect 77646 56590 77698 56642
rect 77870 56590 77922 56642
rect 78206 56590 78258 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 1710 56142 1762 56194
rect 78206 56142 78258 56194
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 1710 55358 1762 55410
rect 2158 55134 2210 55186
rect 77758 55134 77810 55186
rect 78206 55022 78258 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 1710 54574 1762 54626
rect 75630 54462 75682 54514
rect 75406 54350 75458 54402
rect 77870 54350 77922 54402
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 78206 53790 78258 53842
rect 1822 53678 1874 53730
rect 2046 53454 2098 53506
rect 2494 53454 2546 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 1710 53006 1762 53058
rect 78206 52670 78258 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 1710 51886 1762 51938
rect 78206 51886 78258 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 1710 51438 1762 51490
rect 77870 51438 77922 51490
rect 78206 51326 78258 51378
rect 77646 51214 77698 51266
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 1710 50318 1762 50370
rect 2158 50318 2210 50370
rect 77758 50318 77810 50370
rect 78206 50318 78258 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 1710 49870 1762 49922
rect 78206 49870 78258 49922
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 1710 48750 1762 48802
rect 78206 48750 78258 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 39566 48414 39618 48466
rect 39790 48414 39842 48466
rect 43822 48414 43874 48466
rect 44382 48414 44434 48466
rect 1710 48302 1762 48354
rect 78206 48302 78258 48354
rect 40238 48078 40290 48130
rect 43374 48078 43426 48130
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 36430 47518 36482 47570
rect 1710 47182 1762 47234
rect 35534 47182 35586 47234
rect 35870 47182 35922 47234
rect 78206 47182 78258 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 34750 46846 34802 46898
rect 34974 46846 35026 46898
rect 43374 46846 43426 46898
rect 43934 46846 43986 46898
rect 47182 46846 47234 46898
rect 1710 46734 1762 46786
rect 46734 46734 46786 46786
rect 46510 46622 46562 46674
rect 75630 46622 75682 46674
rect 35422 46510 35474 46562
rect 42926 46510 42978 46562
rect 75406 46510 75458 46562
rect 77870 46510 77922 46562
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 2158 45726 2210 45778
rect 77758 45726 77810 45778
rect 1710 45614 1762 45666
rect 78206 45614 78258 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 45614 45278 45666 45330
rect 46174 45278 46226 45330
rect 78206 45166 78258 45218
rect 4286 45054 4338 45106
rect 4846 45054 4898 45106
rect 41470 45054 41522 45106
rect 42030 45054 42082 45106
rect 41022 44942 41074 44994
rect 45166 44942 45218 44994
rect 1934 44830 1986 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 34862 44382 34914 44434
rect 42702 44382 42754 44434
rect 44942 44382 44994 44434
rect 36430 44270 36482 44322
rect 34078 44158 34130 44210
rect 34414 44158 34466 44210
rect 43150 44158 43202 44210
rect 43598 44158 43650 44210
rect 1710 44046 1762 44098
rect 35534 44046 35586 44098
rect 35870 44046 35922 44098
rect 45390 44046 45442 44098
rect 45838 44046 45890 44098
rect 78206 44046 78258 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 78206 43710 78258 43762
rect 1710 43598 1762 43650
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 45838 42702 45890 42754
rect 1710 42478 1762 42530
rect 46398 42478 46450 42530
rect 46846 42478 46898 42530
rect 78206 42478 78258 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 78206 42030 78258 42082
rect 4286 41918 4338 41970
rect 38110 41918 38162 41970
rect 38334 41918 38386 41970
rect 38894 41918 38946 41970
rect 45390 41918 45442 41970
rect 45950 41918 46002 41970
rect 4846 41806 4898 41858
rect 44942 41806 44994 41858
rect 1934 41694 1986 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 34414 41246 34466 41298
rect 1710 41022 1762 41074
rect 78206 41022 78258 41074
rect 2158 40910 2210 40962
rect 33630 40910 33682 40962
rect 33966 40910 34018 40962
rect 77758 40910 77810 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 78206 40462 78258 40514
rect 34414 40350 34466 40402
rect 34638 40350 34690 40402
rect 35198 40350 35250 40402
rect 1710 40126 1762 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 40350 39678 40402 39730
rect 78206 39678 78258 39730
rect 41694 39566 41746 39618
rect 44830 39566 44882 39618
rect 1710 39342 1762 39394
rect 40014 39342 40066 39394
rect 40798 39342 40850 39394
rect 41134 39342 41186 39394
rect 45390 39342 45442 39394
rect 45950 39342 46002 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 2046 38894 2098 38946
rect 1710 38782 1762 38834
rect 35310 38782 35362 38834
rect 38334 38782 38386 38834
rect 39230 38782 39282 38834
rect 44046 38782 44098 38834
rect 2494 38670 2546 38722
rect 34974 38670 35026 38722
rect 35870 38670 35922 38722
rect 37998 38670 38050 38722
rect 38782 38670 38834 38722
rect 39790 38670 39842 38722
rect 41022 38670 41074 38722
rect 43710 38670 43762 38722
rect 44606 38670 44658 38722
rect 78206 38558 78258 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 33406 37998 33458 38050
rect 1710 37774 1762 37826
rect 32622 37774 32674 37826
rect 32846 37774 32898 37826
rect 38894 37774 38946 37826
rect 78206 37774 78258 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 2046 37326 2098 37378
rect 78206 37326 78258 37378
rect 1710 37214 1762 37266
rect 33854 37214 33906 37266
rect 2494 37102 2546 37154
rect 33518 37102 33570 37154
rect 34414 37102 34466 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 77758 36542 77810 36594
rect 34974 36430 35026 36482
rect 1710 36318 1762 36370
rect 2046 36318 2098 36370
rect 2942 36318 2994 36370
rect 78206 36318 78258 36370
rect 2382 36206 2434 36258
rect 34190 36206 34242 36258
rect 34414 36206 34466 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 1710 35758 1762 35810
rect 40126 35646 40178 35698
rect 43150 35646 43202 35698
rect 44158 35646 44210 35698
rect 33630 35534 33682 35586
rect 33854 35534 33906 35586
rect 34078 35534 34130 35586
rect 39566 35534 39618 35586
rect 41022 35534 41074 35586
rect 43598 35534 43650 35586
rect 78206 35422 78258 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 45278 34974 45330 35026
rect 1822 34862 1874 34914
rect 2046 34638 2098 34690
rect 2494 34638 2546 34690
rect 44382 34638 44434 34690
rect 44830 34638 44882 34690
rect 78206 34638 78258 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 1710 34190 1762 34242
rect 77870 34190 77922 34242
rect 34190 34078 34242 34130
rect 34638 34078 34690 34130
rect 46622 34078 46674 34130
rect 78206 34078 78258 34130
rect 35086 33966 35138 34018
rect 46062 33966 46114 34018
rect 47070 33966 47122 34018
rect 77646 33966 77698 34018
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 1710 33406 1762 33458
rect 40462 33294 40514 33346
rect 41022 33070 41074 33122
rect 41582 33070 41634 33122
rect 78206 33070 78258 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 2046 32622 2098 32674
rect 78206 32622 78258 32674
rect 1710 32510 1762 32562
rect 44046 32510 44098 32562
rect 44494 32510 44546 32562
rect 2494 32398 2546 32450
rect 43486 32398 43538 32450
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 77758 31950 77810 32002
rect 1934 31838 1986 31890
rect 4286 31726 4338 31778
rect 4846 31726 4898 31778
rect 78206 31614 78258 31666
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 2942 31166 2994 31218
rect 1710 31054 1762 31106
rect 2046 31054 2098 31106
rect 75630 30942 75682 30994
rect 75294 30830 75346 30882
rect 2382 30718 2434 30770
rect 77982 30718 78034 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 4286 30158 4338 30210
rect 2494 30046 2546 30098
rect 4846 29934 4898 29986
rect 78206 29934 78258 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 78206 29486 78258 29538
rect 1710 29150 1762 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 1934 28702 1986 28754
rect 4286 28590 4338 28642
rect 4846 28590 4898 28642
rect 78206 28366 78258 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 1710 27918 1762 27970
rect 78206 27918 78258 27970
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 77198 27134 77250 27186
rect 77870 26910 77922 26962
rect 78206 26910 78258 26962
rect 1710 26798 1762 26850
rect 2158 26798 2210 26850
rect 77534 26798 77586 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 1710 26350 1762 26402
rect 75630 26238 75682 26290
rect 75294 26126 75346 26178
rect 77982 26014 78034 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 1710 25230 1762 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 1710 24782 1762 24834
rect 75742 24670 75794 24722
rect 75294 24558 75346 24610
rect 77982 24558 78034 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 78206 23774 78258 23826
rect 1710 23662 1762 23714
rect 77758 23662 77810 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 1710 23214 1762 23266
rect 75742 23102 75794 23154
rect 75294 22990 75346 23042
rect 77982 22878 78034 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 1934 22430 1986 22482
rect 4286 22318 4338 22370
rect 4846 22318 4898 22370
rect 78206 22206 78258 22258
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 1710 21758 1762 21810
rect 2942 21758 2994 21810
rect 2046 21646 2098 21698
rect 2382 21646 2434 21698
rect 75630 21534 75682 21586
rect 75294 21422 75346 21474
rect 77982 21422 78034 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 77646 20862 77698 20914
rect 78206 20750 78258 20802
rect 1710 20526 1762 20578
rect 77870 20526 77922 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 2046 20078 2098 20130
rect 1710 19966 1762 20018
rect 75630 19966 75682 20018
rect 2494 19854 2546 19906
rect 75294 19854 75346 19906
rect 77982 19854 78034 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 1710 18958 1762 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 1710 18510 1762 18562
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 1934 17726 1986 17778
rect 4286 17614 4338 17666
rect 4846 17390 4898 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 1710 17054 1762 17106
rect 2942 17054 2994 17106
rect 2046 16942 2098 16994
rect 2382 16942 2434 16994
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 1710 15822 1762 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 1710 15374 1762 15426
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 1710 14254 1762 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 1710 13470 1762 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 1934 13022 1986 13074
rect 4286 12910 4338 12962
rect 4846 12686 4898 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 1710 12350 1762 12402
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 43262 4846 43314 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 36878 4510 36930 4562
rect 42478 4510 42530 4562
rect 46174 4398 46226 4450
rect 46622 4398 46674 4450
rect 29598 4286 29650 4338
rect 35982 4286 36034 4338
rect 43374 4286 43426 4338
rect 51998 4286 52050 4338
rect 30158 4174 30210 4226
rect 41134 4174 41186 4226
rect 41694 4174 41746 4226
rect 43038 4174 43090 4226
rect 47182 4174 47234 4226
rect 50878 4174 50930 4226
rect 51662 4174 51714 4226
rect 27358 4062 27410 4114
rect 34078 4062 34130 4114
rect 42814 4062 42866 4114
rect 43038 4062 43090 4114
rect 44270 4062 44322 4114
rect 53006 4062 53058 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 29150 3614 29202 3666
rect 29822 3614 29874 3666
rect 30494 3614 30546 3666
rect 31614 3614 31666 3666
rect 39902 3614 39954 3666
rect 44606 3614 44658 3666
rect 52222 3614 52274 3666
rect 27246 3502 27298 3554
rect 27582 3502 27634 3554
rect 42142 3502 42194 3554
rect 42814 3502 42866 3554
rect 43710 3502 43762 3554
rect 46734 3502 46786 3554
rect 51214 3502 51266 3554
rect 26798 3390 26850 3442
rect 27806 3390 27858 3442
rect 28478 3390 28530 3442
rect 28814 3390 28866 3442
rect 41246 3390 41298 3442
rect 41582 3390 41634 3442
rect 41918 3390 41970 3442
rect 43038 3390 43090 3442
rect 46510 3390 46562 3442
rect 31054 3278 31106 3330
rect 32510 3278 32562 3330
rect 33182 3278 33234 3330
rect 34526 3278 34578 3330
rect 35198 3278 35250 3330
rect 35982 3278 36034 3330
rect 36542 3278 36594 3330
rect 37214 3278 37266 3330
rect 37886 3278 37938 3330
rect 38558 3278 38610 3330
rect 39118 3278 39170 3330
rect 40574 3278 40626 3330
rect 47406 3278 47458 3330
rect 47854 3278 47906 3330
rect 48302 3278 48354 3330
rect 48750 3278 48802 3330
rect 49310 3278 49362 3330
rect 49982 3278 50034 3330
rect 50654 3278 50706 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 47070 1822 47122 1874
rect 47854 1822 47906 1874
rect 45838 926 45890 978
rect 46622 926 46674 978
<< metal2 >>
rect 0 79200 112 80000
rect 672 79200 784 80000
rect 1344 79200 1456 80000
rect 2016 79200 2128 80000
rect 2688 79200 2800 80000
rect 3360 79200 3472 80000
rect 4032 79200 4144 80000
rect 4704 79200 4816 80000
rect 5376 79200 5488 80000
rect 6048 79200 6160 80000
rect 6720 79200 6832 80000
rect 7392 79200 7504 80000
rect 8064 79200 8176 80000
rect 8736 79200 8848 80000
rect 9408 79200 9520 80000
rect 10080 79200 10192 80000
rect 10752 79200 10864 80000
rect 11424 79200 11536 80000
rect 12096 79200 12208 80000
rect 12768 79200 12880 80000
rect 13440 79200 13552 80000
rect 14112 79200 14224 80000
rect 14784 79200 14896 80000
rect 15456 79200 15568 80000
rect 16128 79200 16240 80000
rect 16800 79200 16912 80000
rect 17472 79200 17584 80000
rect 18144 79200 18256 80000
rect 18816 79200 18928 80000
rect 19488 79200 19600 80000
rect 20160 79200 20272 80000
rect 20832 79200 20944 80000
rect 21504 79200 21616 80000
rect 22176 79200 22288 80000
rect 22848 79200 22960 80000
rect 23520 79200 23632 80000
rect 24192 79200 24304 80000
rect 24864 79200 24976 80000
rect 25536 79200 25648 80000
rect 26208 79200 26320 80000
rect 26880 79200 26992 80000
rect 27552 79200 27664 80000
rect 28224 79200 28336 80000
rect 28896 79200 29008 80000
rect 29568 79200 29680 80000
rect 30240 79200 30352 80000
rect 30912 79200 31024 80000
rect 31584 79200 31696 80000
rect 32256 79200 32368 80000
rect 32928 79200 33040 80000
rect 33600 79200 33712 80000
rect 34272 79200 34384 80000
rect 34944 79200 35056 80000
rect 35616 79200 35728 80000
rect 36288 79200 36400 80000
rect 36960 79200 37072 80000
rect 37632 79200 37744 80000
rect 38304 79200 38416 80000
rect 38976 79200 39088 80000
rect 39648 79200 39760 80000
rect 40320 79200 40432 80000
rect 40992 79200 41104 80000
rect 41664 79200 41776 80000
rect 42336 79200 42448 80000
rect 43008 79200 43120 80000
rect 43680 79200 43792 80000
rect 44352 79200 44464 80000
rect 45024 79200 45136 80000
rect 45696 79200 45808 80000
rect 46368 79200 46480 80000
rect 47040 79200 47152 80000
rect 47712 79200 47824 80000
rect 48384 79200 48496 80000
rect 49056 79200 49168 80000
rect 49728 79200 49840 80000
rect 50400 79200 50512 80000
rect 51072 79200 51184 80000
rect 51744 79200 51856 80000
rect 52416 79200 52528 80000
rect 53088 79200 53200 80000
rect 53760 79200 53872 80000
rect 54432 79200 54544 80000
rect 55104 79200 55216 80000
rect 55776 79200 55888 80000
rect 56448 79200 56560 80000
rect 57120 79200 57232 80000
rect 57792 79200 57904 80000
rect 58464 79200 58576 80000
rect 59136 79200 59248 80000
rect 59808 79200 59920 80000
rect 60480 79200 60592 80000
rect 61152 79200 61264 80000
rect 61824 79200 61936 80000
rect 62496 79200 62608 80000
rect 63168 79200 63280 80000
rect 63840 79200 63952 80000
rect 64512 79200 64624 80000
rect 65184 79200 65296 80000
rect 65856 79200 65968 80000
rect 66528 79200 66640 80000
rect 67200 79200 67312 80000
rect 67872 79200 67984 80000
rect 68544 79200 68656 80000
rect 69216 79200 69328 80000
rect 69888 79200 70000 80000
rect 70560 79200 70672 80000
rect 71232 79200 71344 80000
rect 71904 79200 72016 80000
rect 72576 79200 72688 80000
rect 73248 79200 73360 80000
rect 73920 79200 74032 80000
rect 74592 79200 74704 80000
rect 75264 79200 75376 80000
rect 75936 79200 76048 80000
rect 76608 79200 76720 80000
rect 77280 79200 77392 80000
rect 77952 79200 78064 80000
rect 78624 79200 78736 80000
rect 79296 79200 79408 80000
rect 22204 77364 22260 79200
rect 22204 77308 22708 77364
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 22652 75906 22708 77308
rect 22876 76692 22932 79200
rect 23100 76692 23156 76702
rect 22876 76690 23156 76692
rect 22876 76638 23102 76690
rect 23154 76638 23156 76690
rect 22876 76636 23156 76638
rect 23100 76626 23156 76636
rect 22876 76468 22932 76478
rect 22876 76374 22932 76412
rect 23548 76468 23604 79200
rect 23996 76692 24052 76702
rect 24220 76692 24276 79200
rect 24892 77700 24948 79200
rect 24892 77644 25172 77700
rect 23996 76690 24276 76692
rect 23996 76638 23998 76690
rect 24050 76638 24276 76690
rect 23996 76636 24276 76638
rect 25116 76692 25172 77644
rect 25228 76692 25284 76702
rect 25116 76690 25284 76692
rect 25116 76638 25230 76690
rect 25282 76638 25284 76690
rect 25116 76636 25284 76638
rect 25564 76692 25620 79200
rect 25788 76692 25844 76702
rect 25564 76690 25844 76692
rect 25564 76638 25790 76690
rect 25842 76638 25844 76690
rect 25564 76636 25844 76638
rect 26236 76692 26292 79200
rect 26460 76692 26516 76702
rect 26236 76690 26516 76692
rect 26236 76638 26462 76690
rect 26514 76638 26516 76690
rect 26236 76636 26516 76638
rect 26908 76692 26964 79200
rect 27468 77026 27524 77038
rect 27468 76974 27470 77026
rect 27522 76974 27524 77026
rect 27020 76692 27076 76702
rect 26908 76690 27076 76692
rect 26908 76638 27022 76690
rect 27074 76638 27076 76690
rect 26908 76636 27076 76638
rect 23996 76626 24052 76636
rect 25228 76626 25284 76636
rect 25788 76626 25844 76636
rect 26460 76626 26516 76636
rect 27020 76626 27076 76636
rect 24892 76578 24948 76590
rect 24892 76526 24894 76578
rect 24946 76526 24948 76578
rect 23548 76402 23604 76412
rect 24556 76468 24612 76478
rect 24556 76374 24612 76412
rect 22652 75854 22654 75906
rect 22706 75854 22708 75906
rect 22652 75842 22708 75854
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 1932 67954 1988 67966
rect 1932 67902 1934 67954
rect 1986 67902 1988 67954
rect 1932 67284 1988 67902
rect 4284 67844 4340 67854
rect 4732 67844 4788 67854
rect 4284 67842 4788 67844
rect 4284 67790 4286 67842
rect 4338 67790 4734 67842
rect 4786 67790 4788 67842
rect 4284 67788 4788 67790
rect 4284 67778 4340 67788
rect 1932 67218 1988 67228
rect 4732 67228 4788 67788
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 24892 67228 24948 76526
rect 27468 76578 27524 76974
rect 27468 76526 27470 76578
rect 27522 76526 27524 76578
rect 27468 76514 27524 76526
rect 27580 76356 27636 79200
rect 28252 77028 28308 79200
rect 28140 77026 28308 77028
rect 28140 76974 28254 77026
rect 28306 76974 28308 77026
rect 28140 76972 28308 76974
rect 27580 76290 27636 76300
rect 27804 76578 27860 76590
rect 27804 76526 27806 76578
rect 27858 76526 27860 76578
rect 25004 75684 25060 75694
rect 25452 75684 25508 75694
rect 25004 75682 25508 75684
rect 25004 75630 25006 75682
rect 25058 75630 25454 75682
rect 25506 75630 25508 75682
rect 25004 75628 25508 75630
rect 25004 75618 25060 75628
rect 1708 67170 1764 67182
rect 4732 67172 5012 67228
rect 24892 67172 25060 67228
rect 1708 67118 1710 67170
rect 1762 67118 1764 67170
rect 1708 66612 1764 67118
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 1708 66546 1764 66556
rect 1708 66052 1764 66062
rect 1708 65958 1764 65996
rect 1708 65602 1764 65614
rect 1708 65550 1710 65602
rect 1762 65550 1764 65602
rect 1708 65268 1764 65550
rect 1708 65202 1764 65212
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 2380 64818 2436 64830
rect 2380 64766 2382 64818
rect 2434 64766 2436 64818
rect 1708 64596 1764 64606
rect 1708 64502 1764 64540
rect 2044 64484 2100 64494
rect 1932 64482 2100 64484
rect 1932 64430 2046 64482
rect 2098 64430 2100 64482
rect 1932 64428 2100 64430
rect 1708 64034 1764 64046
rect 1708 63982 1710 64034
rect 1762 63982 1764 64034
rect 1708 63252 1764 63982
rect 1708 63186 1764 63196
rect 1708 62916 1764 62926
rect 1708 62822 1764 62860
rect 1708 62466 1764 62478
rect 1708 62414 1710 62466
rect 1762 62414 1764 62466
rect 1708 61908 1764 62414
rect 1708 61842 1764 61852
rect 1708 61348 1764 61358
rect 1708 61254 1764 61292
rect 1708 60786 1764 60798
rect 1708 60734 1710 60786
rect 1762 60734 1764 60786
rect 1708 60564 1764 60734
rect 1708 60498 1764 60508
rect 1708 59780 1764 59790
rect 1708 59778 1876 59780
rect 1708 59726 1710 59778
rect 1762 59726 1876 59778
rect 1708 59724 1876 59726
rect 1708 59714 1764 59724
rect 1708 59330 1764 59342
rect 1708 59278 1710 59330
rect 1762 59278 1764 59330
rect 1708 58548 1764 59278
rect 1820 59220 1876 59724
rect 1820 59154 1876 59164
rect 1708 58482 1764 58492
rect 1708 58212 1764 58222
rect 1708 58118 1764 58156
rect 1708 57762 1764 57774
rect 1708 57710 1710 57762
rect 1762 57710 1764 57762
rect 1708 57204 1764 57710
rect 1708 57138 1764 57148
rect 1708 56644 1764 56654
rect 1708 56550 1764 56588
rect 1708 56194 1764 56206
rect 1708 56142 1710 56194
rect 1762 56142 1764 56194
rect 1708 55860 1764 56142
rect 1708 55794 1764 55804
rect 1708 55410 1764 55422
rect 1708 55358 1710 55410
rect 1762 55358 1764 55410
rect 1708 54964 1764 55358
rect 1708 54898 1764 54908
rect 1708 54626 1764 54638
rect 1708 54574 1710 54626
rect 1762 54574 1764 54626
rect 1708 53844 1764 54574
rect 1708 53778 1764 53788
rect 1820 53730 1876 53742
rect 1820 53678 1822 53730
rect 1874 53678 1876 53730
rect 1820 53172 1876 53678
rect 1820 53106 1876 53116
rect 1708 53058 1764 53070
rect 1708 53006 1710 53058
rect 1762 53006 1764 53058
rect 1708 52500 1764 53006
rect 1708 52434 1764 52444
rect 1708 51940 1764 51950
rect 1708 51846 1764 51884
rect 1708 51490 1764 51502
rect 1708 51438 1710 51490
rect 1762 51438 1764 51490
rect 1708 51156 1764 51438
rect 1708 51090 1764 51100
rect 1708 50372 1764 50382
rect 1708 50370 1876 50372
rect 1708 50318 1710 50370
rect 1762 50318 1876 50370
rect 1708 50316 1876 50318
rect 1708 50306 1764 50316
rect 1708 49922 1764 49934
rect 1708 49870 1710 49922
rect 1762 49870 1764 49922
rect 1708 49140 1764 49870
rect 1820 49812 1876 50316
rect 1820 49746 1876 49756
rect 1932 49700 1988 64428
rect 2044 64418 2100 64428
rect 2380 63924 2436 64766
rect 2940 64596 2996 64606
rect 2940 64502 2996 64540
rect 2380 63858 2436 63868
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 2044 60898 2100 60910
rect 2044 60846 2046 60898
rect 2098 60846 2100 60898
rect 2044 55468 2100 60846
rect 2492 60674 2548 60686
rect 2492 60622 2494 60674
rect 2546 60622 2548 60674
rect 2492 60564 2548 60622
rect 2492 60498 2548 60508
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 2156 59892 2212 59902
rect 2156 59798 2212 59836
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 2044 55412 2660 55468
rect 2156 55188 2212 55198
rect 2156 55094 2212 55132
rect 2044 53508 2100 53518
rect 2044 53506 2436 53508
rect 2044 53454 2046 53506
rect 2098 53454 2436 53506
rect 2044 53452 2436 53454
rect 2044 53442 2100 53452
rect 2156 50484 2212 50494
rect 2156 50370 2212 50428
rect 2156 50318 2158 50370
rect 2210 50318 2212 50370
rect 2156 50306 2212 50318
rect 1932 49644 2100 49700
rect 1708 49074 1764 49084
rect 1708 48802 1764 48814
rect 1708 48750 1710 48802
rect 1762 48750 1764 48802
rect 1708 48580 1764 48750
rect 1708 48514 1764 48524
rect 1708 48354 1764 48366
rect 1708 48302 1710 48354
rect 1762 48302 1764 48354
rect 1708 47796 1764 48302
rect 1708 47730 1764 47740
rect 1708 47236 1764 47246
rect 1708 47142 1764 47180
rect 1708 46786 1764 46798
rect 1708 46734 1710 46786
rect 1762 46734 1764 46786
rect 1708 46452 1764 46734
rect 1708 46386 1764 46396
rect 1708 45666 1764 45678
rect 1708 45614 1710 45666
rect 1762 45614 1764 45666
rect 1708 45108 1764 45614
rect 1708 45042 1764 45052
rect 1932 44882 1988 44894
rect 1932 44830 1934 44882
rect 1986 44830 1988 44882
rect 1932 44436 1988 44830
rect 1932 44370 1988 44380
rect 1708 44100 1764 44110
rect 1708 44006 1764 44044
rect 2044 43708 2100 49644
rect 2156 45780 2212 45790
rect 2156 45686 2212 45724
rect 2380 44212 2436 53452
rect 2492 53506 2548 53518
rect 2492 53454 2494 53506
rect 2546 53454 2548 53506
rect 2492 53172 2548 53454
rect 2492 53106 2548 53116
rect 2380 44146 2436 44156
rect 1708 43650 1764 43662
rect 2044 43652 2436 43708
rect 1708 43598 1710 43650
rect 1762 43598 1764 43650
rect 1708 43092 1764 43598
rect 1708 43026 1764 43036
rect 1708 42532 1764 42542
rect 1708 42438 1764 42476
rect 1932 41748 1988 41758
rect 1932 41654 1988 41692
rect 1708 41076 1764 41086
rect 1708 40982 1764 41020
rect 2156 40962 2212 40974
rect 2156 40910 2158 40962
rect 2210 40910 2212 40962
rect 2156 40404 2212 40910
rect 2156 40338 2212 40348
rect 2380 40404 2436 43652
rect 2604 40964 2660 55412
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4284 45108 4340 45118
rect 4284 45014 4340 45052
rect 4844 45108 4900 45118
rect 4844 45014 4900 45052
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4284 41970 4340 41982
rect 4284 41918 4286 41970
rect 4338 41918 4340 41970
rect 4284 41860 4340 41918
rect 4284 41794 4340 41804
rect 4844 41860 4900 41870
rect 4844 41766 4900 41804
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 2604 40898 2660 40908
rect 4956 40516 5012 67172
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 25004 46900 25060 67172
rect 25004 46834 25060 46844
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 25452 44324 25508 75628
rect 25452 44258 25508 44268
rect 27804 44100 27860 76526
rect 28140 75794 28196 76972
rect 28252 76962 28308 76972
rect 28588 76356 28644 76366
rect 28588 76262 28644 76300
rect 28140 75742 28142 75794
rect 28194 75742 28196 75794
rect 28140 75730 28196 75742
rect 28700 75796 28756 75806
rect 28924 75796 28980 79200
rect 28700 75794 28980 75796
rect 28700 75742 28702 75794
rect 28754 75742 28980 75794
rect 28700 75740 28980 75742
rect 28700 75730 28756 75740
rect 28924 75684 28980 75740
rect 29148 75684 29204 75694
rect 28924 75682 29204 75684
rect 28924 75630 29150 75682
rect 29202 75630 29204 75682
rect 28924 75628 29204 75630
rect 29148 75618 29204 75628
rect 29596 75572 29652 79200
rect 30268 75908 30324 79200
rect 30828 77026 30884 77038
rect 30828 76974 30830 77026
rect 30882 76974 30884 77026
rect 30828 76466 30884 76974
rect 30828 76414 30830 76466
rect 30882 76414 30884 76466
rect 30828 76402 30884 76414
rect 30492 75908 30548 75918
rect 30268 75906 30548 75908
rect 30268 75854 30494 75906
rect 30546 75854 30548 75906
rect 30268 75852 30548 75854
rect 30492 75842 30548 75852
rect 29820 75572 29876 75582
rect 29596 75570 29876 75572
rect 29596 75518 29822 75570
rect 29874 75518 29876 75570
rect 29596 75516 29876 75518
rect 30940 75572 30996 79200
rect 31612 76354 31668 79200
rect 31612 76302 31614 76354
rect 31666 76302 31668 76354
rect 31612 76290 31668 76302
rect 31724 77026 31780 77038
rect 31724 76974 31726 77026
rect 31778 76974 31780 77026
rect 31724 75682 31780 76974
rect 32284 76692 32340 79200
rect 32508 76692 32564 76702
rect 32284 76690 32564 76692
rect 32284 76638 32510 76690
rect 32562 76638 32564 76690
rect 32284 76636 32564 76638
rect 32956 76692 33012 79200
rect 33628 77364 33684 79200
rect 33628 77308 34132 77364
rect 33180 76692 33236 76702
rect 32956 76690 33236 76692
rect 32956 76638 33182 76690
rect 33234 76638 33236 76690
rect 32956 76636 33236 76638
rect 32508 76626 32564 76636
rect 33180 76626 33236 76636
rect 34076 75906 34132 77308
rect 34300 76580 34356 79200
rect 34972 76692 35028 79200
rect 35644 77476 35700 79200
rect 36316 77924 36372 79200
rect 36316 77868 36708 77924
rect 35644 77420 36036 77476
rect 35196 76692 35252 76702
rect 34972 76690 35252 76692
rect 34972 76638 35198 76690
rect 35250 76638 35252 76690
rect 34972 76636 35252 76638
rect 35196 76626 35252 76636
rect 34300 76524 34580 76580
rect 34300 76356 34356 76366
rect 34300 76262 34356 76300
rect 34524 76354 34580 76524
rect 34524 76302 34526 76354
rect 34578 76302 34580 76354
rect 34524 76290 34580 76302
rect 35980 76578 36036 77420
rect 36652 76690 36708 77868
rect 36652 76638 36654 76690
rect 36706 76638 36708 76690
rect 36652 76626 36708 76638
rect 35980 76526 35982 76578
rect 36034 76526 36036 76578
rect 35980 76356 36036 76526
rect 35980 76290 36036 76300
rect 36316 76578 36372 76590
rect 36316 76526 36318 76578
rect 36370 76526 36372 76578
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 34076 75854 34078 75906
rect 34130 75854 34132 75906
rect 34076 75842 34132 75854
rect 31724 75630 31726 75682
rect 31778 75630 31780 75682
rect 31164 75572 31220 75582
rect 30940 75570 31220 75572
rect 30940 75518 31166 75570
rect 31218 75518 31220 75570
rect 30940 75516 31220 75518
rect 29820 75506 29876 75516
rect 31164 75506 31220 75516
rect 29484 75458 29540 75470
rect 29484 75406 29486 75458
rect 29538 75406 29540 75458
rect 29484 47236 29540 75406
rect 29484 47170 29540 47180
rect 31724 46676 31780 75630
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 36316 48468 36372 76526
rect 36988 76580 37044 79200
rect 37660 76692 37716 79200
rect 37884 76692 37940 76702
rect 37660 76690 37940 76692
rect 37660 76638 37886 76690
rect 37938 76638 37940 76690
rect 37660 76636 37940 76638
rect 37884 76626 37940 76636
rect 37212 76580 37268 76590
rect 36988 76578 37268 76580
rect 36988 76526 37214 76578
rect 37266 76526 37268 76578
rect 36988 76524 37268 76526
rect 37212 75794 37268 76524
rect 37212 75742 37214 75794
rect 37266 75742 37268 75794
rect 37212 75730 37268 75742
rect 37548 76578 37604 76590
rect 37548 76526 37550 76578
rect 37602 76526 37604 76578
rect 36428 75682 36484 75694
rect 36428 75630 36430 75682
rect 36482 75630 36484 75682
rect 36428 74788 36484 75630
rect 36652 74788 36708 74798
rect 36428 74786 36708 74788
rect 36428 74734 36654 74786
rect 36706 74734 36708 74786
rect 36428 74732 36708 74734
rect 36652 55468 36708 74732
rect 37548 67228 37604 76526
rect 38332 75906 38388 79200
rect 39004 76356 39060 79200
rect 39676 76692 39732 79200
rect 39900 76692 39956 76702
rect 39676 76690 39956 76692
rect 39676 76638 39902 76690
rect 39954 76638 39956 76690
rect 39676 76636 39956 76638
rect 39900 76626 39956 76636
rect 39116 76356 39172 76366
rect 39004 76354 39172 76356
rect 39004 76302 39118 76354
rect 39170 76302 39172 76354
rect 39004 76300 39172 76302
rect 39116 76290 39172 76300
rect 38332 75854 38334 75906
rect 38386 75854 38388 75906
rect 38332 75842 38388 75854
rect 40348 75908 40404 79200
rect 41020 76354 41076 79200
rect 41020 76302 41022 76354
rect 41074 76302 41076 76354
rect 41020 76290 41076 76302
rect 40348 75842 40404 75852
rect 41580 75908 41636 75918
rect 41580 75814 41636 75852
rect 39788 75682 39844 75694
rect 39788 75630 39790 75682
rect 39842 75630 39844 75682
rect 39788 74788 39844 75630
rect 40572 75682 40628 75694
rect 40572 75630 40574 75682
rect 40626 75630 40628 75682
rect 40348 74788 40404 74798
rect 40572 74788 40628 75630
rect 41692 75124 41748 79200
rect 42364 77252 42420 79200
rect 43036 77588 43092 79200
rect 43036 77532 43540 77588
rect 42364 77196 43428 77252
rect 42588 76466 42644 76478
rect 42588 76414 42590 76466
rect 42642 76414 42644 76466
rect 41916 75124 41972 75134
rect 41692 75122 41972 75124
rect 41692 75070 41918 75122
rect 41970 75070 41972 75122
rect 41692 75068 41972 75070
rect 41916 75058 41972 75068
rect 38892 74004 38948 74014
rect 37548 67172 38388 67228
rect 36316 48402 36372 48412
rect 36428 55412 36708 55468
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 36428 47570 36484 55412
rect 36428 47518 36430 47570
rect 36482 47518 36484 47570
rect 36428 47506 36484 47518
rect 35532 47236 35588 47246
rect 35868 47236 35924 47246
rect 35588 47234 35924 47236
rect 35588 47182 35870 47234
rect 35922 47182 35924 47234
rect 35588 47180 35924 47182
rect 35532 47142 35588 47180
rect 35868 47170 35924 47180
rect 34748 46900 34804 46910
rect 34972 46900 35028 46910
rect 34804 46898 35028 46900
rect 34804 46846 34974 46898
rect 35026 46846 35028 46898
rect 34804 46844 35028 46846
rect 34748 46806 34804 46844
rect 34972 46834 35028 46844
rect 31724 46610 31780 46620
rect 35420 46676 35476 46686
rect 35420 46562 35476 46620
rect 35420 46510 35422 46562
rect 35474 46510 35476 46562
rect 35420 46498 35476 46510
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34860 45108 34916 45118
rect 34860 44434 34916 45052
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34860 44382 34862 44434
rect 34914 44382 34916 44434
rect 34860 44370 34916 44382
rect 36428 44324 36484 44334
rect 36428 44230 36484 44268
rect 34076 44212 34132 44222
rect 34412 44212 34468 44222
rect 34132 44210 34468 44212
rect 34132 44158 34414 44210
rect 34466 44158 34468 44210
rect 34132 44156 34468 44158
rect 34076 44118 34132 44156
rect 34412 44146 34468 44156
rect 27804 44034 27860 44044
rect 35532 44100 35588 44110
rect 35868 44100 35924 44110
rect 35588 44098 35924 44100
rect 35588 44046 35870 44098
rect 35922 44046 35924 44098
rect 35588 44044 35924 44046
rect 35532 44006 35588 44044
rect 35868 44034 35924 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 38108 41972 38164 41982
rect 38332 41972 38388 67172
rect 38108 41970 38388 41972
rect 38108 41918 38110 41970
rect 38162 41918 38334 41970
rect 38386 41918 38388 41970
rect 38108 41916 38388 41918
rect 38108 41906 38164 41916
rect 38332 41906 38388 41916
rect 38892 41970 38948 73948
rect 39788 74004 39844 74732
rect 39788 73938 39844 73948
rect 40236 74786 40628 74788
rect 40236 74734 40350 74786
rect 40402 74734 40628 74786
rect 40236 74732 40628 74734
rect 41020 74788 41076 74798
rect 39564 48468 39620 48478
rect 39788 48468 39844 48478
rect 39620 48466 39844 48468
rect 39620 48414 39790 48466
rect 39842 48414 39844 48466
rect 39620 48412 39844 48414
rect 39564 48374 39620 48412
rect 39788 48402 39844 48412
rect 40236 48130 40292 74732
rect 40348 74722 40404 74732
rect 41020 74694 41076 74732
rect 41244 74788 41300 74798
rect 41244 55468 41300 74732
rect 42588 74788 42644 76414
rect 43372 75572 43428 77196
rect 43484 77028 43540 77532
rect 43708 77250 43764 79200
rect 44380 77924 44436 79200
rect 44380 77868 44772 77924
rect 43708 77198 43710 77250
rect 43762 77198 43764 77250
rect 43708 77186 43764 77198
rect 44268 77250 44324 77262
rect 44268 77198 44270 77250
rect 44322 77198 44324 77250
rect 43484 76972 43876 77028
rect 43596 76578 43652 76590
rect 43596 76526 43598 76578
rect 43650 76526 43652 76578
rect 43484 75572 43540 75582
rect 43372 75570 43540 75572
rect 43372 75518 43486 75570
rect 43538 75518 43540 75570
rect 43372 75516 43540 75518
rect 43484 75506 43540 75516
rect 42588 74722 42644 74732
rect 43260 74788 43316 74798
rect 43260 74694 43316 74732
rect 43596 55468 43652 76526
rect 43820 76468 43876 76972
rect 44268 76690 44324 77198
rect 44268 76638 44270 76690
rect 44322 76638 44324 76690
rect 44268 76626 44324 76638
rect 44716 76690 44772 77868
rect 44716 76638 44718 76690
rect 44770 76638 44772 76690
rect 44716 76626 44772 76638
rect 45052 76692 45108 79200
rect 45276 76692 45332 76702
rect 45052 76690 45332 76692
rect 45052 76638 45278 76690
rect 45330 76638 45332 76690
rect 45052 76636 45332 76638
rect 45724 76692 45780 79200
rect 45948 76692 46004 76702
rect 45724 76690 46004 76692
rect 45724 76638 45950 76690
rect 46002 76638 46004 76690
rect 45724 76636 46004 76638
rect 45276 76626 45332 76636
rect 45948 76626 46004 76636
rect 43820 76466 44100 76468
rect 43820 76414 43822 76466
rect 43874 76414 44100 76466
rect 43820 76412 44100 76414
rect 43820 76402 43876 76412
rect 44044 75794 44100 76412
rect 46396 76356 46452 79200
rect 46620 76356 46676 76366
rect 46396 76354 46676 76356
rect 46396 76302 46622 76354
rect 46674 76302 46676 76354
rect 46396 76300 46676 76302
rect 46620 76290 46676 76300
rect 44044 75742 44046 75794
rect 44098 75742 44100 75794
rect 44044 75730 44100 75742
rect 40236 48078 40238 48130
rect 40290 48078 40292 48130
rect 40236 48066 40292 48078
rect 41020 55412 41300 55468
rect 43484 55412 43652 55468
rect 44380 70532 44436 70542
rect 41020 44994 41076 55412
rect 43372 48132 43428 48142
rect 43372 48038 43428 48076
rect 42924 47012 42980 47022
rect 42924 46562 42980 46956
rect 43372 46900 43428 46910
rect 43484 46900 43540 55412
rect 43820 48468 43876 48478
rect 44380 48468 44436 70476
rect 47068 67228 47124 79200
rect 47740 76692 47796 79200
rect 47964 76692 48020 76702
rect 47740 76690 48020 76692
rect 47740 76638 47966 76690
rect 48018 76638 48020 76690
rect 47740 76636 48020 76638
rect 47964 76626 48020 76636
rect 47740 76468 47796 76478
rect 47740 76374 47796 76412
rect 48412 76468 48468 79200
rect 48412 76402 48468 76412
rect 48636 76578 48692 76590
rect 48636 76526 48638 76578
rect 48690 76526 48692 76578
rect 48636 70532 48692 76526
rect 48860 76468 48916 76478
rect 48860 76374 48916 76412
rect 49084 76356 49140 79200
rect 49756 76692 49812 79200
rect 49756 76626 49812 76636
rect 50316 76578 50372 76590
rect 50316 76526 50318 76578
rect 50370 76526 50372 76578
rect 49308 76356 49364 76366
rect 49084 76354 49364 76356
rect 49084 76302 49310 76354
rect 49362 76302 49364 76354
rect 49084 76300 49364 76302
rect 49308 76290 49364 76300
rect 50092 76356 50148 76366
rect 48636 70466 48692 70476
rect 47068 67172 47236 67228
rect 43820 48466 44436 48468
rect 43820 48414 43822 48466
rect 43874 48414 44382 48466
rect 44434 48414 44436 48466
rect 43820 48412 44436 48414
rect 43820 48402 43876 48412
rect 44380 48402 44436 48412
rect 43932 46900 43988 46910
rect 43372 46898 43988 46900
rect 43372 46846 43374 46898
rect 43426 46846 43934 46898
rect 43986 46846 43988 46898
rect 43372 46844 43988 46846
rect 43372 46834 43428 46844
rect 43932 46834 43988 46844
rect 46508 46900 46564 46910
rect 46508 46674 46564 46844
rect 47180 46900 47236 67172
rect 50092 47012 50148 76300
rect 50092 46946 50148 46956
rect 47180 46806 47236 46844
rect 46732 46788 46788 46798
rect 46732 46694 46788 46732
rect 46508 46622 46510 46674
rect 46562 46622 46564 46674
rect 46508 46610 46564 46622
rect 42924 46510 42926 46562
rect 42978 46510 42980 46562
rect 42924 46498 42980 46510
rect 45164 46564 45220 46574
rect 41468 45108 41524 45118
rect 41468 45014 41524 45052
rect 42028 45108 42084 45118
rect 42028 45014 42084 45052
rect 41020 44942 41022 44994
rect 41074 44942 41076 44994
rect 41020 44930 41076 44942
rect 45164 44994 45220 46508
rect 45612 45332 45668 45342
rect 45612 45238 45668 45276
rect 46172 45332 46228 45342
rect 46172 45238 46228 45276
rect 50316 45332 50372 76526
rect 50428 76468 50484 79200
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 50540 76468 50596 76478
rect 50428 76466 50932 76468
rect 50428 76414 50542 76466
rect 50594 76414 50932 76466
rect 50428 76412 50932 76414
rect 50540 76402 50596 76412
rect 50876 75794 50932 76412
rect 50876 75742 50878 75794
rect 50930 75742 50932 75794
rect 50876 75730 50932 75742
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 51100 75124 51156 79200
rect 51212 76466 51268 76478
rect 51212 76414 51214 76466
rect 51266 76414 51268 76466
rect 51212 76356 51268 76414
rect 51212 76290 51268 76300
rect 51772 75796 51828 79200
rect 52220 76692 52276 76702
rect 52220 76598 52276 76636
rect 51772 75730 51828 75740
rect 51660 75684 51716 75694
rect 51100 75058 51156 75068
rect 51548 75628 51660 75684
rect 51324 74898 51380 74910
rect 51324 74846 51326 74898
rect 51378 74846 51380 74898
rect 51100 74788 51156 74798
rect 51324 74788 51380 74846
rect 51100 74786 51380 74788
rect 51100 74734 51102 74786
rect 51154 74734 51380 74786
rect 51100 74732 51380 74734
rect 51100 74722 51156 74732
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50316 45266 50372 45276
rect 45164 44942 45166 44994
rect 45218 44942 45220 44994
rect 45164 44930 45220 44942
rect 42700 44548 42756 44558
rect 42700 44434 42756 44492
rect 42700 44382 42702 44434
rect 42754 44382 42756 44434
rect 42700 44370 42756 44382
rect 44940 44436 44996 44446
rect 44940 44342 44996 44380
rect 51324 44436 51380 74732
rect 51548 44548 51604 75628
rect 51660 75590 51716 75628
rect 52108 75572 52164 75582
rect 52444 75572 52500 79200
rect 53116 77252 53172 79200
rect 53116 77186 53172 77196
rect 53788 77026 53844 79200
rect 54460 77250 54516 79200
rect 54460 77198 54462 77250
rect 54514 77198 54516 77250
rect 54460 77186 54516 77198
rect 53788 76974 53790 77026
rect 53842 76974 53844 77026
rect 53788 76962 53844 76974
rect 54460 77026 54516 77038
rect 54460 76974 54462 77026
rect 54514 76974 54516 77026
rect 54460 76692 54516 76974
rect 54348 76690 54516 76692
rect 54348 76638 54462 76690
rect 54514 76638 54516 76690
rect 54348 76636 54516 76638
rect 54124 76578 54180 76590
rect 54124 76526 54126 76578
rect 54178 76526 54180 76578
rect 53788 75796 53844 75806
rect 53788 75702 53844 75740
rect 52668 75684 52724 75694
rect 52668 75590 52724 75628
rect 52108 75570 52500 75572
rect 52108 75518 52110 75570
rect 52162 75518 52500 75570
rect 52108 75516 52500 75518
rect 52108 75506 52164 75516
rect 52332 75124 52388 75134
rect 52332 75030 52388 75068
rect 51548 44482 51604 44492
rect 51324 44370 51380 44380
rect 43148 44212 43204 44222
rect 43148 44118 43204 44156
rect 43596 44212 43652 44222
rect 43596 44118 43652 44156
rect 45388 44100 45444 44110
rect 45388 44006 45444 44044
rect 45836 44100 45892 44110
rect 45836 44006 45892 44044
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 45836 42756 45892 42766
rect 45836 42662 45892 42700
rect 46396 42532 46452 42542
rect 46396 42438 46452 42476
rect 46844 42532 46900 42542
rect 46844 42438 46900 42476
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 38892 41918 38894 41970
rect 38946 41918 38948 41970
rect 38892 41906 38948 41918
rect 45388 41972 45444 41982
rect 45388 41878 45444 41916
rect 45948 41972 46004 41982
rect 45948 41878 46004 41916
rect 54124 41972 54180 76526
rect 54348 75122 54404 76636
rect 54460 76626 54516 76636
rect 55132 76692 55188 79200
rect 55244 77250 55300 77262
rect 55244 77198 55246 77250
rect 55298 77198 55300 77250
rect 55244 76692 55300 77198
rect 55692 77252 55748 77262
rect 55356 76692 55412 76702
rect 55244 76690 55636 76692
rect 55244 76638 55358 76690
rect 55410 76638 55636 76690
rect 55244 76636 55636 76638
rect 55132 76626 55188 76636
rect 55356 76598 55412 76636
rect 54348 75070 54350 75122
rect 54402 75070 54404 75122
rect 54348 75058 54404 75070
rect 55020 76578 55076 76590
rect 55020 76526 55022 76578
rect 55074 76526 55076 76578
rect 55020 44212 55076 76526
rect 55580 75796 55636 76636
rect 55692 76690 55748 77196
rect 55692 76638 55694 76690
rect 55746 76638 55748 76690
rect 55692 76626 55748 76638
rect 55692 75796 55748 75806
rect 55580 75794 55748 75796
rect 55580 75742 55694 75794
rect 55746 75742 55748 75794
rect 55580 75740 55748 75742
rect 55692 75730 55748 75740
rect 55804 75572 55860 79200
rect 56476 77026 56532 79200
rect 56476 76974 56478 77026
rect 56530 76974 56532 77026
rect 56476 76962 56532 76974
rect 57036 77026 57092 77038
rect 57036 76974 57038 77026
rect 57090 76974 57092 77026
rect 56140 76692 56196 76702
rect 57036 76692 57092 76974
rect 56140 76598 56196 76636
rect 56812 76690 57092 76692
rect 56812 76638 57038 76690
rect 57090 76638 57092 76690
rect 56812 76636 57092 76638
rect 57148 76692 57204 79200
rect 57372 76692 57428 76702
rect 57148 76690 57428 76692
rect 57148 76638 57374 76690
rect 57426 76638 57428 76690
rect 57148 76636 57428 76638
rect 57820 76692 57876 79200
rect 58044 76692 58100 76702
rect 57820 76690 58100 76692
rect 57820 76638 58046 76690
rect 58098 76638 58100 76690
rect 57820 76636 58100 76638
rect 56700 76580 56756 76590
rect 56588 76578 56756 76580
rect 56588 76526 56702 76578
rect 56754 76526 56756 76578
rect 56588 76524 56756 76526
rect 56028 75572 56084 75582
rect 55804 75570 56084 75572
rect 55804 75518 56030 75570
rect 56082 75518 56084 75570
rect 55804 75516 56084 75518
rect 56028 75506 56084 75516
rect 56588 45108 56644 76524
rect 56700 76514 56756 76524
rect 56700 75796 56756 75806
rect 56812 75796 56868 76636
rect 57036 76626 57092 76636
rect 57372 76626 57428 76636
rect 58044 76626 58100 76636
rect 58492 76692 58548 79200
rect 58492 76626 58548 76636
rect 59836 76692 59892 76702
rect 59836 76598 59892 76636
rect 56700 75794 56868 75796
rect 56700 75742 56702 75794
rect 56754 75742 56868 75794
rect 56700 75740 56868 75742
rect 58828 76466 58884 76478
rect 58828 76414 58830 76466
rect 58882 76414 58884 76466
rect 56700 75730 56756 75740
rect 58492 75684 58548 75694
rect 58828 75684 58884 76414
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 58492 75682 58884 75684
rect 58492 75630 58494 75682
rect 58546 75630 58884 75682
rect 58492 75628 58884 75630
rect 58492 48132 58548 75628
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 78204 59330 78260 59342
rect 78204 59278 78206 59330
rect 78258 59278 78260 59330
rect 77980 59218 78036 59230
rect 77980 59166 77982 59218
rect 78034 59166 78036 59218
rect 77532 59108 77588 59118
rect 77980 59108 78036 59166
rect 77532 59106 78036 59108
rect 77532 59054 77534 59106
rect 77586 59054 78036 59106
rect 77532 59052 78036 59054
rect 77532 59042 77588 59052
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 77868 57876 77924 57886
rect 75628 57650 75684 57662
rect 75628 57598 75630 57650
rect 75682 57598 75684 57650
rect 75404 57540 75460 57550
rect 75628 57540 75684 57598
rect 75404 57538 75684 57540
rect 75404 57486 75406 57538
rect 75458 57486 75684 57538
rect 75404 57484 75684 57486
rect 77868 57538 77924 57820
rect 77868 57486 77870 57538
rect 77922 57486 77924 57538
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 75404 55468 75460 57484
rect 77868 57474 77924 57486
rect 77644 56642 77700 56654
rect 77644 56590 77646 56642
rect 77698 56590 77700 56642
rect 77644 56532 77700 56590
rect 77644 56466 77700 56476
rect 77868 56642 77924 56654
rect 77868 56590 77870 56642
rect 77922 56590 77924 56642
rect 77868 55468 77924 56590
rect 75068 55412 75460 55468
rect 77532 55412 77924 55468
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 58492 48066 58548 48076
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 56588 45042 56644 45052
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 55020 44146 55076 44156
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 75068 42756 75124 55412
rect 75628 54514 75684 54526
rect 75628 54462 75630 54514
rect 75682 54462 75684 54514
rect 75404 54404 75460 54414
rect 75628 54404 75684 54462
rect 75068 42690 75124 42700
rect 75292 54402 75684 54404
rect 75292 54350 75406 54402
rect 75458 54350 75684 54402
rect 75292 54348 75684 54350
rect 54124 41906 54180 41916
rect 34412 41860 34468 41870
rect 34412 41298 34468 41804
rect 44940 41860 44996 41870
rect 44940 41766 44996 41804
rect 75292 41860 75348 54348
rect 75404 54338 75460 54348
rect 75628 46674 75684 46686
rect 75628 46622 75630 46674
rect 75682 46622 75684 46674
rect 75404 46564 75460 46574
rect 75628 46564 75684 46622
rect 75460 46508 75684 46564
rect 75404 46470 75460 46508
rect 77532 44100 77588 55412
rect 77756 55188 77812 55198
rect 77756 55094 77812 55132
rect 77868 54402 77924 54414
rect 77868 54350 77870 54402
rect 77922 54350 77924 54402
rect 77868 53844 77924 54350
rect 77868 53778 77924 53788
rect 77868 51490 77924 51502
rect 77868 51438 77870 51490
rect 77922 51438 77924 51490
rect 77644 51266 77700 51278
rect 77644 51214 77646 51266
rect 77698 51214 77700 51266
rect 77644 51156 77700 51214
rect 77644 51090 77700 51100
rect 77756 50372 77812 50382
rect 77756 50278 77812 50316
rect 77868 47572 77924 51438
rect 77532 44034 77588 44044
rect 77644 47516 77924 47572
rect 77644 42532 77700 47516
rect 77868 47012 77924 47022
rect 77868 46562 77924 46956
rect 77980 46788 78036 59052
rect 78204 58884 78260 59278
rect 78204 58818 78260 58828
rect 78204 58546 78260 58558
rect 78204 58494 78206 58546
rect 78258 58494 78260 58546
rect 78204 57204 78260 58494
rect 78204 57138 78260 57148
rect 78204 56642 78260 56654
rect 78204 56590 78206 56642
rect 78258 56590 78260 56642
rect 78204 56532 78260 56590
rect 78204 56466 78260 56476
rect 78204 56194 78260 56206
rect 78204 56142 78206 56194
rect 78258 56142 78260 56194
rect 78204 55860 78260 56142
rect 78204 55794 78260 55804
rect 78204 55074 78260 55086
rect 78204 55022 78206 55074
rect 78258 55022 78260 55074
rect 78204 54516 78260 55022
rect 78204 54450 78260 54460
rect 78204 53842 78260 53854
rect 78204 53790 78206 53842
rect 78258 53790 78260 53842
rect 78204 53172 78260 53790
rect 78204 53106 78260 53116
rect 78204 52722 78260 52734
rect 78204 52670 78206 52722
rect 78258 52670 78260 52722
rect 78204 52500 78260 52670
rect 78204 52434 78260 52444
rect 78204 51938 78260 51950
rect 78204 51886 78206 51938
rect 78258 51886 78260 51938
rect 78204 51828 78260 51886
rect 78204 51762 78260 51772
rect 78204 51378 78260 51390
rect 78204 51326 78206 51378
rect 78258 51326 78260 51378
rect 78204 51156 78260 51326
rect 78204 51090 78260 51100
rect 78204 50372 78260 50382
rect 78204 50370 78372 50372
rect 78204 50318 78206 50370
rect 78258 50318 78372 50370
rect 78204 50316 78372 50318
rect 78204 50306 78260 50316
rect 78204 49922 78260 49934
rect 78204 49870 78206 49922
rect 78258 49870 78260 49922
rect 78204 49140 78260 49870
rect 78316 49812 78372 50316
rect 78428 49812 78484 49822
rect 78316 49756 78428 49812
rect 78428 49746 78484 49756
rect 78204 49074 78260 49084
rect 78204 48804 78260 48814
rect 78204 48710 78260 48748
rect 78204 48354 78260 48366
rect 78204 48302 78206 48354
rect 78258 48302 78260 48354
rect 78204 47796 78260 48302
rect 78204 47730 78260 47740
rect 77980 46722 78036 46732
rect 78204 47234 78260 47246
rect 78204 47182 78206 47234
rect 78258 47182 78260 47234
rect 77868 46510 77870 46562
rect 77922 46510 77924 46562
rect 77868 46498 77924 46510
rect 78204 46452 78260 47182
rect 78204 46386 78260 46396
rect 77756 45780 77812 45790
rect 77756 45686 77812 45724
rect 78204 45666 78260 45678
rect 78204 45614 78206 45666
rect 78258 45614 78260 45666
rect 78204 45444 78260 45614
rect 78204 45378 78260 45388
rect 78204 45218 78260 45230
rect 78204 45166 78206 45218
rect 78258 45166 78260 45218
rect 78204 44436 78260 45166
rect 78204 44370 78260 44380
rect 78204 44100 78260 44110
rect 78204 44098 78372 44100
rect 78204 44046 78206 44098
rect 78258 44046 78372 44098
rect 78204 44044 78372 44046
rect 78204 44034 78260 44044
rect 78204 43762 78260 43774
rect 78204 43710 78206 43762
rect 78258 43710 78260 43762
rect 78204 43092 78260 43710
rect 78316 43764 78372 44044
rect 78428 43764 78484 43774
rect 78316 43708 78428 43764
rect 78428 43698 78484 43708
rect 78204 43026 78260 43036
rect 77644 42466 77700 42476
rect 78204 42530 78260 42542
rect 78204 42478 78206 42530
rect 78258 42478 78260 42530
rect 78204 42420 78260 42478
rect 78204 42354 78260 42364
rect 75292 41794 75348 41804
rect 78204 42082 78260 42094
rect 78204 42030 78206 42082
rect 78258 42030 78260 42082
rect 78204 41748 78260 42030
rect 78204 41682 78260 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 34412 41246 34414 41298
rect 34466 41246 34468 41298
rect 34412 41234 34468 41246
rect 78204 41076 78260 41086
rect 78204 40982 78260 41020
rect 33628 40964 33684 40974
rect 33964 40964 34020 40974
rect 33684 40962 34020 40964
rect 33684 40910 33966 40962
rect 34018 40910 34020 40962
rect 33684 40908 34020 40910
rect 33628 40870 33684 40908
rect 33964 40898 34020 40908
rect 77756 40962 77812 40974
rect 77756 40910 77758 40962
rect 77810 40910 77812 40962
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 4956 40450 5012 40460
rect 35084 40516 35140 40526
rect 35140 40460 35252 40516
rect 35084 40450 35140 40460
rect 2380 40338 2436 40348
rect 34412 40404 34468 40414
rect 34636 40404 34692 40414
rect 34468 40402 34692 40404
rect 34468 40350 34638 40402
rect 34690 40350 34692 40402
rect 34468 40348 34692 40350
rect 34412 40310 34468 40348
rect 34636 40338 34692 40348
rect 35196 40402 35252 40460
rect 35196 40350 35198 40402
rect 35250 40350 35252 40402
rect 35196 40338 35252 40350
rect 77756 40404 77812 40910
rect 77756 40338 77812 40348
rect 78204 40514 78260 40526
rect 78204 40462 78206 40514
rect 78258 40462 78260 40514
rect 1708 40178 1764 40190
rect 1708 40126 1710 40178
rect 1762 40126 1764 40178
rect 1708 39732 1764 40126
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 78204 39956 78260 40462
rect 78204 39890 78260 39900
rect 1708 39666 1764 39676
rect 40348 39730 40404 39742
rect 40348 39678 40350 39730
rect 40402 39678 40404 39730
rect 1708 39394 1764 39406
rect 1708 39342 1710 39394
rect 1762 39342 1764 39394
rect 1708 39060 1764 39342
rect 40012 39396 40068 39406
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 1708 38994 1764 39004
rect 2044 38948 2100 38958
rect 2044 38854 2100 38892
rect 40012 38948 40068 39340
rect 40012 38882 40068 38892
rect 1708 38834 1764 38846
rect 1708 38782 1710 38834
rect 1762 38782 1764 38834
rect 1708 38388 1764 38782
rect 35308 38834 35364 38846
rect 35308 38782 35310 38834
rect 35362 38782 35364 38834
rect 1708 38322 1764 38332
rect 2492 38722 2548 38734
rect 34972 38724 35028 38734
rect 35308 38724 35364 38782
rect 38332 38834 38388 38846
rect 38332 38782 38334 38834
rect 38386 38782 38388 38834
rect 2492 38670 2494 38722
rect 2546 38670 2548 38722
rect 2492 38388 2548 38670
rect 34860 38722 35364 38724
rect 34860 38670 34974 38722
rect 35026 38670 35364 38722
rect 34860 38668 35364 38670
rect 35868 38722 35924 38734
rect 35868 38670 35870 38722
rect 35922 38670 35924 38722
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 2492 38322 2548 38332
rect 33404 38050 33460 38062
rect 33404 37998 33406 38050
rect 33458 37998 33460 38050
rect 1708 37828 1764 37838
rect 1708 37734 1764 37772
rect 32620 37828 32676 37838
rect 32844 37828 32900 37838
rect 32620 37826 32900 37828
rect 32620 37774 32622 37826
rect 32674 37774 32846 37826
rect 32898 37774 32900 37826
rect 32620 37772 32900 37774
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 2044 37380 2100 37390
rect 2044 37286 2100 37324
rect 1708 37266 1764 37278
rect 1708 37214 1710 37266
rect 1762 37214 1764 37266
rect 1708 37044 1764 37214
rect 1708 36978 1764 36988
rect 2044 37156 2100 37166
rect 1708 36372 1764 36382
rect 1708 36278 1764 36316
rect 2044 36370 2100 37100
rect 2492 37154 2548 37166
rect 2492 37102 2494 37154
rect 2546 37102 2548 37154
rect 2492 37044 2548 37102
rect 2492 36978 2548 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 2044 36318 2046 36370
rect 2098 36318 2100 36370
rect 2044 36306 2100 36318
rect 2940 36372 2996 36382
rect 2940 36278 2996 36316
rect 2380 36258 2436 36270
rect 2380 36206 2382 36258
rect 2434 36206 2436 36258
rect 1708 35810 1764 35822
rect 1708 35758 1710 35810
rect 1762 35758 1764 35810
rect 1708 35028 1764 35758
rect 2380 35700 2436 36206
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 2380 35634 2436 35644
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 1708 34962 1764 34972
rect 1820 34914 1876 34926
rect 1820 34862 1822 34914
rect 1874 34862 1876 34914
rect 1820 34356 1876 34862
rect 2044 34692 2100 34702
rect 2044 34598 2100 34636
rect 2492 34690 2548 34702
rect 2492 34638 2494 34690
rect 2546 34638 2548 34690
rect 1820 34290 1876 34300
rect 2492 34356 2548 34638
rect 32620 34692 32676 37772
rect 32844 37762 32900 37772
rect 32620 34626 32676 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 2492 34290 2548 34300
rect 1708 34242 1764 34254
rect 1708 34190 1710 34242
rect 1762 34190 1764 34242
rect 1708 33684 1764 34190
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 1708 33618 1764 33628
rect 1708 33458 1764 33470
rect 1708 33406 1710 33458
rect 1762 33406 1764 33458
rect 1708 33012 1764 33406
rect 1708 32946 1764 32956
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 2044 32676 2100 32686
rect 2044 32582 2100 32620
rect 1708 32562 1764 32574
rect 1708 32510 1710 32562
rect 1762 32510 1764 32562
rect 1708 32340 1764 32510
rect 1708 32274 1764 32284
rect 2492 32450 2548 32462
rect 2492 32398 2494 32450
rect 2546 32398 2548 32450
rect 2492 32340 2548 32398
rect 2492 32274 2548 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 1932 31890 1988 31902
rect 1932 31838 1934 31890
rect 1986 31838 1988 31890
rect 1708 31668 1764 31678
rect 1708 31220 1764 31612
rect 1708 31106 1764 31164
rect 1708 31054 1710 31106
rect 1762 31054 1764 31106
rect 1708 31042 1764 31054
rect 1932 30996 1988 31838
rect 4284 31780 4340 31790
rect 4284 31686 4340 31724
rect 4844 31780 4900 31790
rect 4844 31686 4900 31724
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 2940 31220 2996 31230
rect 2940 31126 2996 31164
rect 2044 31108 2100 31118
rect 2044 31014 2100 31052
rect 1932 30930 1988 30940
rect 2380 30770 2436 30782
rect 2380 30718 2382 30770
rect 2434 30718 2436 30770
rect 2380 30324 2436 30718
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 2380 30258 2436 30268
rect 4284 30210 4340 30222
rect 4284 30158 4286 30210
rect 4338 30158 4340 30210
rect 2492 30098 2548 30110
rect 2492 30046 2494 30098
rect 2546 30046 2548 30098
rect 2492 29652 2548 30046
rect 4284 29988 4340 30158
rect 4284 29922 4340 29932
rect 4844 29988 4900 29998
rect 4844 29894 4900 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 2492 29586 2548 29596
rect 1708 29204 1764 29214
rect 1708 29110 1764 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 1932 28754 1988 28766
rect 1932 28702 1934 28754
rect 1986 28702 1988 28754
rect 1932 28308 1988 28702
rect 4284 28644 4340 28654
rect 4284 28550 4340 28588
rect 4844 28644 4900 28654
rect 4844 28550 4900 28588
rect 1932 28242 1988 28252
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 1708 27970 1764 27982
rect 1708 27918 1710 27970
rect 1762 27918 1764 27970
rect 1708 27636 1764 27918
rect 1708 27570 1764 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1708 26964 1764 26974
rect 1708 26850 1764 26908
rect 1708 26798 1710 26850
rect 1762 26798 1764 26850
rect 1708 26786 1764 26798
rect 2156 26850 2212 26862
rect 2156 26798 2158 26850
rect 2210 26798 2212 26850
rect 1708 26402 1764 26414
rect 1708 26350 1710 26402
rect 1762 26350 1764 26402
rect 1708 25620 1764 26350
rect 2156 26292 2212 26798
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 2156 26226 2212 26236
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 1708 25554 1764 25564
rect 1708 25282 1764 25294
rect 1708 25230 1710 25282
rect 1762 25230 1764 25282
rect 1708 25060 1764 25230
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 1708 24994 1764 25004
rect 1708 24834 1764 24846
rect 1708 24782 1710 24834
rect 1762 24782 1764 24834
rect 1708 24276 1764 24782
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 1708 24210 1764 24220
rect 1708 23716 1764 23726
rect 1708 23622 1764 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 1708 23266 1764 23278
rect 1708 23214 1710 23266
rect 1762 23214 1764 23266
rect 1708 22932 1764 23214
rect 1708 22866 1764 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 1932 22482 1988 22494
rect 1932 22430 1934 22482
rect 1986 22430 1988 22482
rect 1708 22260 1764 22270
rect 1708 21810 1764 22204
rect 1708 21758 1710 21810
rect 1762 21758 1764 21810
rect 1708 21746 1764 21758
rect 1932 21588 1988 22430
rect 4284 22372 4340 22382
rect 4284 22278 4340 22316
rect 4844 22372 4900 22382
rect 4844 22278 4900 22316
rect 2940 22260 2996 22270
rect 2940 21810 2996 22204
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 2940 21758 2942 21810
rect 2994 21758 2996 21810
rect 2940 21746 2996 21758
rect 2044 21700 2100 21710
rect 2044 21606 2100 21644
rect 2380 21698 2436 21710
rect 2380 21646 2382 21698
rect 2434 21646 2436 21698
rect 1932 21522 1988 21532
rect 2380 20916 2436 21646
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 2380 20850 2436 20860
rect 1708 20578 1764 20590
rect 1708 20526 1710 20578
rect 1762 20526 1764 20578
rect 1708 20244 1764 20526
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 1708 20178 1764 20188
rect 2044 20132 2100 20142
rect 2044 20038 2100 20076
rect 1708 20018 1764 20030
rect 1708 19966 1710 20018
rect 1762 19966 1764 20018
rect 1708 19572 1764 19966
rect 1708 19506 1764 19516
rect 2492 19906 2548 19918
rect 2492 19854 2494 19906
rect 2546 19854 2548 19906
rect 2492 19572 2548 19854
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 2492 19506 2548 19516
rect 1708 19012 1764 19022
rect 1708 18918 1764 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 1708 18562 1764 18574
rect 1708 18510 1710 18562
rect 1762 18510 1764 18562
rect 1708 18228 1764 18510
rect 1708 18162 1764 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17778 1988 17790
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1708 17556 1764 17566
rect 1708 17108 1764 17500
rect 1708 17014 1764 17052
rect 1932 16884 1988 17726
rect 4284 17666 4340 17678
rect 4284 17614 4286 17666
rect 4338 17614 4340 17666
rect 4284 17444 4340 17614
rect 4284 17378 4340 17388
rect 4844 17444 4900 17454
rect 4844 17350 4900 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 2940 17108 2996 17118
rect 2940 17014 2996 17052
rect 1932 16818 1988 16828
rect 2044 16994 2100 17006
rect 2044 16942 2046 16994
rect 2098 16942 2100 16994
rect 2044 16772 2100 16942
rect 2044 16706 2100 16716
rect 2380 16994 2436 17006
rect 2380 16942 2382 16994
rect 2434 16942 2436 16994
rect 2380 16212 2436 16942
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 2380 16146 2436 16156
rect 1708 15876 1764 15886
rect 1708 15782 1764 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 1708 15426 1764 15438
rect 1708 15374 1710 15426
rect 1762 15374 1764 15426
rect 1708 14868 1764 15374
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 1708 14802 1764 14812
rect 1708 14308 1764 14318
rect 1708 14214 1764 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 1708 13524 1764 13534
rect 1708 13430 1764 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 1932 13074 1988 13086
rect 1932 13022 1934 13074
rect 1986 13022 1988 13074
rect 1708 12852 1764 12862
rect 1708 12402 1764 12796
rect 1708 12350 1710 12402
rect 1762 12350 1764 12402
rect 1708 12338 1764 12350
rect 1932 12180 1988 13022
rect 4284 12962 4340 12974
rect 4284 12910 4286 12962
rect 4338 12910 4340 12962
rect 4284 12740 4340 12910
rect 4284 12674 4340 12684
rect 4844 12740 4900 12750
rect 4844 12646 4900 12684
rect 33404 12740 33460 37998
rect 33852 37266 33908 37278
rect 33852 37214 33854 37266
rect 33906 37214 33908 37266
rect 33516 37156 33572 37166
rect 33852 37156 33908 37214
rect 33572 37100 33908 37156
rect 34412 37156 34468 37166
rect 34412 37154 34580 37156
rect 34412 37102 34414 37154
rect 34466 37102 34580 37154
rect 34412 37100 34580 37102
rect 33516 37062 33572 37100
rect 34412 37090 34468 37100
rect 34188 36260 34244 36270
rect 34412 36260 34468 36270
rect 34188 36258 34468 36260
rect 34188 36206 34190 36258
rect 34242 36206 34414 36258
rect 34466 36206 34468 36258
rect 34188 36204 34468 36206
rect 34188 35812 34244 36204
rect 34412 36194 34468 36204
rect 33964 35756 34244 35812
rect 33628 35588 33684 35598
rect 33852 35588 33908 35598
rect 33628 35586 33908 35588
rect 33628 35534 33630 35586
rect 33682 35534 33854 35586
rect 33906 35534 33908 35586
rect 33628 35532 33908 35534
rect 33628 21700 33684 35532
rect 33852 35522 33908 35532
rect 33964 31108 34020 35756
rect 33964 31042 34020 31052
rect 34076 35586 34132 35598
rect 34076 35534 34078 35586
rect 34130 35534 34132 35586
rect 34076 22372 34132 35534
rect 34188 34132 34244 34142
rect 34188 34038 34244 34076
rect 34524 33908 34580 37100
rect 34076 22306 34132 22316
rect 34412 33852 34580 33908
rect 34636 34132 34692 34142
rect 33628 21634 33684 21644
rect 34412 17444 34468 33852
rect 34636 31948 34692 34076
rect 34860 32676 34916 38668
rect 34972 38658 35028 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 34860 32610 34916 32620
rect 34972 36482 35028 36494
rect 34972 36430 34974 36482
rect 35026 36430 35028 36482
rect 34524 31892 34692 31948
rect 34524 20132 34580 31892
rect 34972 31780 35028 36430
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34972 31714 35028 31724
rect 35084 34018 35140 34030
rect 35084 33966 35086 34018
rect 35138 33966 35140 34018
rect 34524 20066 34580 20076
rect 34412 17378 34468 17388
rect 33404 12674 33460 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 1932 12114 1988 12124
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35084 6804 35140 33966
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35868 29988 35924 38670
rect 37996 38724 38052 38734
rect 38332 38724 38388 38782
rect 39228 38834 39284 38846
rect 39228 38782 39230 38834
rect 39282 38782 39284 38834
rect 37996 38722 38388 38724
rect 37996 38670 37998 38722
rect 38050 38670 38388 38722
rect 37996 38668 38388 38670
rect 37996 38658 38052 38668
rect 35868 29922 35924 29932
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35084 6738 35140 6748
rect 35980 6804 36036 6814
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 35980 4564 36036 6748
rect 36876 4564 36932 4574
rect 35980 4562 36932 4564
rect 35980 4510 36878 4562
rect 36930 4510 36932 4562
rect 35980 4508 36932 4510
rect 29596 4338 29652 4350
rect 29596 4286 29598 4338
rect 29650 4286 29652 4338
rect 29596 4228 29652 4286
rect 35980 4338 36036 4508
rect 36876 4498 36932 4508
rect 35980 4286 35982 4338
rect 36034 4286 36036 4338
rect 35980 4274 36036 4286
rect 29596 4162 29652 4172
rect 30156 4228 30212 4238
rect 30156 4134 30212 4172
rect 27356 4116 27412 4126
rect 34076 4116 34132 4126
rect 26908 4114 27412 4116
rect 26908 4062 27358 4114
rect 27410 4062 27412 4114
rect 26908 4060 27412 4062
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 26796 3444 26852 3454
rect 26796 3350 26852 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 26908 800 26964 4060
rect 27356 4050 27412 4060
rect 33628 4114 34132 4116
rect 33628 4062 34078 4114
rect 34130 4062 34132 4114
rect 33628 4060 34132 4062
rect 29148 3668 29204 3678
rect 29820 3668 29876 3678
rect 30492 3668 30548 3678
rect 28924 3666 29204 3668
rect 28924 3614 29150 3666
rect 29202 3614 29204 3666
rect 28924 3612 29204 3614
rect 27244 3556 27300 3566
rect 27244 3462 27300 3500
rect 27580 3554 27636 3566
rect 27580 3502 27582 3554
rect 27634 3502 27636 3554
rect 27580 3444 27636 3502
rect 28252 3556 28308 3566
rect 27580 800 27636 3388
rect 27804 3444 27860 3454
rect 27804 3350 27860 3388
rect 28252 3444 28308 3500
rect 28812 3556 28868 3566
rect 28476 3444 28532 3454
rect 28252 3442 28532 3444
rect 28252 3390 28478 3442
rect 28530 3390 28532 3442
rect 28252 3388 28532 3390
rect 28252 800 28308 3388
rect 28476 3378 28532 3388
rect 28812 3442 28868 3500
rect 28812 3390 28814 3442
rect 28866 3390 28868 3442
rect 28812 3378 28868 3390
rect 28924 800 28980 3612
rect 29148 3602 29204 3612
rect 29596 3666 29876 3668
rect 29596 3614 29822 3666
rect 29874 3614 29876 3666
rect 29596 3612 29876 3614
rect 29596 800 29652 3612
rect 29820 3602 29876 3612
rect 30268 3666 30548 3668
rect 30268 3614 30494 3666
rect 30546 3614 30548 3666
rect 30268 3612 30548 3614
rect 30268 800 30324 3612
rect 30492 3602 30548 3612
rect 31612 3666 31668 3678
rect 31612 3614 31614 3666
rect 31666 3614 31668 3666
rect 31052 3332 31108 3342
rect 30940 3330 31108 3332
rect 30940 3278 31054 3330
rect 31106 3278 31108 3330
rect 30940 3276 31108 3278
rect 30940 800 30996 3276
rect 31052 3266 31108 3276
rect 31612 800 31668 3614
rect 32508 3332 32564 3342
rect 33180 3332 33236 3342
rect 32284 3330 32564 3332
rect 32284 3278 32510 3330
rect 32562 3278 32564 3330
rect 32284 3276 32564 3278
rect 32284 800 32340 3276
rect 32508 3266 32564 3276
rect 32956 3330 33236 3332
rect 32956 3278 33182 3330
rect 33234 3278 33236 3330
rect 32956 3276 33236 3278
rect 32956 800 33012 3276
rect 33180 3266 33236 3276
rect 33628 800 33684 4060
rect 34076 4050 34132 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 38332 3556 38388 38668
rect 38780 38722 38836 38734
rect 38780 38670 38782 38722
rect 38834 38670 38836 38722
rect 38780 28644 38836 38670
rect 38780 28578 38836 28588
rect 38892 37828 38948 37838
rect 39228 37828 39284 38782
rect 38892 37826 39284 37828
rect 38892 37774 38894 37826
rect 38946 37774 39284 37826
rect 38892 37772 39284 37774
rect 39788 38722 39844 38734
rect 39788 38670 39790 38722
rect 39842 38670 39844 38722
rect 38332 3490 38388 3500
rect 38892 3444 38948 37772
rect 39564 35586 39620 35598
rect 39564 35534 39566 35586
rect 39618 35534 39620 35586
rect 39564 5236 39620 35534
rect 39564 5170 39620 5180
rect 39788 4228 39844 38670
rect 40124 35698 40180 35710
rect 40124 35646 40126 35698
rect 40178 35646 40180 35698
rect 40124 35588 40180 35646
rect 40124 35522 40180 35532
rect 40348 21476 40404 39678
rect 78204 39730 78260 39742
rect 78204 39678 78206 39730
rect 78258 39678 78260 39730
rect 41692 39618 41748 39630
rect 41692 39566 41694 39618
rect 41746 39566 41748 39618
rect 40796 39396 40852 39406
rect 41132 39396 41188 39406
rect 40796 39394 40964 39396
rect 40796 39342 40798 39394
rect 40850 39342 40964 39394
rect 40796 39340 40964 39342
rect 40796 39330 40852 39340
rect 40908 38724 40964 39340
rect 41132 39302 41188 39340
rect 41020 38724 41076 38734
rect 40908 38722 41076 38724
rect 40908 38670 41022 38722
rect 41074 38670 41076 38722
rect 40908 38668 41076 38670
rect 40348 21410 40404 21420
rect 40460 33346 40516 33358
rect 40460 33294 40462 33346
rect 40514 33294 40516 33346
rect 40460 5684 40516 33294
rect 40908 20580 40964 38668
rect 41020 38658 41076 38668
rect 41020 35588 41076 35598
rect 41020 35494 41076 35532
rect 41020 33124 41076 33134
rect 41580 33124 41636 33134
rect 41020 33122 41636 33124
rect 41020 33070 41022 33122
rect 41074 33070 41582 33122
rect 41634 33070 41636 33122
rect 41020 33068 41636 33070
rect 41020 33058 41076 33068
rect 40908 20514 40964 20524
rect 40460 5618 40516 5628
rect 39788 4162 39844 4172
rect 41132 4226 41188 4238
rect 41132 4174 41134 4226
rect 41186 4174 41188 4226
rect 39900 3668 39956 3678
rect 38892 3378 38948 3388
rect 39676 3666 39956 3668
rect 39676 3614 39902 3666
rect 39954 3614 39956 3666
rect 39676 3612 39956 3614
rect 34524 3332 34580 3342
rect 35196 3332 35252 3342
rect 35980 3332 36036 3342
rect 36540 3332 36596 3342
rect 37212 3332 37268 3342
rect 37884 3332 37940 3342
rect 38556 3332 38612 3342
rect 39116 3332 39172 3342
rect 34300 3330 34580 3332
rect 34300 3278 34526 3330
rect 34578 3278 34580 3330
rect 34300 3276 34580 3278
rect 34300 800 34356 3276
rect 34524 3266 34580 3276
rect 34972 3330 35252 3332
rect 34972 3278 35198 3330
rect 35250 3278 35252 3330
rect 34972 3276 35252 3278
rect 34972 800 35028 3276
rect 35196 3266 35252 3276
rect 35644 3330 36036 3332
rect 35644 3278 35982 3330
rect 36034 3278 36036 3330
rect 35644 3276 36036 3278
rect 35644 800 35700 3276
rect 35980 3266 36036 3276
rect 36316 3330 36596 3332
rect 36316 3278 36542 3330
rect 36594 3278 36596 3330
rect 36316 3276 36596 3278
rect 36316 800 36372 3276
rect 36540 3266 36596 3276
rect 36988 3330 37268 3332
rect 36988 3278 37214 3330
rect 37266 3278 37268 3330
rect 36988 3276 37268 3278
rect 36988 800 37044 3276
rect 37212 3266 37268 3276
rect 37660 3330 37940 3332
rect 37660 3278 37886 3330
rect 37938 3278 37940 3330
rect 37660 3276 37940 3278
rect 37660 800 37716 3276
rect 37884 3266 37940 3276
rect 38332 3330 38612 3332
rect 38332 3278 38558 3330
rect 38610 3278 38612 3330
rect 38332 3276 38612 3278
rect 38332 800 38388 3276
rect 38556 3266 38612 3276
rect 39004 3330 39172 3332
rect 39004 3278 39118 3330
rect 39170 3278 39172 3330
rect 39004 3276 39172 3278
rect 39004 800 39060 3276
rect 39116 3266 39172 3276
rect 39676 800 39732 3612
rect 39900 3602 39956 3612
rect 41132 3444 41188 4174
rect 41244 3444 41300 3454
rect 41020 3442 41300 3444
rect 41020 3390 41246 3442
rect 41298 3390 41300 3442
rect 41020 3388 41300 3390
rect 40572 3332 40628 3342
rect 40348 3330 40628 3332
rect 40348 3278 40574 3330
rect 40626 3278 40628 3330
rect 40348 3276 40628 3278
rect 40348 800 40404 3276
rect 40572 3266 40628 3276
rect 41020 800 41076 3388
rect 41244 3378 41300 3388
rect 41580 3442 41636 33068
rect 41692 23044 41748 39566
rect 44828 39620 44884 39630
rect 44828 39618 45108 39620
rect 44828 39566 44830 39618
rect 44882 39566 45108 39618
rect 44828 39564 45108 39566
rect 44828 39554 44884 39564
rect 44044 38834 44100 38846
rect 44044 38782 44046 38834
rect 44098 38782 44100 38834
rect 43708 38724 43764 38734
rect 44044 38724 44100 38782
rect 43708 38722 44100 38724
rect 43708 38670 43710 38722
rect 43762 38670 44100 38722
rect 43708 38668 44100 38670
rect 44604 38724 44660 38734
rect 44604 38722 44996 38724
rect 44604 38670 44606 38722
rect 44658 38670 44996 38722
rect 44604 38668 44996 38670
rect 43708 37380 43764 38668
rect 44604 38658 44660 38668
rect 43708 37314 43764 37324
rect 43148 35700 43204 35710
rect 41692 22978 41748 22988
rect 41916 35588 41972 35598
rect 41580 3390 41582 3442
rect 41634 3390 41636 3442
rect 41580 3378 41636 3390
rect 41692 4226 41748 4238
rect 41692 4174 41694 4226
rect 41746 4174 41748 4226
rect 41692 3556 41748 4174
rect 41692 800 41748 3500
rect 41916 3442 41972 35532
rect 43148 31948 43204 35644
rect 44156 35700 44212 35710
rect 44156 35606 44212 35644
rect 43596 35586 43652 35598
rect 43596 35534 43598 35586
rect 43650 35534 43652 35586
rect 43036 31892 43204 31948
rect 43484 32450 43540 32462
rect 43484 32398 43486 32450
rect 43538 32398 43540 32450
rect 43036 8428 43092 31892
rect 42924 8372 43092 8428
rect 42476 5684 42532 5694
rect 42476 5124 42532 5628
rect 42476 4562 42532 5068
rect 42476 4510 42478 4562
rect 42530 4510 42532 4562
rect 42476 4498 42532 4510
rect 42812 4114 42868 4126
rect 42812 4062 42814 4114
rect 42866 4062 42868 4114
rect 42364 3668 42420 3678
rect 42140 3556 42196 3566
rect 42140 3462 42196 3500
rect 41916 3390 41918 3442
rect 41970 3390 41972 3442
rect 41916 3378 41972 3390
rect 42364 800 42420 3612
rect 42812 3554 42868 4062
rect 42812 3502 42814 3554
rect 42866 3502 42868 3554
rect 42812 3444 42868 3502
rect 42924 3444 42980 8372
rect 43148 5236 43204 5246
rect 43148 4900 43204 5180
rect 43260 5124 43316 5134
rect 43316 5068 43428 5124
rect 43260 5058 43316 5068
rect 43260 4900 43316 4910
rect 43148 4898 43316 4900
rect 43148 4846 43262 4898
rect 43314 4846 43316 4898
rect 43148 4844 43316 4846
rect 43260 4834 43316 4844
rect 43372 4338 43428 5068
rect 43372 4286 43374 4338
rect 43426 4286 43428 4338
rect 43372 4274 43428 4286
rect 43036 4226 43092 4238
rect 43036 4174 43038 4226
rect 43090 4174 43092 4226
rect 43036 4114 43092 4174
rect 43036 4062 43038 4114
rect 43090 4062 43092 4114
rect 43036 4050 43092 4062
rect 43148 4116 43204 4126
rect 43036 3444 43092 3454
rect 42924 3442 43092 3444
rect 42924 3390 43038 3442
rect 43090 3390 43092 3442
rect 42924 3388 43092 3390
rect 42812 3378 42868 3388
rect 43036 3378 43092 3388
rect 43148 2100 43204 4060
rect 43484 3556 43540 32398
rect 43596 4228 43652 35534
rect 44380 34692 44436 34702
rect 44828 34692 44884 34702
rect 44380 34690 44884 34692
rect 44380 34638 44382 34690
rect 44434 34638 44830 34690
rect 44882 34638 44884 34690
rect 44380 34636 44884 34638
rect 44044 32564 44100 32574
rect 44044 32470 44100 32508
rect 44380 16772 44436 34636
rect 44828 34626 44884 34636
rect 44380 16706 44436 16716
rect 44492 32564 44548 32574
rect 44492 5908 44548 32508
rect 44940 26180 44996 38668
rect 44940 26114 44996 26124
rect 45052 24612 45108 39564
rect 45388 39396 45444 39406
rect 45948 39396 46004 39406
rect 45388 39394 46004 39396
rect 45388 39342 45390 39394
rect 45442 39342 45950 39394
rect 46002 39342 46004 39394
rect 45388 39340 46004 39342
rect 45276 35026 45332 35038
rect 45276 34974 45278 35026
rect 45330 34974 45332 35026
rect 45276 30884 45332 34974
rect 45276 30818 45332 30828
rect 45388 27076 45444 39340
rect 45948 39330 46004 39340
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 78204 39060 78260 39678
rect 78204 38994 78260 39004
rect 78204 38610 78260 38622
rect 78204 38558 78206 38610
rect 78258 38558 78260 38610
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 78204 38388 78260 38558
rect 78204 38322 78260 38332
rect 78204 37826 78260 37838
rect 78204 37774 78206 37826
rect 78258 37774 78260 37826
rect 78204 37716 78260 37774
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 78204 37650 78260 37660
rect 50556 37594 50820 37604
rect 78204 37378 78260 37390
rect 78204 37326 78206 37378
rect 78258 37326 78260 37378
rect 78204 37044 78260 37326
rect 78204 36978 78260 36988
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 77756 36594 77812 36606
rect 77756 36542 77758 36594
rect 77810 36542 77812 36594
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 77756 35700 77812 36542
rect 78204 36372 78260 36382
rect 78204 36278 78260 36316
rect 77756 35634 77812 35644
rect 78204 35474 78260 35486
rect 78204 35422 78206 35474
rect 78258 35422 78260 35474
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 78204 35028 78260 35422
rect 78204 34962 78260 34972
rect 78204 34690 78260 34702
rect 78204 34638 78206 34690
rect 78258 34638 78260 34690
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 78204 34356 78260 34638
rect 78204 34290 78260 34300
rect 77868 34244 77924 34254
rect 77868 34150 77924 34188
rect 46620 34130 46676 34142
rect 46620 34078 46622 34130
rect 46674 34078 46676 34130
rect 45388 27010 45444 27020
rect 46060 34018 46116 34030
rect 46060 33966 46062 34018
rect 46114 33966 46116 34018
rect 45052 24546 45108 24556
rect 46060 19908 46116 33966
rect 46620 34020 46676 34078
rect 78204 34130 78260 34142
rect 78204 34078 78206 34130
rect 78258 34078 78260 34130
rect 46620 33954 46676 33964
rect 47068 34020 47124 34030
rect 47068 33926 47124 33964
rect 77644 34020 77700 34030
rect 78204 34020 78260 34078
rect 77644 34018 78260 34020
rect 77644 33966 77646 34018
rect 77698 33966 78260 34018
rect 77644 33964 78260 33966
rect 77644 33954 77700 33964
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 78204 33684 78260 33964
rect 78204 33618 78260 33628
rect 78204 33122 78260 33134
rect 78204 33070 78206 33122
rect 78258 33070 78260 33122
rect 78204 33012 78260 33070
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 78204 32946 78260 32956
rect 50556 32890 50820 32900
rect 78204 32674 78260 32686
rect 78204 32622 78206 32674
rect 78258 32622 78260 32674
rect 78204 32340 78260 32622
rect 78204 32274 78260 32284
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 77756 32002 77812 32014
rect 77756 31950 77758 32002
rect 77810 31950 77812 32002
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 75628 30994 75684 31006
rect 75628 30942 75630 30994
rect 75682 30942 75684 30994
rect 75292 30884 75348 30894
rect 75628 30884 75684 30942
rect 77756 30996 77812 31950
rect 78204 31668 78260 31678
rect 78204 31574 78260 31612
rect 77756 30930 77812 30940
rect 75348 30828 75684 30884
rect 75292 30790 75348 30828
rect 77980 30770 78036 30782
rect 77980 30718 77982 30770
rect 78034 30718 78036 30770
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 77980 30324 78036 30718
rect 77980 30258 78036 30268
rect 78204 29988 78260 29998
rect 78204 29986 78372 29988
rect 78204 29934 78206 29986
rect 78258 29934 78372 29986
rect 78204 29932 78372 29934
rect 78204 29922 78260 29932
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 78316 29652 78372 29932
rect 78428 29652 78484 29662
rect 78316 29596 78428 29652
rect 78428 29586 78484 29596
rect 78204 29538 78260 29550
rect 78204 29486 78206 29538
rect 78258 29486 78260 29538
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 78204 28980 78260 29486
rect 78204 28914 78260 28924
rect 78204 28418 78260 28430
rect 78204 28366 78206 28418
rect 78258 28366 78260 28418
rect 78204 28308 78260 28366
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 78204 28242 78260 28252
rect 50556 28186 50820 28196
rect 78204 27970 78260 27982
rect 78204 27918 78206 27970
rect 78258 27918 78260 27970
rect 78204 27636 78260 27918
rect 78204 27570 78260 27580
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 77196 27188 77252 27198
rect 77196 27094 77252 27132
rect 78204 27188 78260 27198
rect 77868 27076 77924 27086
rect 77868 26962 77924 27020
rect 77868 26910 77870 26962
rect 77922 26910 77924 26962
rect 77868 26898 77924 26910
rect 78204 26962 78260 27132
rect 78204 26910 78206 26962
rect 78258 26910 78260 26962
rect 77532 26852 77588 26862
rect 77532 26758 77588 26796
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 75628 26290 75684 26302
rect 75628 26238 75630 26290
rect 75682 26238 75684 26290
rect 75292 26180 75348 26190
rect 75628 26180 75684 26238
rect 78204 26292 78260 26910
rect 78204 26226 78260 26236
rect 75348 26124 75684 26180
rect 75292 26086 75348 26124
rect 77980 26066 78036 26078
rect 77980 26014 77982 26066
rect 78034 26014 78036 26066
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 77980 25620 78036 26014
rect 77980 25554 78036 25564
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 77980 24948 78036 24958
rect 75740 24722 75796 24734
rect 75740 24670 75742 24722
rect 75794 24670 75796 24722
rect 75292 24612 75348 24622
rect 75292 24518 75348 24556
rect 75740 24612 75796 24670
rect 75740 24546 75796 24556
rect 77980 24610 78036 24892
rect 77980 24558 77982 24610
rect 78034 24558 78036 24610
rect 77980 24546 78036 24558
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 78204 24276 78260 24286
rect 78204 23826 78260 24220
rect 78204 23774 78206 23826
rect 78258 23774 78260 23826
rect 78204 23762 78260 23774
rect 77756 23714 77812 23726
rect 77756 23662 77758 23714
rect 77810 23662 77812 23714
rect 77756 23604 77812 23662
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 77756 23538 77812 23548
rect 50556 23482 50820 23492
rect 75740 23154 75796 23166
rect 75740 23102 75742 23154
rect 75794 23102 75796 23154
rect 75292 23044 75348 23054
rect 75292 22950 75348 22988
rect 75740 23044 75796 23102
rect 75740 22978 75796 22988
rect 77980 22932 78036 22942
rect 77980 22838 78036 22876
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 78204 22260 78260 22270
rect 78204 22166 78260 22204
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 75628 21588 75684 21598
rect 75292 21586 75684 21588
rect 75292 21534 75630 21586
rect 75682 21534 75684 21586
rect 75292 21532 75684 21534
rect 75292 21476 75348 21532
rect 75628 21522 75684 21532
rect 77980 21588 78036 21598
rect 75292 21382 75348 21420
rect 77980 21474 78036 21532
rect 77980 21422 77982 21474
rect 78034 21422 78036 21474
rect 77980 21410 78036 21422
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 77644 20916 77700 20926
rect 77644 20822 77700 20860
rect 78204 20916 78260 20926
rect 78204 20802 78260 20860
rect 78204 20750 78206 20802
rect 78258 20750 78260 20802
rect 78204 20738 78260 20750
rect 77868 20580 77924 20590
rect 77868 20486 77924 20524
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 77980 20132 78036 20142
rect 75628 20018 75684 20030
rect 75628 19966 75630 20018
rect 75682 19966 75684 20018
rect 46060 19842 46116 19852
rect 75292 19908 75348 19918
rect 75628 19908 75684 19966
rect 75348 19852 75684 19908
rect 77980 19906 78036 20076
rect 77980 19854 77982 19906
rect 78034 19854 78036 19906
rect 75292 19814 75348 19852
rect 77980 19842 78036 19854
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 44492 5842 44548 5852
rect 46396 5908 46452 5918
rect 43596 4162 43652 4172
rect 43708 5236 43764 5246
rect 43484 3490 43540 3500
rect 43708 3554 43764 5180
rect 45052 4452 45108 4462
rect 44268 4116 44324 4126
rect 44268 4022 44324 4060
rect 44604 3668 44660 3678
rect 44604 3574 44660 3612
rect 43708 3502 43710 3554
rect 43762 3502 43764 3554
rect 43708 3490 43764 3502
rect 43036 2044 43204 2100
rect 43820 3444 43876 3454
rect 43036 800 43092 2044
rect 43820 1316 43876 3388
rect 43708 1260 43876 1316
rect 44380 3444 44436 3454
rect 43708 800 43764 1260
rect 44380 800 44436 3388
rect 45052 800 45108 4396
rect 46172 4452 46228 4462
rect 46172 4358 46228 4396
rect 46396 4340 46452 5852
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 46620 4450 46676 4462
rect 46620 4398 46622 4450
rect 46674 4398 46676 4450
rect 46396 4284 46564 4340
rect 46508 3442 46564 4284
rect 46508 3390 46510 3442
rect 46562 3390 46564 3442
rect 46508 3378 46564 3390
rect 46396 3332 46452 3342
rect 45836 980 45892 990
rect 45724 978 45892 980
rect 45724 926 45838 978
rect 45890 926 45892 978
rect 45724 924 45892 926
rect 45724 800 45780 924
rect 45836 914 45892 924
rect 46396 800 46452 3276
rect 46620 978 46676 4398
rect 51996 4340 52052 4350
rect 51660 4338 52052 4340
rect 51660 4286 51998 4338
rect 52050 4286 52052 4338
rect 51660 4284 52052 4286
rect 47180 4226 47236 4238
rect 47180 4174 47182 4226
rect 47234 4174 47236 4226
rect 46732 3556 46788 3566
rect 47180 3556 47236 4174
rect 50876 4226 50932 4238
rect 50876 4174 50878 4226
rect 50930 4174 50932 4226
rect 46732 3554 47236 3556
rect 46732 3502 46734 3554
rect 46786 3502 47236 3554
rect 46732 3500 47236 3502
rect 50428 3668 50484 3678
rect 46732 3444 46788 3500
rect 46732 3378 46788 3388
rect 47404 3332 47460 3342
rect 47404 3238 47460 3276
rect 47852 3330 47908 3342
rect 48300 3332 48356 3342
rect 48748 3332 48804 3342
rect 49308 3332 49364 3342
rect 49980 3332 50036 3342
rect 47852 3278 47854 3330
rect 47906 3278 47908 3330
rect 46620 926 46622 978
rect 46674 926 46676 978
rect 46620 914 46676 926
rect 47068 1874 47124 1886
rect 47068 1822 47070 1874
rect 47122 1822 47124 1874
rect 47068 800 47124 1822
rect 47852 1874 47908 3278
rect 47852 1822 47854 1874
rect 47906 1822 47908 1874
rect 47852 1810 47908 1822
rect 47964 3330 48356 3332
rect 47964 3278 48302 3330
rect 48354 3278 48356 3330
rect 47964 3276 48356 3278
rect 47964 1652 48020 3276
rect 48300 3266 48356 3276
rect 48412 3330 48804 3332
rect 48412 3278 48750 3330
rect 48802 3278 48804 3330
rect 48412 3276 48804 3278
rect 47740 1596 48020 1652
rect 47740 800 47796 1596
rect 48412 800 48468 3276
rect 48748 3266 48804 3276
rect 49084 3330 49364 3332
rect 49084 3278 49310 3330
rect 49362 3278 49364 3330
rect 49084 3276 49364 3278
rect 49084 800 49140 3276
rect 49308 3266 49364 3276
rect 49756 3330 50036 3332
rect 49756 3278 49982 3330
rect 50034 3278 50036 3330
rect 49756 3276 50036 3278
rect 49756 800 49812 3276
rect 49980 3266 50036 3276
rect 50428 800 50484 3612
rect 50876 3556 50932 4174
rect 51660 4228 51716 4284
rect 51996 4274 52052 4284
rect 51660 4134 51716 4172
rect 51772 4116 51828 4126
rect 50876 3490 50932 3500
rect 51212 3556 51268 3566
rect 51212 3462 51268 3500
rect 50652 3332 50708 3342
rect 50652 3330 51156 3332
rect 50652 3278 50654 3330
rect 50706 3278 51156 3330
rect 50652 3276 51156 3278
rect 50652 3266 50708 3276
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 51100 800 51156 3276
rect 51772 800 51828 4060
rect 53004 4116 53060 4126
rect 53004 4022 53060 4060
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 52220 3668 52276 3678
rect 52220 3574 52276 3612
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32256 0 32368 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 34272 0 34384 800
rect 34944 0 35056 800
rect 35616 0 35728 800
rect 36288 0 36400 800
rect 36960 0 37072 800
rect 37632 0 37744 800
rect 38304 0 38416 800
rect 38976 0 39088 800
rect 39648 0 39760 800
rect 40320 0 40432 800
rect 40992 0 41104 800
rect 41664 0 41776 800
rect 42336 0 42448 800
rect 43008 0 43120 800
rect 43680 0 43792 800
rect 44352 0 44464 800
rect 45024 0 45136 800
rect 45696 0 45808 800
rect 46368 0 46480 800
rect 47040 0 47152 800
rect 47712 0 47824 800
rect 48384 0 48496 800
rect 49056 0 49168 800
rect 49728 0 49840 800
rect 50400 0 50512 800
rect 51072 0 51184 800
rect 51744 0 51856 800
rect 52416 0 52528 800
rect 53088 0 53200 800
rect 53760 0 53872 800
rect 54432 0 54544 800
rect 55104 0 55216 800
rect 55776 0 55888 800
rect 56448 0 56560 800
rect 57120 0 57232 800
rect 57792 0 57904 800
rect 58464 0 58576 800
rect 59136 0 59248 800
rect 59808 0 59920 800
rect 60480 0 60592 800
rect 61152 0 61264 800
rect 61824 0 61936 800
rect 62496 0 62608 800
rect 63168 0 63280 800
rect 63840 0 63952 800
rect 64512 0 64624 800
rect 65184 0 65296 800
rect 65856 0 65968 800
rect 66528 0 66640 800
rect 67200 0 67312 800
rect 67872 0 67984 800
rect 68544 0 68656 800
rect 69216 0 69328 800
rect 69888 0 70000 800
rect 70560 0 70672 800
rect 71232 0 71344 800
rect 71904 0 72016 800
rect 72576 0 72688 800
rect 73248 0 73360 800
rect 73920 0 74032 800
rect 74592 0 74704 800
rect 75264 0 75376 800
rect 75936 0 76048 800
rect 76608 0 76720 800
rect 77280 0 77392 800
rect 77952 0 78064 800
rect 78624 0 78736 800
rect 79296 0 79408 800
<< via2 >>
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 22876 76466 22932 76468
rect 22876 76414 22878 76466
rect 22878 76414 22930 76466
rect 22930 76414 22932 76466
rect 22876 76412 22932 76414
rect 23548 76412 23604 76468
rect 24556 76466 24612 76468
rect 24556 76414 24558 76466
rect 24558 76414 24610 76466
rect 24610 76414 24612 76466
rect 24556 76412 24612 76414
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 1932 67228 1988 67284
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 27580 76300 27636 76356
rect 1708 66556 1764 66612
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 1708 66050 1764 66052
rect 1708 65998 1710 66050
rect 1710 65998 1762 66050
rect 1762 65998 1764 66050
rect 1708 65996 1764 65998
rect 1708 65212 1764 65268
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 1708 64594 1764 64596
rect 1708 64542 1710 64594
rect 1710 64542 1762 64594
rect 1762 64542 1764 64594
rect 1708 64540 1764 64542
rect 1708 63196 1764 63252
rect 1708 62914 1764 62916
rect 1708 62862 1710 62914
rect 1710 62862 1762 62914
rect 1762 62862 1764 62914
rect 1708 62860 1764 62862
rect 1708 61852 1764 61908
rect 1708 61346 1764 61348
rect 1708 61294 1710 61346
rect 1710 61294 1762 61346
rect 1762 61294 1764 61346
rect 1708 61292 1764 61294
rect 1708 60508 1764 60564
rect 1820 59164 1876 59220
rect 1708 58492 1764 58548
rect 1708 58210 1764 58212
rect 1708 58158 1710 58210
rect 1710 58158 1762 58210
rect 1762 58158 1764 58210
rect 1708 58156 1764 58158
rect 1708 57148 1764 57204
rect 1708 56642 1764 56644
rect 1708 56590 1710 56642
rect 1710 56590 1762 56642
rect 1762 56590 1764 56642
rect 1708 56588 1764 56590
rect 1708 55804 1764 55860
rect 1708 54908 1764 54964
rect 1708 53788 1764 53844
rect 1820 53116 1876 53172
rect 1708 52444 1764 52500
rect 1708 51938 1764 51940
rect 1708 51886 1710 51938
rect 1710 51886 1762 51938
rect 1762 51886 1764 51938
rect 1708 51884 1764 51886
rect 1708 51100 1764 51156
rect 1820 49756 1876 49812
rect 2940 64594 2996 64596
rect 2940 64542 2942 64594
rect 2942 64542 2994 64594
rect 2994 64542 2996 64594
rect 2940 64540 2996 64542
rect 2380 63868 2436 63924
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 2492 60508 2548 60564
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 2156 59890 2212 59892
rect 2156 59838 2158 59890
rect 2158 59838 2210 59890
rect 2210 59838 2212 59890
rect 2156 59836 2212 59838
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 2156 55186 2212 55188
rect 2156 55134 2158 55186
rect 2158 55134 2210 55186
rect 2210 55134 2212 55186
rect 2156 55132 2212 55134
rect 2156 50428 2212 50484
rect 1708 49084 1764 49140
rect 1708 48524 1764 48580
rect 1708 47740 1764 47796
rect 1708 47234 1764 47236
rect 1708 47182 1710 47234
rect 1710 47182 1762 47234
rect 1762 47182 1764 47234
rect 1708 47180 1764 47182
rect 1708 46396 1764 46452
rect 1708 45052 1764 45108
rect 1932 44380 1988 44436
rect 1708 44098 1764 44100
rect 1708 44046 1710 44098
rect 1710 44046 1762 44098
rect 1762 44046 1764 44098
rect 1708 44044 1764 44046
rect 2156 45778 2212 45780
rect 2156 45726 2158 45778
rect 2158 45726 2210 45778
rect 2210 45726 2212 45778
rect 2156 45724 2212 45726
rect 2492 53116 2548 53172
rect 2380 44156 2436 44212
rect 1708 43036 1764 43092
rect 1708 42530 1764 42532
rect 1708 42478 1710 42530
rect 1710 42478 1762 42530
rect 1762 42478 1764 42530
rect 1708 42476 1764 42478
rect 1932 41746 1988 41748
rect 1932 41694 1934 41746
rect 1934 41694 1986 41746
rect 1986 41694 1988 41746
rect 1932 41692 1988 41694
rect 1708 41074 1764 41076
rect 1708 41022 1710 41074
rect 1710 41022 1762 41074
rect 1762 41022 1764 41074
rect 1708 41020 1764 41022
rect 2156 40348 2212 40404
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4284 45106 4340 45108
rect 4284 45054 4286 45106
rect 4286 45054 4338 45106
rect 4338 45054 4340 45106
rect 4284 45052 4340 45054
rect 4844 45106 4900 45108
rect 4844 45054 4846 45106
rect 4846 45054 4898 45106
rect 4898 45054 4900 45106
rect 4844 45052 4900 45054
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4284 41804 4340 41860
rect 4844 41858 4900 41860
rect 4844 41806 4846 41858
rect 4846 41806 4898 41858
rect 4898 41806 4900 41858
rect 4844 41804 4900 41806
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 2604 40908 2660 40964
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 25004 46844 25060 46900
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 25452 44268 25508 44324
rect 28588 76354 28644 76356
rect 28588 76302 28590 76354
rect 28590 76302 28642 76354
rect 28642 76302 28644 76354
rect 28588 76300 28644 76302
rect 34300 76354 34356 76356
rect 34300 76302 34302 76354
rect 34302 76302 34354 76354
rect 34354 76302 34356 76354
rect 34300 76300 34356 76302
rect 35980 76300 36036 76356
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 29484 47180 29540 47236
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 40348 75852 40404 75908
rect 41580 75906 41636 75908
rect 41580 75854 41582 75906
rect 41582 75854 41634 75906
rect 41634 75854 41636 75906
rect 41580 75852 41636 75854
rect 39788 74732 39844 74788
rect 38892 73948 38948 74004
rect 36316 48412 36372 48468
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35532 47234 35588 47236
rect 35532 47182 35534 47234
rect 35534 47182 35586 47234
rect 35586 47182 35588 47234
rect 35532 47180 35588 47182
rect 34748 46898 34804 46900
rect 34748 46846 34750 46898
rect 34750 46846 34802 46898
rect 34802 46846 34804 46898
rect 34748 46844 34804 46846
rect 31724 46620 31780 46676
rect 35420 46620 35476 46676
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 34860 45052 34916 45108
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 36428 44322 36484 44324
rect 36428 44270 36430 44322
rect 36430 44270 36482 44322
rect 36482 44270 36484 44322
rect 36428 44268 36484 44270
rect 34076 44210 34132 44212
rect 34076 44158 34078 44210
rect 34078 44158 34130 44210
rect 34130 44158 34132 44210
rect 34076 44156 34132 44158
rect 27804 44044 27860 44100
rect 35532 44098 35588 44100
rect 35532 44046 35534 44098
rect 35534 44046 35586 44098
rect 35586 44046 35588 44098
rect 35532 44044 35588 44046
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 39788 73948 39844 74004
rect 41020 74786 41076 74788
rect 41020 74734 41022 74786
rect 41022 74734 41074 74786
rect 41074 74734 41076 74786
rect 41020 74732 41076 74734
rect 39564 48466 39620 48468
rect 39564 48414 39566 48466
rect 39566 48414 39618 48466
rect 39618 48414 39620 48466
rect 39564 48412 39620 48414
rect 41244 74732 41300 74788
rect 42588 74732 42644 74788
rect 43260 74786 43316 74788
rect 43260 74734 43262 74786
rect 43262 74734 43314 74786
rect 43314 74734 43316 74786
rect 43260 74732 43316 74734
rect 44380 70476 44436 70532
rect 43372 48130 43428 48132
rect 43372 48078 43374 48130
rect 43374 48078 43426 48130
rect 43426 48078 43428 48130
rect 43372 48076 43428 48078
rect 42924 46956 42980 47012
rect 47740 76466 47796 76468
rect 47740 76414 47742 76466
rect 47742 76414 47794 76466
rect 47794 76414 47796 76466
rect 47740 76412 47796 76414
rect 48412 76412 48468 76468
rect 48860 76466 48916 76468
rect 48860 76414 48862 76466
rect 48862 76414 48914 76466
rect 48914 76414 48916 76466
rect 48860 76412 48916 76414
rect 49756 76636 49812 76692
rect 50092 76354 50148 76356
rect 50092 76302 50094 76354
rect 50094 76302 50146 76354
rect 50146 76302 50148 76354
rect 50092 76300 50148 76302
rect 48636 70476 48692 70532
rect 46508 46844 46564 46900
rect 50092 46956 50148 47012
rect 47180 46898 47236 46900
rect 47180 46846 47182 46898
rect 47182 46846 47234 46898
rect 47234 46846 47236 46898
rect 47180 46844 47236 46846
rect 46732 46786 46788 46788
rect 46732 46734 46734 46786
rect 46734 46734 46786 46786
rect 46786 46734 46788 46786
rect 46732 46732 46788 46734
rect 45164 46508 45220 46564
rect 41468 45106 41524 45108
rect 41468 45054 41470 45106
rect 41470 45054 41522 45106
rect 41522 45054 41524 45106
rect 41468 45052 41524 45054
rect 42028 45106 42084 45108
rect 42028 45054 42030 45106
rect 42030 45054 42082 45106
rect 42082 45054 42084 45106
rect 42028 45052 42084 45054
rect 45612 45330 45668 45332
rect 45612 45278 45614 45330
rect 45614 45278 45666 45330
rect 45666 45278 45668 45330
rect 45612 45276 45668 45278
rect 46172 45330 46228 45332
rect 46172 45278 46174 45330
rect 46174 45278 46226 45330
rect 46226 45278 46228 45330
rect 46172 45276 46228 45278
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 51212 76300 51268 76356
rect 52220 76690 52276 76692
rect 52220 76638 52222 76690
rect 52222 76638 52274 76690
rect 52274 76638 52276 76690
rect 52220 76636 52276 76638
rect 51772 75740 51828 75796
rect 51100 75068 51156 75124
rect 51660 75682 51716 75684
rect 51660 75630 51662 75682
rect 51662 75630 51714 75682
rect 51714 75630 51716 75682
rect 51660 75628 51716 75630
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50316 45276 50372 45332
rect 42700 44492 42756 44548
rect 44940 44434 44996 44436
rect 44940 44382 44942 44434
rect 44942 44382 44994 44434
rect 44994 44382 44996 44434
rect 44940 44380 44996 44382
rect 53116 77196 53172 77252
rect 53788 75794 53844 75796
rect 53788 75742 53790 75794
rect 53790 75742 53842 75794
rect 53842 75742 53844 75794
rect 53788 75740 53844 75742
rect 52668 75682 52724 75684
rect 52668 75630 52670 75682
rect 52670 75630 52722 75682
rect 52722 75630 52724 75682
rect 52668 75628 52724 75630
rect 52332 75122 52388 75124
rect 52332 75070 52334 75122
rect 52334 75070 52386 75122
rect 52386 75070 52388 75122
rect 52332 75068 52388 75070
rect 51548 44492 51604 44548
rect 51324 44380 51380 44436
rect 43148 44210 43204 44212
rect 43148 44158 43150 44210
rect 43150 44158 43202 44210
rect 43202 44158 43204 44210
rect 43148 44156 43204 44158
rect 43596 44210 43652 44212
rect 43596 44158 43598 44210
rect 43598 44158 43650 44210
rect 43650 44158 43652 44210
rect 43596 44156 43652 44158
rect 45388 44098 45444 44100
rect 45388 44046 45390 44098
rect 45390 44046 45442 44098
rect 45442 44046 45444 44098
rect 45388 44044 45444 44046
rect 45836 44098 45892 44100
rect 45836 44046 45838 44098
rect 45838 44046 45890 44098
rect 45890 44046 45892 44098
rect 45836 44044 45892 44046
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 45836 42754 45892 42756
rect 45836 42702 45838 42754
rect 45838 42702 45890 42754
rect 45890 42702 45892 42754
rect 45836 42700 45892 42702
rect 46396 42530 46452 42532
rect 46396 42478 46398 42530
rect 46398 42478 46450 42530
rect 46450 42478 46452 42530
rect 46396 42476 46452 42478
rect 46844 42530 46900 42532
rect 46844 42478 46846 42530
rect 46846 42478 46898 42530
rect 46898 42478 46900 42530
rect 46844 42476 46900 42478
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 45388 41970 45444 41972
rect 45388 41918 45390 41970
rect 45390 41918 45442 41970
rect 45442 41918 45444 41970
rect 45388 41916 45444 41918
rect 45948 41970 46004 41972
rect 45948 41918 45950 41970
rect 45950 41918 46002 41970
rect 46002 41918 46004 41970
rect 45948 41916 46004 41918
rect 55132 76636 55188 76692
rect 55692 77196 55748 77252
rect 56140 76690 56196 76692
rect 56140 76638 56142 76690
rect 56142 76638 56194 76690
rect 56194 76638 56196 76690
rect 56140 76636 56196 76638
rect 58492 76636 58548 76692
rect 59836 76690 59892 76692
rect 59836 76638 59838 76690
rect 59838 76638 59890 76690
rect 59890 76638 59892 76690
rect 59836 76636 59892 76638
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 77868 57820 77924 57876
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 77644 56476 77700 56532
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 58492 48076 58548 48132
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 56588 45052 56644 45108
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 55020 44156 55076 44212
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 75068 42700 75124 42756
rect 54124 41916 54180 41972
rect 34412 41804 34468 41860
rect 44940 41858 44996 41860
rect 44940 41806 44942 41858
rect 44942 41806 44994 41858
rect 44994 41806 44996 41858
rect 44940 41804 44996 41806
rect 75404 46562 75460 46564
rect 75404 46510 75406 46562
rect 75406 46510 75458 46562
rect 75458 46510 75460 46562
rect 75404 46508 75460 46510
rect 77756 55186 77812 55188
rect 77756 55134 77758 55186
rect 77758 55134 77810 55186
rect 77810 55134 77812 55186
rect 77756 55132 77812 55134
rect 77868 53788 77924 53844
rect 77644 51100 77700 51156
rect 77756 50370 77812 50372
rect 77756 50318 77758 50370
rect 77758 50318 77810 50370
rect 77810 50318 77812 50370
rect 77756 50316 77812 50318
rect 77532 44044 77588 44100
rect 77868 46956 77924 47012
rect 78204 58828 78260 58884
rect 78204 57148 78260 57204
rect 78204 56476 78260 56532
rect 78204 55804 78260 55860
rect 78204 54460 78260 54516
rect 78204 53116 78260 53172
rect 78204 52444 78260 52500
rect 78204 51772 78260 51828
rect 78204 51100 78260 51156
rect 78428 49756 78484 49812
rect 78204 49084 78260 49140
rect 78204 48802 78260 48804
rect 78204 48750 78206 48802
rect 78206 48750 78258 48802
rect 78258 48750 78260 48802
rect 78204 48748 78260 48750
rect 78204 47740 78260 47796
rect 77980 46732 78036 46788
rect 78204 46396 78260 46452
rect 77756 45778 77812 45780
rect 77756 45726 77758 45778
rect 77758 45726 77810 45778
rect 77810 45726 77812 45778
rect 77756 45724 77812 45726
rect 78204 45388 78260 45444
rect 78204 44380 78260 44436
rect 78428 43708 78484 43764
rect 78204 43036 78260 43092
rect 77644 42476 77700 42532
rect 78204 42364 78260 42420
rect 75292 41804 75348 41860
rect 78204 41692 78260 41748
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 78204 41074 78260 41076
rect 78204 41022 78206 41074
rect 78206 41022 78258 41074
rect 78258 41022 78260 41074
rect 78204 41020 78260 41022
rect 33628 40962 33684 40964
rect 33628 40910 33630 40962
rect 33630 40910 33682 40962
rect 33682 40910 33684 40962
rect 33628 40908 33684 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 4956 40460 5012 40516
rect 35084 40460 35140 40516
rect 2380 40348 2436 40404
rect 34412 40402 34468 40404
rect 34412 40350 34414 40402
rect 34414 40350 34466 40402
rect 34466 40350 34468 40402
rect 34412 40348 34468 40350
rect 77756 40348 77812 40404
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 78204 39900 78260 39956
rect 1708 39676 1764 39732
rect 40012 39394 40068 39396
rect 40012 39342 40014 39394
rect 40014 39342 40066 39394
rect 40066 39342 40068 39394
rect 40012 39340 40068 39342
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 1708 39004 1764 39060
rect 2044 38946 2100 38948
rect 2044 38894 2046 38946
rect 2046 38894 2098 38946
rect 2098 38894 2100 38946
rect 2044 38892 2100 38894
rect 40012 38892 40068 38948
rect 1708 38332 1764 38388
rect 2492 38332 2548 38388
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 1708 37826 1764 37828
rect 1708 37774 1710 37826
rect 1710 37774 1762 37826
rect 1762 37774 1764 37826
rect 1708 37772 1764 37774
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 2044 37378 2100 37380
rect 2044 37326 2046 37378
rect 2046 37326 2098 37378
rect 2098 37326 2100 37378
rect 2044 37324 2100 37326
rect 1708 36988 1764 37044
rect 2044 37100 2100 37156
rect 1708 36370 1764 36372
rect 1708 36318 1710 36370
rect 1710 36318 1762 36370
rect 1762 36318 1764 36370
rect 1708 36316 1764 36318
rect 2492 36988 2548 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 2940 36370 2996 36372
rect 2940 36318 2942 36370
rect 2942 36318 2994 36370
rect 2994 36318 2996 36370
rect 2940 36316 2996 36318
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 2380 35644 2436 35700
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 1708 34972 1764 35028
rect 2044 34690 2100 34692
rect 2044 34638 2046 34690
rect 2046 34638 2098 34690
rect 2098 34638 2100 34690
rect 2044 34636 2100 34638
rect 1820 34300 1876 34356
rect 32620 34636 32676 34692
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 2492 34300 2548 34356
rect 1708 33628 1764 33684
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 1708 32956 1764 33012
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 2044 32674 2100 32676
rect 2044 32622 2046 32674
rect 2046 32622 2098 32674
rect 2098 32622 2100 32674
rect 2044 32620 2100 32622
rect 1708 32284 1764 32340
rect 2492 32284 2548 32340
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 1708 31612 1764 31668
rect 1708 31164 1764 31220
rect 4284 31778 4340 31780
rect 4284 31726 4286 31778
rect 4286 31726 4338 31778
rect 4338 31726 4340 31778
rect 4284 31724 4340 31726
rect 4844 31778 4900 31780
rect 4844 31726 4846 31778
rect 4846 31726 4898 31778
rect 4898 31726 4900 31778
rect 4844 31724 4900 31726
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 2940 31218 2996 31220
rect 2940 31166 2942 31218
rect 2942 31166 2994 31218
rect 2994 31166 2996 31218
rect 2940 31164 2996 31166
rect 2044 31106 2100 31108
rect 2044 31054 2046 31106
rect 2046 31054 2098 31106
rect 2098 31054 2100 31106
rect 2044 31052 2100 31054
rect 1932 30940 1988 30996
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 2380 30268 2436 30324
rect 4284 29932 4340 29988
rect 4844 29986 4900 29988
rect 4844 29934 4846 29986
rect 4846 29934 4898 29986
rect 4898 29934 4900 29986
rect 4844 29932 4900 29934
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 2492 29596 2548 29652
rect 1708 29202 1764 29204
rect 1708 29150 1710 29202
rect 1710 29150 1762 29202
rect 1762 29150 1764 29202
rect 1708 29148 1764 29150
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4284 28642 4340 28644
rect 4284 28590 4286 28642
rect 4286 28590 4338 28642
rect 4338 28590 4340 28642
rect 4284 28588 4340 28590
rect 4844 28642 4900 28644
rect 4844 28590 4846 28642
rect 4846 28590 4898 28642
rect 4898 28590 4900 28642
rect 4844 28588 4900 28590
rect 1932 28252 1988 28308
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 1708 27580 1764 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 1708 26908 1764 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 2156 26236 2212 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 1708 25564 1764 25620
rect 1708 25004 1764 25060
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 1708 24220 1764 24276
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 1708 23714 1764 23716
rect 1708 23662 1710 23714
rect 1710 23662 1762 23714
rect 1762 23662 1764 23714
rect 1708 23660 1764 23662
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 1708 22876 1764 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 1708 22204 1764 22260
rect 4284 22370 4340 22372
rect 4284 22318 4286 22370
rect 4286 22318 4338 22370
rect 4338 22318 4340 22370
rect 4284 22316 4340 22318
rect 4844 22370 4900 22372
rect 4844 22318 4846 22370
rect 4846 22318 4898 22370
rect 4898 22318 4900 22370
rect 4844 22316 4900 22318
rect 2940 22204 2996 22260
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 2044 21698 2100 21700
rect 2044 21646 2046 21698
rect 2046 21646 2098 21698
rect 2098 21646 2100 21698
rect 2044 21644 2100 21646
rect 1932 21532 1988 21588
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 2380 20860 2436 20916
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 1708 20188 1764 20244
rect 2044 20130 2100 20132
rect 2044 20078 2046 20130
rect 2046 20078 2098 20130
rect 2098 20078 2100 20130
rect 2044 20076 2100 20078
rect 1708 19516 1764 19572
rect 2492 19516 2548 19572
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 1708 19010 1764 19012
rect 1708 18958 1710 19010
rect 1710 18958 1762 19010
rect 1762 18958 1764 19010
rect 1708 18956 1764 18958
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 1708 18172 1764 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1708 17500 1764 17556
rect 1708 17106 1764 17108
rect 1708 17054 1710 17106
rect 1710 17054 1762 17106
rect 1762 17054 1764 17106
rect 1708 17052 1764 17054
rect 4284 17388 4340 17444
rect 4844 17442 4900 17444
rect 4844 17390 4846 17442
rect 4846 17390 4898 17442
rect 4898 17390 4900 17442
rect 4844 17388 4900 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 2940 17106 2996 17108
rect 2940 17054 2942 17106
rect 2942 17054 2994 17106
rect 2994 17054 2996 17106
rect 2940 17052 2996 17054
rect 1932 16828 1988 16884
rect 2044 16716 2100 16772
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 2380 16156 2436 16212
rect 1708 15874 1764 15876
rect 1708 15822 1710 15874
rect 1710 15822 1762 15874
rect 1762 15822 1764 15874
rect 1708 15820 1764 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 1708 14812 1764 14868
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 1708 14306 1764 14308
rect 1708 14254 1710 14306
rect 1710 14254 1762 14306
rect 1762 14254 1764 14306
rect 1708 14252 1764 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 1708 13522 1764 13524
rect 1708 13470 1710 13522
rect 1710 13470 1762 13522
rect 1762 13470 1764 13522
rect 1708 13468 1764 13470
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 1708 12796 1764 12852
rect 4284 12684 4340 12740
rect 4844 12738 4900 12740
rect 4844 12686 4846 12738
rect 4846 12686 4898 12738
rect 4898 12686 4900 12738
rect 4844 12684 4900 12686
rect 33516 37154 33572 37156
rect 33516 37102 33518 37154
rect 33518 37102 33570 37154
rect 33570 37102 33572 37154
rect 33516 37100 33572 37102
rect 33964 31052 34020 31108
rect 34188 34130 34244 34132
rect 34188 34078 34190 34130
rect 34190 34078 34242 34130
rect 34242 34078 34244 34130
rect 34188 34076 34244 34078
rect 34076 22316 34132 22372
rect 34636 34130 34692 34132
rect 34636 34078 34638 34130
rect 34638 34078 34690 34130
rect 34690 34078 34692 34130
rect 34636 34076 34692 34078
rect 33628 21644 33684 21700
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 34860 32620 34916 32676
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34972 31724 35028 31780
rect 34524 20076 34580 20132
rect 34412 17388 34468 17444
rect 33404 12684 33460 12740
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 1932 12124 1988 12180
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35868 29932 35924 29988
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35084 6748 35140 6804
rect 35980 6748 36036 6804
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 29596 4172 29652 4228
rect 30156 4226 30212 4228
rect 30156 4174 30158 4226
rect 30158 4174 30210 4226
rect 30210 4174 30212 4226
rect 30156 4172 30212 4174
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 26796 3442 26852 3444
rect 26796 3390 26798 3442
rect 26798 3390 26850 3442
rect 26850 3390 26852 3442
rect 26796 3388 26852 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 27244 3554 27300 3556
rect 27244 3502 27246 3554
rect 27246 3502 27298 3554
rect 27298 3502 27300 3554
rect 27244 3500 27300 3502
rect 28252 3500 28308 3556
rect 27580 3388 27636 3444
rect 27804 3442 27860 3444
rect 27804 3390 27806 3442
rect 27806 3390 27858 3442
rect 27858 3390 27860 3442
rect 27804 3388 27860 3390
rect 28812 3500 28868 3556
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 38780 28588 38836 28644
rect 38332 3500 38388 3556
rect 39564 5180 39620 5236
rect 40124 35532 40180 35588
rect 41132 39394 41188 39396
rect 41132 39342 41134 39394
rect 41134 39342 41186 39394
rect 41186 39342 41188 39394
rect 41132 39340 41188 39342
rect 40348 21420 40404 21476
rect 41020 35586 41076 35588
rect 41020 35534 41022 35586
rect 41022 35534 41074 35586
rect 41074 35534 41076 35586
rect 41020 35532 41076 35534
rect 40908 20524 40964 20580
rect 40460 5628 40516 5684
rect 39788 4172 39844 4228
rect 38892 3388 38948 3444
rect 43708 37324 43764 37380
rect 43148 35698 43204 35700
rect 43148 35646 43150 35698
rect 43150 35646 43202 35698
rect 43202 35646 43204 35698
rect 43148 35644 43204 35646
rect 41692 22988 41748 23044
rect 41916 35532 41972 35588
rect 41692 3500 41748 3556
rect 44156 35698 44212 35700
rect 44156 35646 44158 35698
rect 44158 35646 44210 35698
rect 44210 35646 44212 35698
rect 44156 35644 44212 35646
rect 42476 5628 42532 5684
rect 42476 5068 42532 5124
rect 42364 3612 42420 3668
rect 42140 3554 42196 3556
rect 42140 3502 42142 3554
rect 42142 3502 42194 3554
rect 42194 3502 42196 3554
rect 42140 3500 42196 3502
rect 42812 3388 42868 3444
rect 43148 5180 43204 5236
rect 43260 5068 43316 5124
rect 43148 4060 43204 4116
rect 44044 32562 44100 32564
rect 44044 32510 44046 32562
rect 44046 32510 44098 32562
rect 44098 32510 44100 32562
rect 44044 32508 44100 32510
rect 44380 16716 44436 16772
rect 44492 32562 44548 32564
rect 44492 32510 44494 32562
rect 44494 32510 44546 32562
rect 44546 32510 44548 32562
rect 44492 32508 44548 32510
rect 44940 26124 44996 26180
rect 45276 30828 45332 30884
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 78204 39004 78260 39060
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 78204 38332 78260 38388
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 78204 37660 78260 37716
rect 50764 37604 50820 37606
rect 78204 36988 78260 37044
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 78204 36370 78260 36372
rect 78204 36318 78206 36370
rect 78206 36318 78258 36370
rect 78258 36318 78260 36370
rect 78204 36316 78260 36318
rect 77756 35644 77812 35700
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 78204 34972 78260 35028
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 78204 34300 78260 34356
rect 77868 34242 77924 34244
rect 77868 34190 77870 34242
rect 77870 34190 77922 34242
rect 77922 34190 77924 34242
rect 77868 34188 77924 34190
rect 45388 27020 45444 27076
rect 45052 24556 45108 24612
rect 46620 33964 46676 34020
rect 47068 34018 47124 34020
rect 47068 33966 47070 34018
rect 47070 33966 47122 34018
rect 47122 33966 47124 34018
rect 47068 33964 47124 33966
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 78204 33628 78260 33684
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 78204 32956 78260 33012
rect 50764 32900 50820 32902
rect 78204 32284 78260 32340
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 78204 31666 78260 31668
rect 78204 31614 78206 31666
rect 78206 31614 78258 31666
rect 78258 31614 78260 31666
rect 78204 31612 78260 31614
rect 77756 30940 77812 30996
rect 75292 30882 75348 30884
rect 75292 30830 75294 30882
rect 75294 30830 75346 30882
rect 75346 30830 75348 30882
rect 75292 30828 75348 30830
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 77980 30268 78036 30324
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 78428 29596 78484 29652
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 78204 28924 78260 28980
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 78204 28252 78260 28308
rect 50764 28196 50820 28198
rect 78204 27580 78260 27636
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 77196 27186 77252 27188
rect 77196 27134 77198 27186
rect 77198 27134 77250 27186
rect 77250 27134 77252 27186
rect 77196 27132 77252 27134
rect 78204 27132 78260 27188
rect 77868 27020 77924 27076
rect 77532 26850 77588 26852
rect 77532 26798 77534 26850
rect 77534 26798 77586 26850
rect 77586 26798 77588 26850
rect 77532 26796 77588 26798
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 78204 26236 78260 26292
rect 75292 26178 75348 26180
rect 75292 26126 75294 26178
rect 75294 26126 75346 26178
rect 75346 26126 75348 26178
rect 75292 26124 75348 26126
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 77980 25564 78036 25620
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 77980 24892 78036 24948
rect 75292 24610 75348 24612
rect 75292 24558 75294 24610
rect 75294 24558 75346 24610
rect 75346 24558 75348 24610
rect 75292 24556 75348 24558
rect 75740 24556 75796 24612
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 78204 24220 78260 24276
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 77756 23548 77812 23604
rect 50764 23492 50820 23494
rect 75292 23042 75348 23044
rect 75292 22990 75294 23042
rect 75294 22990 75346 23042
rect 75346 22990 75348 23042
rect 75292 22988 75348 22990
rect 75740 22988 75796 23044
rect 77980 22930 78036 22932
rect 77980 22878 77982 22930
rect 77982 22878 78034 22930
rect 78034 22878 78036 22930
rect 77980 22876 78036 22878
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 78204 22258 78260 22260
rect 78204 22206 78206 22258
rect 78206 22206 78258 22258
rect 78258 22206 78260 22258
rect 78204 22204 78260 22206
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 77980 21532 78036 21588
rect 75292 21474 75348 21476
rect 75292 21422 75294 21474
rect 75294 21422 75346 21474
rect 75346 21422 75348 21474
rect 75292 21420 75348 21422
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 77644 20914 77700 20916
rect 77644 20862 77646 20914
rect 77646 20862 77698 20914
rect 77698 20862 77700 20914
rect 77644 20860 77700 20862
rect 78204 20860 78260 20916
rect 77868 20578 77924 20580
rect 77868 20526 77870 20578
rect 77870 20526 77922 20578
rect 77922 20526 77924 20578
rect 77868 20524 77924 20526
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 77980 20076 78036 20132
rect 46060 19852 46116 19908
rect 75292 19906 75348 19908
rect 75292 19854 75294 19906
rect 75294 19854 75346 19906
rect 75346 19854 75348 19906
rect 75292 19852 75348 19854
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 44492 5852 44548 5908
rect 46396 5852 46452 5908
rect 43596 4172 43652 4228
rect 43708 5180 43764 5236
rect 43484 3500 43540 3556
rect 45052 4396 45108 4452
rect 44268 4114 44324 4116
rect 44268 4062 44270 4114
rect 44270 4062 44322 4114
rect 44322 4062 44324 4114
rect 44268 4060 44324 4062
rect 44604 3666 44660 3668
rect 44604 3614 44606 3666
rect 44606 3614 44658 3666
rect 44658 3614 44660 3666
rect 44604 3612 44660 3614
rect 43820 3388 43876 3444
rect 44380 3388 44436 3444
rect 46172 4450 46228 4452
rect 46172 4398 46174 4450
rect 46174 4398 46226 4450
rect 46226 4398 46228 4450
rect 46172 4396 46228 4398
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 46396 3276 46452 3332
rect 50428 3612 50484 3668
rect 46732 3388 46788 3444
rect 47404 3330 47460 3332
rect 47404 3278 47406 3330
rect 47406 3278 47458 3330
rect 47458 3278 47460 3330
rect 47404 3276 47460 3278
rect 51660 4226 51716 4228
rect 51660 4174 51662 4226
rect 51662 4174 51714 4226
rect 51714 4174 51716 4226
rect 51660 4172 51716 4174
rect 51772 4060 51828 4116
rect 50876 3500 50932 3556
rect 51212 3554 51268 3556
rect 51212 3502 51214 3554
rect 51214 3502 51266 3554
rect 51266 3502 51268 3554
rect 51212 3500 51268 3502
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 53004 4114 53060 4116
rect 53004 4062 53006 4114
rect 53006 4062 53058 4114
rect 53058 4062 53060 4114
rect 53004 4060 53060 4062
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 52220 3666 52276 3668
rect 52220 3614 52222 3666
rect 52222 3614 52274 3666
rect 52274 3614 52276 3666
rect 52220 3612 52276 3614
<< metal3 >>
rect 0 79296 800 79408
rect 79200 79296 80000 79408
rect 0 78624 800 78736
rect 79200 78624 80000 78736
rect 0 77952 800 78064
rect 79200 77952 80000 78064
rect 0 77280 800 77392
rect 79200 77280 80000 77392
rect 53106 77196 53116 77252
rect 53172 77196 55692 77252
rect 55748 77196 55758 77252
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 0 76608 800 76720
rect 49746 76636 49756 76692
rect 49812 76636 52220 76692
rect 52276 76636 52286 76692
rect 55122 76636 55132 76692
rect 55188 76636 56140 76692
rect 56196 76636 56206 76692
rect 58482 76636 58492 76692
rect 58548 76636 59836 76692
rect 59892 76636 59902 76692
rect 79200 76608 80000 76720
rect 22866 76412 22876 76468
rect 22932 76412 23548 76468
rect 23604 76412 24556 76468
rect 24612 76412 24622 76468
rect 47730 76412 47740 76468
rect 47796 76412 48412 76468
rect 48468 76412 48860 76468
rect 48916 76412 48926 76468
rect 27570 76300 27580 76356
rect 27636 76300 28588 76356
rect 28644 76300 28654 76356
rect 34290 76300 34300 76356
rect 34356 76300 35980 76356
rect 36036 76300 36046 76356
rect 50082 76300 50092 76356
rect 50148 76300 51212 76356
rect 51268 76300 51278 76356
rect 0 75936 800 76048
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 79200 75936 80000 76048
rect 40338 75852 40348 75908
rect 40404 75852 41580 75908
rect 41636 75852 41646 75908
rect 51762 75740 51772 75796
rect 51828 75740 53788 75796
rect 53844 75740 53854 75796
rect 51650 75628 51660 75684
rect 51716 75628 52668 75684
rect 52724 75628 52734 75684
rect 0 75264 800 75376
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 79200 75264 80000 75376
rect 51090 75068 51100 75124
rect 51156 75068 52332 75124
rect 52388 75068 52398 75124
rect 39778 74732 39788 74788
rect 39844 74732 41020 74788
rect 41076 74732 41086 74788
rect 41234 74732 41244 74788
rect 41300 74732 42588 74788
rect 42644 74732 43260 74788
rect 43316 74732 43326 74788
rect 0 74592 800 74704
rect 79200 74592 80000 74704
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 0 73920 800 74032
rect 38882 73948 38892 74004
rect 38948 73948 39788 74004
rect 39844 73948 39854 74004
rect 79200 73920 80000 74032
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 0 73248 800 73360
rect 79200 73248 80000 73360
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 0 72576 800 72688
rect 79200 72576 80000 72688
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 79200 71904 80000 72016
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 79200 71232 80000 71344
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 79200 70560 80000 70672
rect 44370 70476 44380 70532
rect 44436 70476 48636 70532
rect 48692 70476 48702 70532
rect 79200 69888 80000 70000
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 79200 69216 80000 69328
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 79200 68544 80000 68656
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 79200 67872 80000 67984
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 0 67284 800 67312
rect 0 67228 1932 67284
rect 1988 67228 1998 67284
rect 0 67200 800 67228
rect 79200 67200 80000 67312
rect 0 66612 800 66640
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 0 66556 1708 66612
rect 1764 66556 1774 66612
rect 0 66528 800 66556
rect 79200 66528 80000 66640
rect 1698 65996 1708 66052
rect 1764 65996 1774 66052
rect 0 65940 800 65968
rect 1708 65940 1764 65996
rect 0 65884 1764 65940
rect 0 65856 800 65884
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 79200 65856 80000 65968
rect 0 65268 800 65296
rect 0 65212 1708 65268
rect 1764 65212 1774 65268
rect 0 65184 800 65212
rect 79200 65184 80000 65296
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 0 64596 800 64624
rect 0 64540 1708 64596
rect 1764 64540 2940 64596
rect 2996 64540 3006 64596
rect 0 64512 800 64540
rect 79200 64512 80000 64624
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 0 63924 800 63952
rect 0 63868 2380 63924
rect 2436 63868 2446 63924
rect 0 63840 800 63868
rect 79200 63840 80000 63952
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 0 63252 800 63280
rect 0 63196 1708 63252
rect 1764 63196 1774 63252
rect 0 63168 800 63196
rect 79200 63168 80000 63280
rect 1698 62860 1708 62916
rect 1764 62860 1774 62916
rect 0 62580 800 62608
rect 1708 62580 1764 62860
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 0 62524 1764 62580
rect 0 62496 800 62524
rect 79200 62496 80000 62608
rect 0 61908 800 61936
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 0 61852 1708 61908
rect 1764 61852 1774 61908
rect 0 61824 800 61852
rect 79200 61824 80000 61936
rect 1698 61292 1708 61348
rect 1764 61292 1774 61348
rect 0 61236 800 61264
rect 1708 61236 1764 61292
rect 0 61180 1764 61236
rect 0 61152 800 61180
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 79200 61152 80000 61264
rect 0 60564 800 60592
rect 0 60508 1708 60564
rect 1764 60508 2492 60564
rect 2548 60508 2558 60564
rect 0 60480 800 60508
rect 79200 60480 80000 60592
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 0 59892 800 59920
rect 0 59836 2156 59892
rect 2212 59836 2222 59892
rect 0 59808 800 59836
rect 79200 59808 80000 59920
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 0 59220 800 59248
rect 0 59164 1820 59220
rect 1876 59164 1886 59220
rect 0 59136 800 59164
rect 79200 59136 80000 59248
rect 78194 58828 78204 58884
rect 78260 58828 78270 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 0 58548 800 58576
rect 78204 58548 78260 58828
rect 79200 58548 80000 58576
rect 0 58492 1708 58548
rect 1764 58492 1774 58548
rect 78204 58492 80000 58548
rect 0 58464 800 58492
rect 79200 58464 80000 58492
rect 1698 58156 1708 58212
rect 1764 58156 1774 58212
rect 1708 57988 1764 58156
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 924 57932 1764 57988
rect 0 57876 800 57904
rect 924 57876 980 57932
rect 79200 57876 80000 57904
rect 0 57820 980 57876
rect 77858 57820 77868 57876
rect 77924 57820 80000 57876
rect 0 57792 800 57820
rect 79200 57792 80000 57820
rect 0 57204 800 57232
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 79200 57204 80000 57232
rect 0 57148 1708 57204
rect 1764 57148 1774 57204
rect 78194 57148 78204 57204
rect 78260 57148 80000 57204
rect 0 57120 800 57148
rect 79200 57120 80000 57148
rect 1698 56588 1708 56644
rect 1764 56588 1774 56644
rect 0 56532 800 56560
rect 1708 56532 1764 56588
rect 79200 56532 80000 56560
rect 0 56476 1764 56532
rect 77634 56476 77644 56532
rect 77700 56476 78204 56532
rect 78260 56476 80000 56532
rect 0 56448 800 56476
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 79200 56448 80000 56476
rect 0 55860 800 55888
rect 79200 55860 80000 55888
rect 0 55804 1708 55860
rect 1764 55804 1774 55860
rect 78194 55804 78204 55860
rect 78260 55804 80000 55860
rect 0 55776 800 55804
rect 79200 55776 80000 55804
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 0 55188 800 55216
rect 79200 55188 80000 55216
rect 0 55132 2156 55188
rect 2212 55132 2222 55188
rect 77746 55132 77756 55188
rect 77812 55132 80000 55188
rect 0 55104 800 55132
rect 79200 55104 80000 55132
rect 1698 54908 1708 54964
rect 1764 54908 1774 54964
rect 1708 54852 1764 54908
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 924 54796 1764 54852
rect 0 54516 800 54544
rect 924 54516 980 54796
rect 79200 54516 80000 54544
rect 0 54460 980 54516
rect 78194 54460 78204 54516
rect 78260 54460 80000 54516
rect 0 54432 800 54460
rect 79200 54432 80000 54460
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 0 53844 800 53872
rect 79200 53844 80000 53872
rect 0 53788 1708 53844
rect 1764 53788 1774 53844
rect 77858 53788 77868 53844
rect 77924 53788 80000 53844
rect 0 53760 800 53788
rect 79200 53760 80000 53788
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 0 53172 800 53200
rect 79200 53172 80000 53200
rect 0 53116 1820 53172
rect 1876 53116 2492 53172
rect 2548 53116 2558 53172
rect 78194 53116 78204 53172
rect 78260 53116 80000 53172
rect 0 53088 800 53116
rect 79200 53088 80000 53116
rect 0 52500 800 52528
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 79200 52500 80000 52528
rect 0 52444 1708 52500
rect 1764 52444 1774 52500
rect 78194 52444 78204 52500
rect 78260 52444 80000 52500
rect 0 52416 800 52444
rect 79200 52416 80000 52444
rect 1698 51884 1708 51940
rect 1764 51884 1774 51940
rect 0 51828 800 51856
rect 1708 51828 1764 51884
rect 79200 51828 80000 51856
rect 0 51772 1764 51828
rect 78194 51772 78204 51828
rect 78260 51772 80000 51828
rect 0 51744 800 51772
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 79200 51744 80000 51772
rect 0 51156 800 51184
rect 79200 51156 80000 51184
rect 0 51100 1708 51156
rect 1764 51100 1774 51156
rect 77634 51100 77644 51156
rect 77700 51100 78204 51156
rect 78260 51100 80000 51156
rect 0 51072 800 51100
rect 79200 51072 80000 51100
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 0 50484 800 50512
rect 79200 50484 80000 50512
rect 0 50428 2156 50484
rect 2212 50428 2222 50484
rect 77756 50428 80000 50484
rect 0 50400 800 50428
rect 77756 50372 77812 50428
rect 79200 50400 80000 50428
rect 77746 50316 77756 50372
rect 77812 50316 77822 50372
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 0 49812 800 49840
rect 79200 49812 80000 49840
rect 0 49756 1820 49812
rect 1876 49756 1886 49812
rect 78418 49756 78428 49812
rect 78484 49756 80000 49812
rect 0 49728 800 49756
rect 79200 49728 80000 49756
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 0 49140 800 49168
rect 79200 49140 80000 49168
rect 0 49084 1708 49140
rect 1764 49084 1774 49140
rect 78194 49084 78204 49140
rect 78260 49084 80000 49140
rect 0 49056 800 49084
rect 79200 49056 80000 49084
rect 78194 48748 78204 48804
rect 78260 48748 78270 48804
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 1698 48524 1708 48580
rect 1764 48524 1774 48580
rect 0 48468 800 48496
rect 1708 48468 1764 48524
rect 78204 48468 78260 48748
rect 79200 48468 80000 48496
rect 0 48412 1764 48468
rect 36306 48412 36316 48468
rect 36372 48412 39564 48468
rect 39620 48412 39630 48468
rect 78204 48412 80000 48468
rect 0 48384 800 48412
rect 79200 48384 80000 48412
rect 43362 48076 43372 48132
rect 43428 48076 58492 48132
rect 58548 48076 58558 48132
rect 0 47796 800 47824
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 79200 47796 80000 47824
rect 0 47740 1708 47796
rect 1764 47740 1774 47796
rect 78194 47740 78204 47796
rect 78260 47740 80000 47796
rect 0 47712 800 47740
rect 79200 47712 80000 47740
rect 1698 47180 1708 47236
rect 1764 47180 1774 47236
rect 29474 47180 29484 47236
rect 29540 47180 35532 47236
rect 35588 47180 35598 47236
rect 0 47124 800 47152
rect 1708 47124 1764 47180
rect 79200 47124 80000 47152
rect 0 47068 1764 47124
rect 77868 47068 80000 47124
rect 0 47040 800 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 77868 47012 77924 47068
rect 79200 47040 80000 47068
rect 42914 46956 42924 47012
rect 42980 46956 50092 47012
rect 50148 46956 50158 47012
rect 77858 46956 77868 47012
rect 77924 46956 77934 47012
rect 24994 46844 25004 46900
rect 25060 46844 34748 46900
rect 34804 46844 34814 46900
rect 46498 46844 46508 46900
rect 46564 46844 47180 46900
rect 47236 46844 47246 46900
rect 46722 46732 46732 46788
rect 46788 46732 77980 46788
rect 78036 46732 78046 46788
rect 31714 46620 31724 46676
rect 31780 46620 35420 46676
rect 35476 46620 35486 46676
rect 45154 46508 45164 46564
rect 45220 46508 75404 46564
rect 75460 46508 75470 46564
rect 0 46452 800 46480
rect 79200 46452 80000 46480
rect 0 46396 1708 46452
rect 1764 46396 1774 46452
rect 78194 46396 78204 46452
rect 78260 46396 80000 46452
rect 0 46368 800 46396
rect 79200 46368 80000 46396
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 0 45780 800 45808
rect 79200 45780 80000 45808
rect 0 45724 2156 45780
rect 2212 45724 2222 45780
rect 77746 45724 77756 45780
rect 77812 45724 80000 45780
rect 0 45696 800 45724
rect 79200 45696 80000 45724
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 78194 45388 78204 45444
rect 78260 45388 78270 45444
rect 45602 45276 45612 45332
rect 45668 45276 46172 45332
rect 46228 45276 50316 45332
rect 50372 45276 50382 45332
rect 0 45108 800 45136
rect 78204 45108 78260 45388
rect 79200 45108 80000 45136
rect 0 45052 1708 45108
rect 1764 45052 1774 45108
rect 4274 45052 4284 45108
rect 4340 45052 4844 45108
rect 4900 45052 34860 45108
rect 34916 45052 34926 45108
rect 41458 45052 41468 45108
rect 41524 45052 42028 45108
rect 42084 45052 56588 45108
rect 56644 45052 56654 45108
rect 78204 45052 80000 45108
rect 0 45024 800 45052
rect 79200 45024 80000 45052
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 42690 44492 42700 44548
rect 42756 44492 51548 44548
rect 51604 44492 51614 44548
rect 0 44436 800 44464
rect 79200 44436 80000 44464
rect 0 44380 1932 44436
rect 1988 44380 1998 44436
rect 44930 44380 44940 44436
rect 44996 44380 51324 44436
rect 51380 44380 51390 44436
rect 78194 44380 78204 44436
rect 78260 44380 80000 44436
rect 0 44352 800 44380
rect 79200 44352 80000 44380
rect 25442 44268 25452 44324
rect 25508 44268 36428 44324
rect 36484 44268 36494 44324
rect 2370 44156 2380 44212
rect 2436 44156 34076 44212
rect 34132 44156 34142 44212
rect 43138 44156 43148 44212
rect 43204 44156 43596 44212
rect 43652 44156 55020 44212
rect 55076 44156 55086 44212
rect 1698 44044 1708 44100
rect 1764 44044 1774 44100
rect 27794 44044 27804 44100
rect 27860 44044 35532 44100
rect 35588 44044 35598 44100
rect 45378 44044 45388 44100
rect 45444 44044 45836 44100
rect 45892 44044 77532 44100
rect 77588 44044 77598 44100
rect 1708 43876 1764 44044
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 924 43820 1764 43876
rect 0 43764 800 43792
rect 924 43764 980 43820
rect 79200 43764 80000 43792
rect 0 43708 980 43764
rect 78418 43708 78428 43764
rect 78484 43708 80000 43764
rect 0 43680 800 43708
rect 79200 43680 80000 43708
rect 0 43092 800 43120
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 79200 43092 80000 43120
rect 0 43036 1708 43092
rect 1764 43036 1774 43092
rect 78194 43036 78204 43092
rect 78260 43036 80000 43092
rect 0 43008 800 43036
rect 79200 43008 80000 43036
rect 45826 42700 45836 42756
rect 45892 42700 75068 42756
rect 75124 42700 75134 42756
rect 1698 42476 1708 42532
rect 1764 42476 1774 42532
rect 46386 42476 46396 42532
rect 46452 42476 46844 42532
rect 46900 42476 77644 42532
rect 77700 42476 77710 42532
rect 0 42420 800 42448
rect 1708 42420 1764 42476
rect 79200 42420 80000 42448
rect 0 42364 1764 42420
rect 78194 42364 78204 42420
rect 78260 42364 80000 42420
rect 0 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 79200 42336 80000 42364
rect 45378 41916 45388 41972
rect 45444 41916 45948 41972
rect 46004 41916 54124 41972
rect 54180 41916 54190 41972
rect 4274 41804 4284 41860
rect 4340 41804 4844 41860
rect 4900 41804 34412 41860
rect 34468 41804 34478 41860
rect 44930 41804 44940 41860
rect 44996 41804 75292 41860
rect 75348 41804 75358 41860
rect 0 41748 800 41776
rect 79200 41748 80000 41776
rect 0 41692 1932 41748
rect 1988 41692 1998 41748
rect 78194 41692 78204 41748
rect 78260 41692 80000 41748
rect 0 41664 800 41692
rect 79200 41664 80000 41692
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 0 41076 800 41104
rect 79200 41076 80000 41104
rect 0 41020 1708 41076
rect 1764 41020 1774 41076
rect 78194 41020 78204 41076
rect 78260 41020 80000 41076
rect 0 40992 800 41020
rect 79200 40992 80000 41020
rect 2594 40908 2604 40964
rect 2660 40908 33628 40964
rect 33684 40908 33694 40964
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 4946 40460 4956 40516
rect 5012 40460 35084 40516
rect 35140 40460 35150 40516
rect 0 40404 800 40432
rect 79200 40404 80000 40432
rect 0 40348 2156 40404
rect 2212 40348 2222 40404
rect 2370 40348 2380 40404
rect 2436 40348 34412 40404
rect 34468 40348 34478 40404
rect 77746 40348 77756 40404
rect 77812 40348 80000 40404
rect 0 40320 800 40348
rect 79200 40320 80000 40348
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 78194 39900 78204 39956
rect 78260 39900 78270 39956
rect 0 39732 800 39760
rect 78204 39732 78260 39900
rect 79200 39732 80000 39760
rect 0 39676 1708 39732
rect 1764 39676 1774 39732
rect 78204 39676 80000 39732
rect 0 39648 800 39676
rect 79200 39648 80000 39676
rect 40002 39340 40012 39396
rect 40068 39340 41132 39396
rect 41188 39340 41198 39396
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 0 39060 800 39088
rect 79200 39060 80000 39088
rect 0 39004 1708 39060
rect 1764 39004 1774 39060
rect 78194 39004 78204 39060
rect 78260 39004 80000 39060
rect 0 38976 800 39004
rect 79200 38976 80000 39004
rect 2034 38892 2044 38948
rect 2100 38892 40012 38948
rect 40068 38892 40078 38948
rect 0 38388 800 38416
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 79200 38388 80000 38416
rect 0 38332 1708 38388
rect 1764 38332 2492 38388
rect 2548 38332 2558 38388
rect 78194 38332 78204 38388
rect 78260 38332 80000 38388
rect 0 38304 800 38332
rect 79200 38304 80000 38332
rect 1698 37772 1708 37828
rect 1764 37772 1774 37828
rect 0 37716 800 37744
rect 1708 37716 1764 37772
rect 79200 37716 80000 37744
rect 0 37660 1764 37716
rect 78194 37660 78204 37716
rect 78260 37660 80000 37716
rect 0 37632 800 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 79200 37632 80000 37660
rect 2034 37324 2044 37380
rect 2100 37324 43708 37380
rect 43764 37324 43774 37380
rect 2034 37100 2044 37156
rect 2100 37100 33516 37156
rect 33572 37100 33582 37156
rect 0 37044 800 37072
rect 79200 37044 80000 37072
rect 0 36988 1708 37044
rect 1764 36988 2492 37044
rect 2548 36988 2558 37044
rect 78194 36988 78204 37044
rect 78260 36988 80000 37044
rect 0 36960 800 36988
rect 79200 36960 80000 36988
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 0 36372 800 36400
rect 79200 36372 80000 36400
rect 0 36316 1708 36372
rect 1764 36316 2940 36372
rect 2996 36316 3006 36372
rect 78194 36316 78204 36372
rect 78260 36316 80000 36372
rect 0 36288 800 36316
rect 79200 36288 80000 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 0 35700 800 35728
rect 79200 35700 80000 35728
rect 0 35644 2380 35700
rect 2436 35644 2446 35700
rect 43138 35644 43148 35700
rect 43204 35644 44156 35700
rect 44212 35644 44222 35700
rect 77746 35644 77756 35700
rect 77812 35644 80000 35700
rect 0 35616 800 35644
rect 79200 35616 80000 35644
rect 40114 35532 40124 35588
rect 40180 35532 41020 35588
rect 41076 35532 41916 35588
rect 41972 35532 41982 35588
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 0 35028 800 35056
rect 79200 35028 80000 35056
rect 0 34972 1708 35028
rect 1764 34972 1774 35028
rect 78194 34972 78204 35028
rect 78260 34972 80000 35028
rect 0 34944 800 34972
rect 79200 34944 80000 34972
rect 2034 34636 2044 34692
rect 2100 34636 32620 34692
rect 32676 34636 32686 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 0 34356 800 34384
rect 79200 34356 80000 34384
rect 0 34300 1820 34356
rect 1876 34300 2492 34356
rect 2548 34300 2558 34356
rect 78194 34300 78204 34356
rect 78260 34300 80000 34356
rect 0 34272 800 34300
rect 79200 34272 80000 34300
rect 55412 34188 77868 34244
rect 77924 34188 77934 34244
rect 34178 34076 34188 34132
rect 34244 34076 34636 34132
rect 34692 34076 34702 34132
rect 55412 34020 55468 34188
rect 46610 33964 46620 34020
rect 46676 33964 47068 34020
rect 47124 33964 55468 34020
rect 0 33684 800 33712
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 79200 33684 80000 33712
rect 0 33628 1708 33684
rect 1764 33628 1774 33684
rect 78194 33628 78204 33684
rect 78260 33628 80000 33684
rect 0 33600 800 33628
rect 79200 33600 80000 33628
rect 0 33012 800 33040
rect 79200 33012 80000 33040
rect 0 32956 1708 33012
rect 1764 32956 1774 33012
rect 78194 32956 78204 33012
rect 78260 32956 80000 33012
rect 0 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 79200 32928 80000 32956
rect 2034 32620 2044 32676
rect 2100 32620 34860 32676
rect 34916 32620 34926 32676
rect 44034 32508 44044 32564
rect 44100 32508 44492 32564
rect 44548 32508 44558 32564
rect 0 32340 800 32368
rect 79200 32340 80000 32368
rect 0 32284 1708 32340
rect 1764 32284 2492 32340
rect 2548 32284 2558 32340
rect 78194 32284 78204 32340
rect 78260 32284 80000 32340
rect 0 32256 800 32284
rect 79200 32256 80000 32284
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 4274 31724 4284 31780
rect 4340 31724 4844 31780
rect 4900 31724 34972 31780
rect 35028 31724 35038 31780
rect 0 31668 800 31696
rect 79200 31668 80000 31696
rect 0 31612 1708 31668
rect 1764 31612 1774 31668
rect 78194 31612 78204 31668
rect 78260 31612 80000 31668
rect 0 31584 800 31612
rect 79200 31584 80000 31612
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 1698 31164 1708 31220
rect 1764 31164 2940 31220
rect 2996 31164 3006 31220
rect 2034 31052 2044 31108
rect 2100 31052 33964 31108
rect 34020 31052 34030 31108
rect 0 30996 800 31024
rect 79200 30996 80000 31024
rect 0 30940 1932 30996
rect 1988 30940 1998 30996
rect 77746 30940 77756 30996
rect 77812 30940 80000 30996
rect 0 30912 800 30940
rect 79200 30912 80000 30940
rect 45266 30828 45276 30884
rect 45332 30828 75292 30884
rect 75348 30828 75358 30884
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 0 30324 800 30352
rect 79200 30324 80000 30352
rect 0 30268 2380 30324
rect 2436 30268 2446 30324
rect 77970 30268 77980 30324
rect 78036 30268 80000 30324
rect 0 30240 800 30268
rect 79200 30240 80000 30268
rect 4274 29932 4284 29988
rect 4340 29932 4844 29988
rect 4900 29932 35868 29988
rect 35924 29932 35934 29988
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 0 29652 800 29680
rect 79200 29652 80000 29680
rect 0 29596 2492 29652
rect 2548 29596 2558 29652
rect 78418 29596 78428 29652
rect 78484 29596 80000 29652
rect 0 29568 800 29596
rect 79200 29568 80000 29596
rect 1698 29148 1708 29204
rect 1764 29148 1774 29204
rect 0 28980 800 29008
rect 1708 28980 1764 29148
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 79200 28980 80000 29008
rect 0 28924 1764 28980
rect 78194 28924 78204 28980
rect 78260 28924 80000 28980
rect 0 28896 800 28924
rect 79200 28896 80000 28924
rect 4274 28588 4284 28644
rect 4340 28588 4844 28644
rect 4900 28588 38780 28644
rect 38836 28588 38846 28644
rect 0 28308 800 28336
rect 79200 28308 80000 28336
rect 0 28252 1932 28308
rect 1988 28252 1998 28308
rect 78194 28252 78204 28308
rect 78260 28252 80000 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 79200 28224 80000 28252
rect 0 27636 800 27664
rect 79200 27636 80000 27664
rect 0 27580 1708 27636
rect 1764 27580 1774 27636
rect 78194 27580 78204 27636
rect 78260 27580 80000 27636
rect 0 27552 800 27580
rect 79200 27552 80000 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 77186 27132 77196 27188
rect 77252 27132 78204 27188
rect 78260 27132 78270 27188
rect 45378 27020 45388 27076
rect 45444 27020 77868 27076
rect 77924 27020 77934 27076
rect 0 26964 800 26992
rect 79200 26964 80000 26992
rect 0 26908 1708 26964
rect 1764 26908 1774 26964
rect 77532 26908 80000 26964
rect 0 26880 800 26908
rect 77532 26852 77588 26908
rect 79200 26880 80000 26908
rect 77522 26796 77532 26852
rect 77588 26796 77598 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 0 26292 800 26320
rect 79200 26292 80000 26320
rect 0 26236 2156 26292
rect 2212 26236 2222 26292
rect 78194 26236 78204 26292
rect 78260 26236 80000 26292
rect 0 26208 800 26236
rect 79200 26208 80000 26236
rect 44930 26124 44940 26180
rect 44996 26124 75292 26180
rect 75348 26124 75358 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 0 25620 800 25648
rect 79200 25620 80000 25648
rect 0 25564 1708 25620
rect 1764 25564 1774 25620
rect 77970 25564 77980 25620
rect 78036 25564 80000 25620
rect 0 25536 800 25564
rect 79200 25536 80000 25564
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 1698 25004 1708 25060
rect 1764 25004 1774 25060
rect 0 24948 800 24976
rect 1708 24948 1764 25004
rect 79200 24948 80000 24976
rect 0 24892 1764 24948
rect 77970 24892 77980 24948
rect 78036 24892 80000 24948
rect 0 24864 800 24892
rect 79200 24864 80000 24892
rect 45042 24556 45052 24612
rect 45108 24556 75292 24612
rect 75348 24556 75740 24612
rect 75796 24556 75806 24612
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 79200 24276 80000 24304
rect 0 24220 1708 24276
rect 1764 24220 1774 24276
rect 78194 24220 78204 24276
rect 78260 24220 80000 24276
rect 0 24192 800 24220
rect 79200 24192 80000 24220
rect 1698 23660 1708 23716
rect 1764 23660 1774 23716
rect 0 23604 800 23632
rect 1708 23604 1764 23660
rect 79200 23604 80000 23632
rect 0 23548 1764 23604
rect 77746 23548 77756 23604
rect 77812 23548 80000 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 79200 23520 80000 23548
rect 41682 22988 41692 23044
rect 41748 22988 75292 23044
rect 75348 22988 75740 23044
rect 75796 22988 75806 23044
rect 0 22932 800 22960
rect 79200 22932 80000 22960
rect 0 22876 1708 22932
rect 1764 22876 1774 22932
rect 77970 22876 77980 22932
rect 78036 22876 80000 22932
rect 0 22848 800 22876
rect 79200 22848 80000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 4274 22316 4284 22372
rect 4340 22316 4844 22372
rect 4900 22316 34076 22372
rect 34132 22316 34142 22372
rect 0 22260 800 22288
rect 79200 22260 80000 22288
rect 0 22204 1708 22260
rect 1764 22204 2940 22260
rect 2996 22204 3006 22260
rect 78194 22204 78204 22260
rect 78260 22204 80000 22260
rect 0 22176 800 22204
rect 79200 22176 80000 22204
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 2034 21644 2044 21700
rect 2100 21644 33628 21700
rect 33684 21644 33694 21700
rect 0 21588 800 21616
rect 79200 21588 80000 21616
rect 0 21532 1932 21588
rect 1988 21532 1998 21588
rect 77970 21532 77980 21588
rect 78036 21532 80000 21588
rect 0 21504 800 21532
rect 79200 21504 80000 21532
rect 40338 21420 40348 21476
rect 40404 21420 75292 21476
rect 75348 21420 75358 21476
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 0 20916 800 20944
rect 79200 20916 80000 20944
rect 0 20860 2380 20916
rect 2436 20860 2446 20916
rect 77634 20860 77644 20916
rect 77700 20860 78204 20916
rect 78260 20860 80000 20916
rect 0 20832 800 20860
rect 79200 20832 80000 20860
rect 40898 20524 40908 20580
rect 40964 20524 77868 20580
rect 77924 20524 77934 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 0 20244 800 20272
rect 79200 20244 80000 20272
rect 0 20188 1708 20244
rect 1764 20188 1774 20244
rect 77980 20188 80000 20244
rect 0 20160 800 20188
rect 77980 20132 78036 20188
rect 79200 20160 80000 20188
rect 2034 20076 2044 20132
rect 2100 20076 34524 20132
rect 34580 20076 34590 20132
rect 77970 20076 77980 20132
rect 78036 20076 78046 20132
rect 46050 19852 46060 19908
rect 46116 19852 75292 19908
rect 75348 19852 75358 19908
rect 0 19572 800 19600
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 0 19516 1708 19572
rect 1764 19516 2492 19572
rect 2548 19516 2558 19572
rect 0 19488 800 19516
rect 79200 19488 80000 19600
rect 1698 18956 1708 19012
rect 1764 18956 1774 19012
rect 0 18900 800 18928
rect 1708 18900 1764 18956
rect 0 18844 1764 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 79200 18816 80000 18928
rect 0 18228 800 18256
rect 0 18172 1708 18228
rect 1764 18172 1774 18228
rect 0 18144 800 18172
rect 79200 18144 80000 18256
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 0 17556 800 17584
rect 0 17500 1708 17556
rect 1764 17500 1774 17556
rect 0 17472 800 17500
rect 79200 17472 80000 17584
rect 4274 17388 4284 17444
rect 4340 17388 4844 17444
rect 4900 17388 34412 17444
rect 34468 17388 34478 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 1698 17052 1708 17108
rect 1764 17052 2940 17108
rect 2996 17052 3006 17108
rect 0 16884 800 16912
rect 0 16828 1932 16884
rect 1988 16828 1998 16884
rect 0 16800 800 16828
rect 79200 16800 80000 16912
rect 2034 16716 2044 16772
rect 2100 16716 44380 16772
rect 44436 16716 44446 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 0 16212 800 16240
rect 0 16156 2380 16212
rect 2436 16156 2446 16212
rect 0 16128 800 16156
rect 79200 16128 80000 16240
rect 1698 15820 1708 15876
rect 1764 15820 1774 15876
rect 1708 15652 1764 15820
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 924 15596 1764 15652
rect 0 15540 800 15568
rect 924 15540 980 15596
rect 0 15484 980 15540
rect 0 15456 800 15484
rect 79200 15456 80000 15568
rect 0 14868 800 14896
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 0 14812 1708 14868
rect 1764 14812 1774 14868
rect 0 14784 800 14812
rect 79200 14784 80000 14896
rect 1698 14252 1708 14308
rect 1764 14252 1774 14308
rect 0 14196 800 14224
rect 1708 14196 1764 14252
rect 0 14140 1764 14196
rect 0 14112 800 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 79200 14112 80000 14224
rect 0 13524 800 13552
rect 0 13468 1708 13524
rect 1764 13468 1774 13524
rect 0 13440 800 13468
rect 79200 13440 80000 13552
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 0 12852 800 12880
rect 0 12796 1708 12852
rect 1764 12796 1774 12852
rect 0 12768 800 12796
rect 79200 12768 80000 12880
rect 4274 12684 4284 12740
rect 4340 12684 4844 12740
rect 4900 12684 33404 12740
rect 33460 12684 33470 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 0 12180 800 12208
rect 0 12124 1932 12180
rect 1988 12124 1998 12180
rect 0 12096 800 12124
rect 79200 12096 80000 12208
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 79200 11424 80000 11536
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 79200 10752 80000 10864
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 79200 10080 80000 10192
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 79200 9408 80000 9520
rect 79200 8736 80000 8848
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 79200 8064 80000 8176
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 79200 7392 80000 7504
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 35074 6748 35084 6804
rect 35140 6748 35980 6804
rect 36036 6748 36046 6804
rect 79200 6720 80000 6832
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 79200 6048 80000 6160
rect 44482 5852 44492 5908
rect 44548 5852 46396 5908
rect 46452 5852 46462 5908
rect 40450 5628 40460 5684
rect 40516 5628 42476 5684
rect 42532 5628 42542 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 79200 5376 80000 5488
rect 39554 5180 39564 5236
rect 39620 5180 43148 5236
rect 43204 5180 43708 5236
rect 43764 5180 43774 5236
rect 42466 5068 42476 5124
rect 42532 5068 43260 5124
rect 43316 5068 43326 5124
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 79200 4704 80000 4816
rect 45042 4396 45052 4452
rect 45108 4396 46172 4452
rect 46228 4396 46238 4452
rect 29586 4172 29596 4228
rect 29652 4172 30156 4228
rect 30212 4172 39788 4228
rect 39844 4172 39854 4228
rect 43586 4172 43596 4228
rect 43652 4172 51660 4228
rect 51716 4172 51726 4228
rect 43138 4060 43148 4116
rect 43204 4060 44268 4116
rect 44324 4060 44334 4116
rect 51762 4060 51772 4116
rect 51828 4060 53004 4116
rect 53060 4060 53070 4116
rect 79200 4032 80000 4144
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 42354 3612 42364 3668
rect 42420 3612 44604 3668
rect 44660 3612 44670 3668
rect 50418 3612 50428 3668
rect 50484 3612 52220 3668
rect 52276 3612 52286 3668
rect 27234 3500 27244 3556
rect 27300 3500 28252 3556
rect 28308 3500 28318 3556
rect 28802 3500 28812 3556
rect 28868 3500 38332 3556
rect 38388 3500 38398 3556
rect 41682 3500 41692 3556
rect 41748 3500 42140 3556
rect 42196 3500 42206 3556
rect 43474 3500 43484 3556
rect 43540 3500 50876 3556
rect 50932 3500 51212 3556
rect 51268 3500 51278 3556
rect 26786 3388 26796 3444
rect 26852 3388 27580 3444
rect 27636 3388 27646 3444
rect 27794 3388 27804 3444
rect 27860 3388 38892 3444
rect 38948 3388 38958 3444
rect 42802 3388 42812 3444
rect 42868 3388 43820 3444
rect 43876 3388 43886 3444
rect 44370 3388 44380 3444
rect 44436 3388 46732 3444
rect 46788 3388 46798 3444
rect 79200 3360 80000 3472
rect 46386 3276 46396 3332
rect 46452 3276 47404 3332
rect 47460 3276 47470 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 79200 2688 80000 2800
rect 79200 2016 80000 2128
rect 79200 1344 80000 1456
rect 79200 672 80000 784
rect 79200 0 80000 112
<< via3 >>
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 76076 35488 76892
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 76860 50848 76892
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 76076 66208 76892
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _000_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33712 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46256 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _166_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46816 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _167_
timestamp 1698431365
transform -1 0 43344 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _168_
timestamp 1698431365
transform -1 0 40320 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _169_
timestamp 1698431365
transform -1 0 41216 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _170_
timestamp 1698431365
transform -1 0 45584 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _171_
timestamp 1698431365
transform 1 0 38192 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _172_
timestamp 1698431365
transform 1 0 39648 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _173_
timestamp 1698431365
transform -1 0 40992 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _174_
timestamp 1698431365
transform 1 0 33712 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _175_
timestamp 1698431365
transform 1 0 35168 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _176_
timestamp 1698431365
transform -1 0 46592 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _177_
timestamp 1698431365
transform 1 0 34496 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _178_
timestamp 1698431365
transform 1 0 43008 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _179_
timestamp 1698431365
transform 1 0 35728 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _180_
timestamp 1698431365
transform 1 0 32704 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _181_
timestamp 1698431365
transform -1 0 44240 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _182_
timestamp 1698431365
transform 1 0 39088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _183_
timestamp 1698431365
transform -1 0 44016 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _184_
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _185_
timestamp 1698431365
transform 1 0 33824 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _186_
timestamp 1698431365
transform -1 0 45584 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _187_
timestamp 1698431365
transform 1 0 34272 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _188_
timestamp 1698431365
transform -1 0 41664 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _189_
timestamp 1698431365
transform -1 0 45808 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _190_
timestamp 1698431365
transform 1 0 34384 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _191_
timestamp 1698431365
transform 1 0 34832 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _192_
timestamp 1698431365
transform 1 0 43904 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _193_
timestamp 1698431365
transform 1 0 40992 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _194_
timestamp 1698431365
transform -1 0 43568 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _195_
timestamp 1698431365
transform 1 0 34272 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _196_
timestamp 1698431365
transform 1 0 35728 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _197_
timestamp 1698431365
transform -1 0 45584 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _198_
timestamp 1698431365
transform 1 0 38192 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__000__I test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 33712 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__I
timestamp 1698431365
transform 1 0 47152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__I
timestamp 1698431365
transform 1 0 47040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__I
timestamp 1698431365
transform 1 0 43568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__I
timestamp 1698431365
transform 1 0 40992 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__I
timestamp 1698431365
transform -1 0 41664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__I
timestamp 1698431365
transform -1 0 46032 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__I
timestamp 1698431365
transform -1 0 38192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I
timestamp 1698431365
transform -1 0 39648 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__I
timestamp 1698431365
transform 1 0 40992 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__I
timestamp 1698431365
transform 1 0 33488 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I
timestamp 1698431365
transform 1 0 34944 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__I
timestamp 1698431365
transform 1 0 46816 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1698431365
transform -1 0 34496 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1698431365
transform 1 0 44128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I
timestamp 1698431365
transform 1 0 35504 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I
timestamp 1698431365
transform -1 0 32704 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1698431365
transform 1 0 44464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I
timestamp 1698431365
transform 1 0 38864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I
timestamp 1698431365
transform -1 0 44464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__I
timestamp 1698431365
transform -1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I
timestamp 1698431365
transform 1 0 33600 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1698431365
transform -1 0 46032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__I
timestamp 1698431365
transform -1 0 34272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__I
timestamp 1698431365
transform -1 0 42112 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I
timestamp 1698431365
transform -1 0 46256 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__I
timestamp 1698431365
transform 1 0 34160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__I
timestamp 1698431365
transform -1 0 34832 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__I
timestamp 1698431365
transform 1 0 43680 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__I
timestamp 1698431365
transform -1 0 40096 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I
timestamp 1698431365
transform -1 0 44016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__I
timestamp 1698431365
transform 1 0 34048 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I
timestamp 1698431365
transform 1 0 35504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I
timestamp 1698431365
transform 1 0 45808 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__I
timestamp 1698431365
transform 1 0 37968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 41776 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 41216 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 77280 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 37296 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 34384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 77728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 2912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 2464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 77728 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 2912 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 43120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 28224 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 47152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 26880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 47824 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 77728 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 27328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 77728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 55664 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 44016 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 2464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 2464 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 54320 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 2912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 56784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 50848 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 22960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 2464 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 2912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1698431365
transform 1 0 77504 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1698431365
transform 1 0 75264 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output37_I
timestamp 1698431365
transform -1 0 75488 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output38_I
timestamp 1698431365
transform 1 0 4704 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output39_I
timestamp 1698431365
transform 1 0 51632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output40_I
timestamp 1698431365
transform 1 0 25424 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output41_I
timestamp 1698431365
transform -1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output42_I
timestamp 1698431365
transform 1 0 50848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output43_I
timestamp 1698431365
transform 1 0 30128 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output44_I
timestamp 1698431365
transform 1 0 58464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output45_I
timestamp 1698431365
transform 1 0 51632 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output46_I
timestamp 1698431365
transform 1 0 43232 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output47_I
timestamp 1698431365
transform 1 0 42448 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output48_I
timestamp 1698431365
transform 1 0 75264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output49_I
timestamp 1698431365
transform 1 0 40992 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output50_I
timestamp 1698431365
transform -1 0 40432 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output51_I
timestamp 1698431365
transform 1 0 75264 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output52_I
timestamp 1698431365
transform -1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output53_I
timestamp 1698431365
transform -1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output54_I
timestamp 1698431365
transform 1 0 75264 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output55_I
timestamp 1698431365
transform -1 0 4928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output56_I
timestamp 1698431365
transform -1 0 75488 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output57_I
timestamp 1698431365
transform -1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output58_I
timestamp 1698431365
transform 1 0 43232 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output59_I
timestamp 1698431365
transform -1 0 75488 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output60_I
timestamp 1698431365
transform 1 0 36848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output61_I
timestamp 1698431365
transform 1 0 31696 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output62_I
timestamp 1698431365
transform 1 0 75264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output63_I
timestamp 1698431365
transform 1 0 75264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output64_I
timestamp 1698431365
transform -1 0 50176 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output65_I
timestamp 1698431365
transform -1 0 4928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output66_I
timestamp 1698431365
transform -1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output67_I
timestamp 1698431365
transform 1 0 36624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output68_I
timestamp 1698431365
transform -1 0 51184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output69_I
timestamp 1698431365
transform -1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_70 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 77952 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_71
timestamp 1698431365
transform 1 0 77952 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_72
timestamp 1698431365
transform -1 0 56000 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_73
timestamp 1698431365
transform -1 0 25536 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_74
timestamp 1698431365
transform 1 0 77504 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_75
timestamp 1698431365
transform -1 0 33488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_76
timestamp 1698431365
transform 1 0 77952 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_77
timestamp 1698431365
transform 1 0 77952 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_78
timestamp 1698431365
transform 1 0 77952 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_79
timestamp 1698431365
transform -1 0 32816 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_80
timestamp 1698431365
transform -1 0 31472 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_81
timestamp 1698431365
transform -1 0 2016 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_82
timestamp 1698431365
transform 1 0 77952 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_83
timestamp 1698431365
transform 1 0 77952 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_84
timestamp 1698431365
transform 1 0 77504 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_85
timestamp 1698431365
transform 1 0 77952 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_86
timestamp 1698431365
transform 1 0 77504 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_87
timestamp 1698431365
transform 1 0 77952 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_88
timestamp 1698431365
transform 1 0 50400 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_89
timestamp 1698431365
transform 1 0 77952 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_90
timestamp 1698431365
transform -1 0 46256 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_91
timestamp 1698431365
transform 1 0 77952 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_92
timestamp 1698431365
transform -1 0 2464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_93
timestamp 1698431365
transform -1 0 2016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_94
timestamp 1698431365
transform -1 0 2016 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_95
timestamp 1698431365
transform 1 0 77952 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_96
timestamp 1698431365
transform -1 0 40880 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_97
timestamp 1698431365
transform -1 0 2016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_98
timestamp 1698431365
transform -1 0 38864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_99
timestamp 1698431365
transform 1 0 77952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_100
timestamp 1698431365
transform -1 0 56448 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_101
timestamp 1698431365
transform -1 0 2016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_102
timestamp 1698431365
transform -1 0 26096 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_103
timestamp 1698431365
transform -1 0 23408 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_104
timestamp 1698431365
transform -1 0 27328 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_105
timestamp 1698431365
transform -1 0 31360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_106
timestamp 1698431365
transform 1 0 77952 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_107
timestamp 1698431365
transform -1 0 47712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_108
timestamp 1698431365
transform 1 0 77952 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_109
timestamp 1698431365
transform -1 0 48272 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_110
timestamp 1698431365
transform -1 0 2016 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_111
timestamp 1698431365
transform -1 0 42224 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_112
timestamp 1698431365
transform 1 0 77504 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_113
timestamp 1698431365
transform -1 0 2016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_114
timestamp 1698431365
transform 1 0 77952 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_115
timestamp 1698431365
transform -1 0 2016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_116
timestamp 1698431365
transform 1 0 77952 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_117
timestamp 1698431365
transform -1 0 2016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_118
timestamp 1698431365
transform 1 0 77504 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_119
timestamp 1698431365
transform -1 0 2016 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_120
timestamp 1698431365
transform -1 0 57680 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_121
timestamp 1698431365
transform 1 0 77952 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_122
timestamp 1698431365
transform 1 0 77952 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_123
timestamp 1698431365
transform -1 0 40208 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_124
timestamp 1698431365
transform 1 0 77952 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_125
timestamp 1698431365
transform -1 0 50288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_126
timestamp 1698431365
transform -1 0 32816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_127
timestamp 1698431365
transform -1 0 48608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_128
timestamp 1698431365
transform -1 0 45584 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_129
timestamp 1698431365
transform -1 0 2464 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_130
timestamp 1698431365
transform -1 0 30128 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_131
timestamp 1698431365
transform -1 0 2016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_132
timestamp 1698431365
transform -1 0 49616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_133
timestamp 1698431365
transform -1 0 38192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_134
timestamp 1698431365
transform 1 0 77952 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_135
timestamp 1698431365
transform 1 0 77952 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_136
timestamp 1698431365
transform -1 0 2016 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_137
timestamp 1698431365
transform -1 0 43792 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_138
timestamp 1698431365
transform -1 0 2016 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_139
timestamp 1698431365
transform -1 0 39424 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_140
timestamp 1698431365
transform -1 0 49056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_141
timestamp 1698431365
transform -1 0 35504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_142
timestamp 1698431365
transform -1 0 33488 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_143
timestamp 1698431365
transform -1 0 36848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_144
timestamp 1698431365
transform 1 0 77952 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_145
timestamp 1698431365
transform -1 0 46480 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_146
timestamp 1698431365
transform -1 0 56336 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_147
timestamp 1698431365
transform -1 0 37520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_148
timestamp 1698431365
transform 1 0 77952 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_149
timestamp 1698431365
transform -1 0 2016 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_150
timestamp 1698431365
transform -1 0 36288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_151
timestamp 1698431365
transform 1 0 77280 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_152
timestamp 1698431365
transform 1 0 77952 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_153
timestamp 1698431365
transform 1 0 23744 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_154
timestamp 1698431365
transform 1 0 51856 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_155
timestamp 1698431365
transform 1 0 77952 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_156
timestamp 1698431365
transform -1 0 46928 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_157
timestamp 1698431365
transform -1 0 48160 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_158
timestamp 1698431365
transform -1 0 34832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_159
timestamp 1698431365
transform -1 0 26768 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_160
timestamp 1698431365
transform -1 0 45024 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_161
timestamp 1698431365
transform -1 0 2016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_162
timestamp 1698431365
transform 1 0 77952 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_163
timestamp 1698431365
transform -1 0 38192 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_164
timestamp 1698431365
transform -1 0 2016 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_165
timestamp 1698431365
transform -1 0 2016 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_166
timestamp 1698431365
transform -1 0 44576 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_167
timestamp 1698431365
transform 1 0 77952 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_168
timestamp 1698431365
transform -1 0 2016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_169
timestamp 1698431365
transform -1 0 58352 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_170
timestamp 1698431365
transform 1 0 77952 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_171
timestamp 1698431365
transform -1 0 35504 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_172
timestamp 1698431365
transform -1 0 2016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_173
timestamp 1698431365
transform -1 0 2016 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_174
timestamp 1698431365
transform -1 0 2016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_175
timestamp 1698431365
transform -1 0 36960 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_176
timestamp 1698431365
transform -1 0 2464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_177
timestamp 1698431365
transform -1 0 2016 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_178
timestamp 1698431365
transform -1 0 2016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_179
timestamp 1698431365
transform -1 0 2016 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_180
timestamp 1698431365
transform -1 0 2016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_181
timestamp 1698431365
transform -1 0 2016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_182
timestamp 1698431365
transform -1 0 2016 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_183
timestamp 1698431365
transform -1 0 2688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_184
timestamp 1698431365
transform -1 0 2688 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_185
timestamp 1698431365
transform -1 0 2016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_186
timestamp 1698431365
transform -1 0 2016 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_187
timestamp 1698431365
transform -1 0 2016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_188
timestamp 1698431365
transform -1 0 2016 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_189
timestamp 1698431365
transform -1 0 2016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_190
timestamp 1698431365
transform -1 0 2016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_191
timestamp 1698431365
transform -1 0 2016 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_192
timestamp 1698431365
transform -1 0 2464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_193
timestamp 1698431365
transform -1 0 2016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_194
timestamp 1698431365
transform -1 0 2016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_195
timestamp 1698431365
transform -1 0 2016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_196
timestamp 1698431365
transform -1 0 2464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_197
timestamp 1698431365
transform -1 0 2016 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_198
timestamp 1698431365
transform -1 0 2016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_199
timestamp 1698431365
transform -1 0 2016 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_200
timestamp 1698431365
transform -1 0 2016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_201
timestamp 1698431365
transform -1 0 2016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_202
timestamp 1698431365
transform -1 0 2016 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_203
timestamp 1698431365
transform -1 0 2016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_204
timestamp 1698431365
transform -1 0 2016 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_205
timestamp 1698431365
transform -1 0 2688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_206
timestamp 1698431365
transform -1 0 2016 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  caravel_if_207
timestamp 1698431365
transform -1 0 2464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_208 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34832 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_209
timestamp 1698431365
transform 1 0 77952 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_210
timestamp 1698431365
transform -1 0 49616 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_211
timestamp 1698431365
transform 1 0 31360 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_212
timestamp 1698431365
transform 1 0 77952 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_213
timestamp 1698431365
transform 1 0 77952 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_214
timestamp 1698431365
transform -1 0 2688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_215
timestamp 1698431365
transform -1 0 29456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_216
timestamp 1698431365
transform -1 0 2016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_217
timestamp 1698431365
transform -1 0 40208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_218
timestamp 1698431365
transform 1 0 77952 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_219
timestamp 1698431365
transform 1 0 77952 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_220
timestamp 1698431365
transform -1 0 30800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_221
timestamp 1698431365
transform -1 0 2016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_222
timestamp 1698431365
transform 1 0 31360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_223
timestamp 1698431365
transform -1 0 2016 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_224
timestamp 1698431365
transform 1 0 77504 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_225
timestamp 1698431365
transform -1 0 2016 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_226
timestamp 1698431365
transform 1 0 77504 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_227
timestamp 1698431365
transform -1 0 46928 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_228
timestamp 1698431365
transform -1 0 2688 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_229
timestamp 1698431365
transform -1 0 39424 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_230
timestamp 1698431365
transform -1 0 30800 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_231
timestamp 1698431365
transform 1 0 77952 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_232
timestamp 1698431365
transform -1 0 2016 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  caravel_if_233
timestamp 1698431365
transform -1 0 30128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_206 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_222 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_228 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_240 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_251
timestamp 1698431365
transform 1 0 29456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_257
timestamp 1698431365
transform 1 0 30128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_263
timestamp 1698431365
transform 1 0 30800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_276
timestamp 1698431365
transform 1 0 32256 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_281
timestamp 1698431365
transform 1 0 32816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_287 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_299
timestamp 1698431365
transform 1 0 34832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_312
timestamp 1698431365
transform 1 0 36288 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_317
timestamp 1698431365
transform 1 0 36848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_323
timestamp 1698431365
transform 1 0 37520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_329
timestamp 1698431365
transform 1 0 38192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_335
timestamp 1698431365
transform 1 0 38864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_347
timestamp 1698431365
transform 1 0 40208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_353
timestamp 1698431365
transform 1 0 40880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_367
timestamp 1698431365
transform 1 0 42448 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_426
timestamp 1698431365
transform 1 0 49056 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_431
timestamp 1698431365
transform 1 0 49616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_437
timestamp 1698431365
transform 1 0 50288 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_470
timestamp 1698431365
transform 1 0 53984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_474
timestamp 1698431365
transform 1 0 54432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_512
timestamp 1698431365
transform 1 0 58688 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_546
timestamp 1698431365
transform 1 0 62496 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_580
timestamp 1698431365
transform 1 0 66304 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_614
timestamp 1698431365
transform 1 0 70112 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_648
timestamp 1698431365
transform 1 0 73920 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_682
timestamp 1698431365
transform 1 0 77728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_686
timestamp 1698431365
transform 1 0 78176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_228
timestamp 1698431365
transform 1 0 26880 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_255
timestamp 1698431365
transform 1 0 29904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_259
timestamp 1698431365
transform 1 0 30352 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698431365
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_286
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_288
timestamp 1698431365
transform 1 0 33600 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_315
timestamp 1698431365
transform 1 0 36624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_319
timestamp 1698431365
transform 1 0 37072 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_335
timestamp 1698431365
transform 1 0 38864 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_343
timestamp 1698431365
transform 1 0 39760 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_347
timestamp 1698431365
transform 1 0 40208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_356
timestamp 1698431365
transform 1 0 41216 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_358
timestamp 1698431365
transform 1 0 41440 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_361
timestamp 1698431365
transform 1 0 41776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_365
timestamp 1698431365
transform 1 0 42224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_369
timestamp 1698431365
transform 1 0 42672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_407
timestamp 1698431365
transform 1 0 46928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_411
timestamp 1698431365
transform 1 0 47376 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_419
timestamp 1698431365
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_438
timestamp 1698431365
transform 1 0 50400 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_444
timestamp 1698431365
transform 1 0 51072 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_448
timestamp 1698431365
transform 1 0 51520 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_477
timestamp 1698431365
transform 1 0 54768 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_485
timestamp 1698431365
transform 1 0 55664 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1698431365
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_556
timestamp 1698431365
transform 1 0 63616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_562
timestamp 1698431365
transform 1 0 64288 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_626
timestamp 1698431365
transform 1 0 71456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_632
timestamp 1698431365
transform 1 0 72128 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_664
timestamp 1698431365
transform 1 0 75712 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_680
timestamp 1698431365
transform 1 0 77504 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_349
timestamp 1698431365
transform 1 0 40432 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_365
timestamp 1698431365
transform 1 0 42224 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_373
timestamp 1698431365
transform 1 0 43120 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_376
timestamp 1698431365
transform 1 0 43456 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_384
timestamp 1698431365
transform 1 0 44352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698431365
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_521
timestamp 1698431365
transform 1 0 59696 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_527
timestamp 1698431365
transform 1 0 60368 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_591
timestamp 1698431365
transform 1 0 67536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_597
timestamp 1698431365
transform 1 0 68208 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_661
timestamp 1698431365
transform 1 0 75376 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_667
timestamp 1698431365
transform 1 0 76048 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_683
timestamp 1698431365
transform 1 0 77840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_687
timestamp 1698431365
transform 1 0 78288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_556
timestamp 1698431365
transform 1 0 63616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_562
timestamp 1698431365
transform 1 0 64288 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_626
timestamp 1698431365
transform 1 0 71456 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_632
timestamp 1698431365
transform 1 0 72128 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_664
timestamp 1698431365
transform 1 0 75712 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_680
timestamp 1698431365
transform 1 0 77504 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_521
timestamp 1698431365
transform 1 0 59696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_527
timestamp 1698431365
transform 1 0 60368 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_591
timestamp 1698431365
transform 1 0 67536 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_597
timestamp 1698431365
transform 1 0 68208 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_661
timestamp 1698431365
transform 1 0 75376 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_667
timestamp 1698431365
transform 1 0 76048 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_683
timestamp 1698431365
transform 1 0 77840 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_687
timestamp 1698431365
transform 1 0 78288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698431365
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_556
timestamp 1698431365
transform 1 0 63616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_562
timestamp 1698431365
transform 1 0 64288 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_626
timestamp 1698431365
transform 1 0 71456 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_632
timestamp 1698431365
transform 1 0 72128 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_664
timestamp 1698431365
transform 1 0 75712 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_680
timestamp 1698431365
transform 1 0 77504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_521
timestamp 1698431365
transform 1 0 59696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_527
timestamp 1698431365
transform 1 0 60368 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_591
timestamp 1698431365
transform 1 0 67536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_597
timestamp 1698431365
transform 1 0 68208 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_661
timestamp 1698431365
transform 1 0 75376 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_667
timestamp 1698431365
transform 1 0 76048 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_683
timestamp 1698431365
transform 1 0 77840 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_687
timestamp 1698431365
transform 1 0 78288 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_556
timestamp 1698431365
transform 1 0 63616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_562
timestamp 1698431365
transform 1 0 64288 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_626
timestamp 1698431365
transform 1 0 71456 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_632
timestamp 1698431365
transform 1 0 72128 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_664
timestamp 1698431365
transform 1 0 75712 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_680
timestamp 1698431365
transform 1 0 77504 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698431365
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_521
timestamp 1698431365
transform 1 0 59696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_527
timestamp 1698431365
transform 1 0 60368 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_591
timestamp 1698431365
transform 1 0 67536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_597
timestamp 1698431365
transform 1 0 68208 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_661
timestamp 1698431365
transform 1 0 75376 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_667
timestamp 1698431365
transform 1 0 76048 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_683
timestamp 1698431365
transform 1 0 77840 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_687
timestamp 1698431365
transform 1 0 78288 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698431365
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_556
timestamp 1698431365
transform 1 0 63616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_562
timestamp 1698431365
transform 1 0 64288 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_626
timestamp 1698431365
transform 1 0 71456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_632
timestamp 1698431365
transform 1 0 72128 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_664
timestamp 1698431365
transform 1 0 75712 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_680
timestamp 1698431365
transform 1 0 77504 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698431365
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_521
timestamp 1698431365
transform 1 0 59696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_527
timestamp 1698431365
transform 1 0 60368 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_591
timestamp 1698431365
transform 1 0 67536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_597
timestamp 1698431365
transform 1 0 68208 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_661
timestamp 1698431365
transform 1 0 75376 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_667
timestamp 1698431365
transform 1 0 76048 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_683
timestamp 1698431365
transform 1 0 77840 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_687
timestamp 1698431365
transform 1 0 78288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_6
timestamp 1698431365
transform 1 0 2016 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698431365
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_556
timestamp 1698431365
transform 1 0 63616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_562
timestamp 1698431365
transform 1 0 64288 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_626
timestamp 1698431365
transform 1 0 71456 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_632
timestamp 1698431365
transform 1 0 72128 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_664
timestamp 1698431365
transform 1 0 75712 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_680
timestamp 1698431365
transform 1 0 77504 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_28
timestamp 1698431365
transform 1 0 4480 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698431365
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_521
timestamp 1698431365
transform 1 0 59696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_527
timestamp 1698431365
transform 1 0 60368 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_591
timestamp 1698431365
transform 1 0 67536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_597
timestamp 1698431365
transform 1 0 68208 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_661
timestamp 1698431365
transform 1 0 75376 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_667
timestamp 1698431365
transform 1 0 76048 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_683
timestamp 1698431365
transform 1 0 77840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_687
timestamp 1698431365
transform 1 0 78288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_6
timestamp 1698431365
transform 1 0 2016 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698431365
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698431365
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_556
timestamp 1698431365
transform 1 0 63616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_562
timestamp 1698431365
transform 1 0 64288 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_626
timestamp 1698431365
transform 1 0 71456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_632
timestamp 1698431365
transform 1 0 72128 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_664
timestamp 1698431365
transform 1 0 75712 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_680
timestamp 1698431365
transform 1 0 77504 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_6
timestamp 1698431365
transform 1 0 2016 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_22
timestamp 1698431365
transform 1 0 3808 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_30
timestamp 1698431365
transform 1 0 4704 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_521
timestamp 1698431365
transform 1 0 59696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_527
timestamp 1698431365
transform 1 0 60368 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_591
timestamp 1698431365
transform 1 0 67536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_597
timestamp 1698431365
transform 1 0 68208 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_661
timestamp 1698431365
transform 1 0 75376 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_667
timestamp 1698431365
transform 1 0 76048 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_683
timestamp 1698431365
transform 1 0 77840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_687
timestamp 1698431365
transform 1 0 78288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_6
timestamp 1698431365
transform 1 0 2016 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698431365
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_556
timestamp 1698431365
transform 1 0 63616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_562
timestamp 1698431365
transform 1 0 64288 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_626
timestamp 1698431365
transform 1 0 71456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_632
timestamp 1698431365
transform 1 0 72128 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_664
timestamp 1698431365
transform 1 0 75712 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_680
timestamp 1698431365
transform 1 0 77504 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_6
timestamp 1698431365
transform 1 0 2016 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_22
timestamp 1698431365
transform 1 0 3808 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_30
timestamp 1698431365
transform 1 0 4704 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_521
timestamp 1698431365
transform 1 0 59696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_527
timestamp 1698431365
transform 1 0 60368 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_591
timestamp 1698431365
transform 1 0 67536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_597
timestamp 1698431365
transform 1 0 68208 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_661
timestamp 1698431365
transform 1 0 75376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_667
timestamp 1698431365
transform 1 0 76048 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_683
timestamp 1698431365
transform 1 0 77840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_687
timestamp 1698431365
transform 1 0 78288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_12
timestamp 1698431365
transform 1 0 2688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_16
timestamp 1698431365
transform 1 0 3136 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_48
timestamp 1698431365
transform 1 0 6720 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_64
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698431365
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_556
timestamp 1698431365
transform 1 0 63616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_562
timestamp 1698431365
transform 1 0 64288 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_626
timestamp 1698431365
transform 1 0 71456 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_632
timestamp 1698431365
transform 1 0 72128 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_664
timestamp 1698431365
transform 1 0 75712 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_680
timestamp 1698431365
transform 1 0 77504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_28
timestamp 1698431365
transform 1 0 4480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_521
timestamp 1698431365
transform 1 0 59696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_527
timestamp 1698431365
transform 1 0 60368 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_591
timestamp 1698431365
transform 1 0 67536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_597
timestamp 1698431365
transform 1 0 68208 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_661
timestamp 1698431365
transform 1 0 75376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_667
timestamp 1698431365
transform 1 0 76048 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_683
timestamp 1698431365
transform 1 0 77840 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_687
timestamp 1698431365
transform 1 0 78288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_6
timestamp 1698431365
transform 1 0 2016 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698431365
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698431365
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698431365
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_556
timestamp 1698431365
transform 1 0 63616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_562
timestamp 1698431365
transform 1 0 64288 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_626
timestamp 1698431365
transform 1 0 71456 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_632
timestamp 1698431365
transform 1 0 72128 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_664
timestamp 1698431365
transform 1 0 75712 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_680
timestamp 1698431365
transform 1 0 77504 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_6
timestamp 1698431365
transform 1 0 2016 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_22
timestamp 1698431365
transform 1 0 3808 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_30
timestamp 1698431365
transform 1 0 4704 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_381
timestamp 1698431365
transform 1 0 44016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698431365
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_521
timestamp 1698431365
transform 1 0 59696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_527
timestamp 1698431365
transform 1 0 60368 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_591
timestamp 1698431365
transform 1 0 67536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_597
timestamp 1698431365
transform 1 0 68208 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_661
timestamp 1698431365
transform 1 0 75376 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_667
timestamp 1698431365
transform 1 0 76048 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_683
timestamp 1698431365
transform 1 0 77840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_687
timestamp 1698431365
transform 1 0 78288 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_12
timestamp 1698431365
transform 1 0 2688 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_44
timestamp 1698431365
transform 1 0 6272 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698431365
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698431365
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_346
timestamp 1698431365
transform 1 0 40096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698431365
transform 1 0 47936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_556
timestamp 1698431365
transform 1 0 63616 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_562
timestamp 1698431365
transform 1 0 64288 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_626
timestamp 1698431365
transform 1 0 71456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_632
timestamp 1698431365
transform 1 0 72128 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_648
timestamp 1698431365
transform 1 0 73920 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_656
timestamp 1698431365
transform 1 0 74816 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_6
timestamp 1698431365
transform 1 0 2016 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_22
timestamp 1698431365
transform 1 0 3808 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_30
timestamp 1698431365
transform 1 0 4704 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_381
timestamp 1698431365
transform 1 0 44016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698431365
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_521
timestamp 1698431365
transform 1 0 59696 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_527
timestamp 1698431365
transform 1 0 60368 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_591
timestamp 1698431365
transform 1 0 67536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_597
timestamp 1698431365
transform 1 0 68208 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_661
timestamp 1698431365
transform 1 0 75376 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_667
timestamp 1698431365
transform 1 0 76048 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_675
timestamp 1698431365
transform 1 0 76944 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_679
timestamp 1698431365
transform 1 0 77392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_12
timestamp 1698431365
transform 1 0 2688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_16
timestamp 1698431365
transform 1 0 3136 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_48
timestamp 1698431365
transform 1 0 6720 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698431365
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_346
timestamp 1698431365
transform 1 0 40096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698431365
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698431365
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_556
timestamp 1698431365
transform 1 0 63616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_562
timestamp 1698431365
transform 1 0 64288 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_626
timestamp 1698431365
transform 1 0 71456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_632
timestamp 1698431365
transform 1 0 72128 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_648
timestamp 1698431365
transform 1 0 73920 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_656
timestamp 1698431365
transform 1 0 74816 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698431365
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_451
timestamp 1698431365
transform 1 0 51856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_521
timestamp 1698431365
transform 1 0 59696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_527
timestamp 1698431365
transform 1 0 60368 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_591
timestamp 1698431365
transform 1 0 67536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_597
timestamp 1698431365
transform 1 0 68208 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_661
timestamp 1698431365
transform 1 0 75376 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_667
timestamp 1698431365
transform 1 0 76048 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_683
timestamp 1698431365
transform 1 0 77840 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_6
timestamp 1698431365
transform 1 0 2016 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698431365
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_556
timestamp 1698431365
transform 1 0 63616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_562
timestamp 1698431365
transform 1 0 64288 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_626
timestamp 1698431365
transform 1 0 71456 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_632
timestamp 1698431365
transform 1 0 72128 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_648
timestamp 1698431365
transform 1 0 73920 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_656
timestamp 1698431365
transform 1 0 74816 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_6
timestamp 1698431365
transform 1 0 2016 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_22
timestamp 1698431365
transform 1 0 3808 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_30
timestamp 1698431365
transform 1 0 4704 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_381
timestamp 1698431365
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_451
timestamp 1698431365
transform 1 0 51856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_521
timestamp 1698431365
transform 1 0 59696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_527
timestamp 1698431365
transform 1 0 60368 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_591
timestamp 1698431365
transform 1 0 67536 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_597
timestamp 1698431365
transform 1 0 68208 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_661
timestamp 1698431365
transform 1 0 75376 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_667
timestamp 1698431365
transform 1 0 76048 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_675
timestamp 1698431365
transform 1 0 76944 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_679
timestamp 1698431365
transform 1 0 77392 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_6
timestamp 1698431365
transform 1 0 2016 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698431365
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_556
timestamp 1698431365
transform 1 0 63616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_562
timestamp 1698431365
transform 1 0 64288 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_626
timestamp 1698431365
transform 1 0 71456 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_632
timestamp 1698431365
transform 1 0 72128 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_648
timestamp 1698431365
transform 1 0 73920 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_656
timestamp 1698431365
transform 1 0 74816 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_6
timestamp 1698431365
transform 1 0 2016 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_22
timestamp 1698431365
transform 1 0 3808 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_30
timestamp 1698431365
transform 1 0 4704 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698431365
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_521
timestamp 1698431365
transform 1 0 59696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_527
timestamp 1698431365
transform 1 0 60368 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_591
timestamp 1698431365
transform 1 0 67536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_597
timestamp 1698431365
transform 1 0 68208 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_661
timestamp 1698431365
transform 1 0 75376 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_667
timestamp 1698431365
transform 1 0 76048 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_683
timestamp 1698431365
transform 1 0 77840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_687
timestamp 1698431365
transform 1 0 78288 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_6
timestamp 1698431365
transform 1 0 2016 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_416
timestamp 1698431365
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698431365
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_556
timestamp 1698431365
transform 1 0 63616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_562
timestamp 1698431365
transform 1 0 64288 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_626
timestamp 1698431365
transform 1 0 71456 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_632
timestamp 1698431365
transform 1 0 72128 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_648
timestamp 1698431365
transform 1 0 73920 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_656
timestamp 1698431365
transform 1 0 74816 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_10
timestamp 1698431365
transform 1 0 2464 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_381
timestamp 1698431365
transform 1 0 44016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698431365
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_521
timestamp 1698431365
transform 1 0 59696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_527
timestamp 1698431365
transform 1 0 60368 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_591
timestamp 1698431365
transform 1 0 67536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_597
timestamp 1698431365
transform 1 0 68208 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_661
timestamp 1698431365
transform 1 0 75376 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_667
timestamp 1698431365
transform 1 0 76048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_675
timestamp 1698431365
transform 1 0 76944 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_6
timestamp 1698431365
transform 1 0 2016 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698431365
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_556
timestamp 1698431365
transform 1 0 63616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_562
timestamp 1698431365
transform 1 0 64288 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_626
timestamp 1698431365
transform 1 0 71456 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_632
timestamp 1698431365
transform 1 0 72128 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_664
timestamp 1698431365
transform 1 0 75712 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_680
timestamp 1698431365
transform 1 0 77504 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_28
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_381
timestamp 1698431365
transform 1 0 44016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698431365
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_521
timestamp 1698431365
transform 1 0 59696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_527
timestamp 1698431365
transform 1 0 60368 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_591
timestamp 1698431365
transform 1 0 67536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_597
timestamp 1698431365
transform 1 0 68208 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_661
timestamp 1698431365
transform 1 0 75376 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_667
timestamp 1698431365
transform 1 0 76048 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_683
timestamp 1698431365
transform 1 0 77840 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_6
timestamp 1698431365
transform 1 0 2016 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698431365
transform 1 0 47936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_556
timestamp 1698431365
transform 1 0 63616 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_562
timestamp 1698431365
transform 1 0 64288 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_626
timestamp 1698431365
transform 1 0 71456 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_632
timestamp 1698431365
transform 1 0 72128 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_664
timestamp 1698431365
transform 1 0 75712 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_680
timestamp 1698431365
transform 1 0 77504 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_28
timestamp 1698431365
transform 1 0 4480 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_32
timestamp 1698431365
transform 1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698431365
transform 1 0 44016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698431365
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_521
timestamp 1698431365
transform 1 0 59696 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_527
timestamp 1698431365
transform 1 0 60368 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_591
timestamp 1698431365
transform 1 0 67536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_597
timestamp 1698431365
transform 1 0 68208 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_661
timestamp 1698431365
transform 1 0 75376 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_667
timestamp 1698431365
transform 1 0 76048 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_683
timestamp 1698431365
transform 1 0 77840 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_12
timestamp 1698431365
transform 1 0 2688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_16
timestamp 1698431365
transform 1 0 3136 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_48
timestamp 1698431365
transform 1 0 6720 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_64
timestamp 1698431365
transform 1 0 8512 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_68
timestamp 1698431365
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698431365
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_416
timestamp 1698431365
transform 1 0 47936 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698431365
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_556
timestamp 1698431365
transform 1 0 63616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_562
timestamp 1698431365
transform 1 0 64288 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_626
timestamp 1698431365
transform 1 0 71456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_632
timestamp 1698431365
transform 1 0 72128 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_648
timestamp 1698431365
transform 1 0 73920 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_656
timestamp 1698431365
transform 1 0 74816 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_28
timestamp 1698431365
transform 1 0 4480 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_32
timestamp 1698431365
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_381
timestamp 1698431365
transform 1 0 44016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1698431365
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_521
timestamp 1698431365
transform 1 0 59696 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_527
timestamp 1698431365
transform 1 0 60368 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_591
timestamp 1698431365
transform 1 0 67536 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_597
timestamp 1698431365
transform 1 0 68208 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_661
timestamp 1698431365
transform 1 0 75376 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_667
timestamp 1698431365
transform 1 0 76048 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_675
timestamp 1698431365
transform 1 0 76944 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_679
timestamp 1698431365
transform 1 0 77392 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_8
timestamp 1698431365
transform 1 0 2240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_12
timestamp 1698431365
transform 1 0 2688 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_44
timestamp 1698431365
transform 1 0 6272 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_60
timestamp 1698431365
transform 1 0 8064 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_68
timestamp 1698431365
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_368
timestamp 1698431365
transform 1 0 42560 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_372
timestamp 1698431365
transform 1 0 43008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_374
timestamp 1698431365
transform 1 0 43232 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_383
timestamp 1698431365
transform 1 0 44240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_387
timestamp 1698431365
transform 1 0 44688 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1698431365
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698431365
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_556
timestamp 1698431365
transform 1 0 63616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_562
timestamp 1698431365
transform 1 0 64288 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_626
timestamp 1698431365
transform 1 0 71456 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_632
timestamp 1698431365
transform 1 0 72128 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_664
timestamp 1698431365
transform 1 0 75712 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_680
timestamp 1698431365
transform 1 0 77504 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_6
timestamp 1698431365
transform 1 0 2016 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_22
timestamp 1698431365
transform 1 0 3808 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_30
timestamp 1698431365
transform 1 0 4704 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_333
timestamp 1698431365
transform 1 0 38640 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_341
timestamp 1698431365
transform 1 0 39536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_345
timestamp 1698431365
transform 1 0 39984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_347
timestamp 1698431365
transform 1 0 40208 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_356
timestamp 1698431365
transform 1 0 41216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_360
timestamp 1698431365
transform 1 0 41664 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_376
timestamp 1698431365
transform 1 0 43456 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_384
timestamp 1698431365
transform 1 0 44352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_451
timestamp 1698431365
transform 1 0 51856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_521
timestamp 1698431365
transform 1 0 59696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_527
timestamp 1698431365
transform 1 0 60368 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_591
timestamp 1698431365
transform 1 0 67536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_597
timestamp 1698431365
transform 1 0 68208 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_661
timestamp 1698431365
transform 1 0 75376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_667
timestamp 1698431365
transform 1 0 76048 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_683
timestamp 1698431365
transform 1 0 77840 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_6
timestamp 1698431365
transform 1 0 2016 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_290
timestamp 1698431365
transform 1 0 33824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_292
timestamp 1698431365
transform 1 0 34048 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_303
timestamp 1698431365
transform 1 0 35280 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_335
timestamp 1698431365
transform 1 0 38864 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_343
timestamp 1698431365
transform 1 0 39760 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_347
timestamp 1698431365
transform 1 0 40208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_384
timestamp 1698431365
transform 1 0 44352 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_392
timestamp 1698431365
transform 1 0 45248 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_396
timestamp 1698431365
transform 1 0 45696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_406
timestamp 1698431365
transform 1 0 46816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_410
timestamp 1698431365
transform 1 0 47264 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_418
timestamp 1698431365
transform 1 0 48160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_556
timestamp 1698431365
transform 1 0 63616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_562
timestamp 1698431365
transform 1 0 64288 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_626
timestamp 1698431365
transform 1 0 71456 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_632
timestamp 1698431365
transform 1 0 72128 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_664
timestamp 1698431365
transform 1 0 75712 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_8
timestamp 1698431365
transform 1 0 2240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_12
timestamp 1698431365
transform 1 0 2688 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_28
timestamp 1698431365
transform 1 0 4480 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_395
timestamp 1698431365
transform 1 0 45584 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_427
timestamp 1698431365
transform 1 0 49168 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_443
timestamp 1698431365
transform 1 0 50960 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_451
timestamp 1698431365
transform 1 0 51856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_521
timestamp 1698431365
transform 1 0 59696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_527
timestamp 1698431365
transform 1 0 60368 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_591
timestamp 1698431365
transform 1 0 67536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_597
timestamp 1698431365
transform 1 0 68208 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_661
timestamp 1698431365
transform 1 0 75376 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_667
timestamp 1698431365
transform 1 0 76048 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_683
timestamp 1698431365
transform 1 0 77840 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_6
timestamp 1698431365
transform 1 0 2016 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_295
timestamp 1698431365
transform 1 0 34384 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_327
timestamp 1698431365
transform 1 0 37968 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_335
timestamp 1698431365
transform 1 0 38864 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_339
timestamp 1698431365
transform 1 0 39312 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_348
timestamp 1698431365
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_356
timestamp 1698431365
transform 1 0 41216 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_380
timestamp 1698431365
transform 1 0 43904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_384
timestamp 1698431365
transform 1 0 44352 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698431365
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698431365
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_556
timestamp 1698431365
transform 1 0 63616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_562
timestamp 1698431365
transform 1 0 64288 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_626
timestamp 1698431365
transform 1 0 71456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_632
timestamp 1698431365
transform 1 0 72128 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_664
timestamp 1698431365
transform 1 0 75712 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_680
timestamp 1698431365
transform 1 0 77504 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_12
timestamp 1698431365
transform 1 0 2688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_16
timestamp 1698431365
transform 1 0 3136 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_32
timestamp 1698431365
transform 1 0 4928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_279
timestamp 1698431365
transform 1 0 32592 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_287
timestamp 1698431365
transform 1 0 33488 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_291
timestamp 1698431365
transform 1 0 33936 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_302
timestamp 1698431365
transform 1 0 35168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_310
timestamp 1698431365
transform 1 0 36064 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698431365
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_381
timestamp 1698431365
transform 1 0 44016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_451
timestamp 1698431365
transform 1 0 51856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_521
timestamp 1698431365
transform 1 0 59696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_527
timestamp 1698431365
transform 1 0 60368 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_591
timestamp 1698431365
transform 1 0 67536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_597
timestamp 1698431365
transform 1 0 68208 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_661
timestamp 1698431365
transform 1 0 75376 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_667
timestamp 1698431365
transform 1 0 76048 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_675
timestamp 1698431365
transform 1 0 76944 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_679
timestamp 1698431365
transform 1 0 77392 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_8
timestamp 1698431365
transform 1 0 2240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_12
timestamp 1698431365
transform 1 0 2688 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_44
timestamp 1698431365
transform 1 0 6272 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_60
timestamp 1698431365
transform 1 0 8064 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_286
timestamp 1698431365
transform 1 0 33376 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_297
timestamp 1698431365
transform 1 0 34608 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_329
timestamp 1698431365
transform 1 0 38192 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_345
timestamp 1698431365
transform 1 0 39984 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698431365
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698431365
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_556
timestamp 1698431365
transform 1 0 63616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_562
timestamp 1698431365
transform 1 0 64288 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_626
timestamp 1698431365
transform 1 0 71456 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_632
timestamp 1698431365
transform 1 0 72128 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_664
timestamp 1698431365
transform 1 0 75712 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_680
timestamp 1698431365
transform 1 0 77504 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_6
timestamp 1698431365
transform 1 0 2016 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_22
timestamp 1698431365
transform 1 0 3808 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_30
timestamp 1698431365
transform 1 0 4704 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_263
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_271
timestamp 1698431365
transform 1 0 31696 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_275
timestamp 1698431365
transform 1 0 32144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_277
timestamp 1698431365
transform 1 0 32368 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_288
timestamp 1698431365
transform 1 0 33600 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_304
timestamp 1698431365
transform 1 0 35392 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_312
timestamp 1698431365
transform 1 0 36288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1698431365
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_333
timestamp 1698431365
transform 1 0 38640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_337
timestamp 1698431365
transform 1 0 39088 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_369
timestamp 1698431365
transform 1 0 42672 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698431365
transform 1 0 51856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_521
timestamp 1698431365
transform 1 0 59696 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_527
timestamp 1698431365
transform 1 0 60368 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_591
timestamp 1698431365
transform 1 0 67536 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_597
timestamp 1698431365
transform 1 0 68208 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_661
timestamp 1698431365
transform 1 0 75376 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_667
timestamp 1698431365
transform 1 0 76048 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_683
timestamp 1698431365
transform 1 0 77840 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_8
timestamp 1698431365
transform 1 0 2240 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_12
timestamp 1698431365
transform 1 0 2688 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_44
timestamp 1698431365
transform 1 0 6272 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_60
timestamp 1698431365
transform 1 0 8064 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_68
timestamp 1698431365
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_298
timestamp 1698431365
transform 1 0 34720 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_310
timestamp 1698431365
transform 1 0 36064 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_326
timestamp 1698431365
transform 1 0 37856 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_345
timestamp 1698431365
transform 1 0 39984 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_349
timestamp 1698431365
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_356
timestamp 1698431365
transform 1 0 41216 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_372
timestamp 1698431365
transform 1 0 43008 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_376
timestamp 1698431365
transform 1 0 43456 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_388
timestamp 1698431365
transform 1 0 44800 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698431365
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_556
timestamp 1698431365
transform 1 0 63616 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_562
timestamp 1698431365
transform 1 0 64288 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_626
timestamp 1698431365
transform 1 0 71456 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_632
timestamp 1698431365
transform 1 0 72128 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_664
timestamp 1698431365
transform 1 0 75712 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_680
timestamp 1698431365
transform 1 0 77504 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_6
timestamp 1698431365
transform 1 0 2016 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_22
timestamp 1698431365
transform 1 0 3808 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_30
timestamp 1698431365
transform 1 0 4704 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_333
timestamp 1698431365
transform 1 0 38640 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_341
timestamp 1698431365
transform 1 0 39536 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_343
timestamp 1698431365
transform 1 0 39760 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_362
timestamp 1698431365
transform 1 0 41888 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_378
timestamp 1698431365
transform 1 0 43680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_382
timestamp 1698431365
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_395
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_399
timestamp 1698431365
transform 1 0 46032 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_431
timestamp 1698431365
transform 1 0 49616 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_447
timestamp 1698431365
transform 1 0 51408 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_521
timestamp 1698431365
transform 1 0 59696 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_527
timestamp 1698431365
transform 1 0 60368 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_591
timestamp 1698431365
transform 1 0 67536 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_597
timestamp 1698431365
transform 1 0 68208 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_661
timestamp 1698431365
transform 1 0 75376 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_667
timestamp 1698431365
transform 1 0 76048 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_683
timestamp 1698431365
transform 1 0 77840 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_6
timestamp 1698431365
transform 1 0 2016 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_290
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_304
timestamp 1698431365
transform 1 0 35392 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_336
timestamp 1698431365
transform 1 0 38976 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_344
timestamp 1698431365
transform 1 0 39872 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_348
timestamp 1698431365
transform 1 0 40320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698431365
transform 1 0 55776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_556
timestamp 1698431365
transform 1 0 63616 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_562
timestamp 1698431365
transform 1 0 64288 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_626
timestamp 1698431365
transform 1 0 71456 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_632
timestamp 1698431365
transform 1 0 72128 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_664
timestamp 1698431365
transform 1 0 75712 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_680
timestamp 1698431365
transform 1 0 77504 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_10
timestamp 1698431365
transform 1 0 2464 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_26
timestamp 1698431365
transform 1 0 4256 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_279
timestamp 1698431365
transform 1 0 32592 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_287
timestamp 1698431365
transform 1 0 33488 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_298
timestamp 1698431365
transform 1 0 34720 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698431365
transform 1 0 51856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_521
timestamp 1698431365
transform 1 0 59696 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_527
timestamp 1698431365
transform 1 0 60368 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_591
timestamp 1698431365
transform 1 0 67536 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_597
timestamp 1698431365
transform 1 0 68208 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_661
timestamp 1698431365
transform 1 0 75376 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_667
timestamp 1698431365
transform 1 0 76048 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_675
timestamp 1698431365
transform 1 0 76944 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_679
timestamp 1698431365
transform 1 0 77392 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_28
timestamp 1698431365
transform 1 0 4480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_32
timestamp 1698431365
transform 1 0 4928 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_64
timestamp 1698431365
transform 1 0 8512 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_314
timestamp 1698431365
transform 1 0 36512 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_322
timestamp 1698431365
transform 1 0 37408 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_326
timestamp 1698431365
transform 1 0 37856 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_337
timestamp 1698431365
transform 1 0 39088 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_345
timestamp 1698431365
transform 1 0 39984 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_349
timestamp 1698431365
transform 1 0 40432 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_384
timestamp 1698431365
transform 1 0 44352 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_386
timestamp 1698431365
transform 1 0 44576 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_395
timestamp 1698431365
transform 1 0 45584 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_399
timestamp 1698431365
transform 1 0 46032 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_415
timestamp 1698431365
transform 1 0 47824 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698431365
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_486
timestamp 1698431365
transform 1 0 55776 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_556
timestamp 1698431365
transform 1 0 63616 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_562
timestamp 1698431365
transform 1 0 64288 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_626
timestamp 1698431365
transform 1 0 71456 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_632
timestamp 1698431365
transform 1 0 72128 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_664
timestamp 1698431365
transform 1 0 75712 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_680
timestamp 1698431365
transform 1 0 77504 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_6
timestamp 1698431365
transform 1 0 2016 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_22
timestamp 1698431365
transform 1 0 3808 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_30
timestamp 1698431365
transform 1 0 4704 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698431365
transform 1 0 20496 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_395
timestamp 1698431365
transform 1 0 45584 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_404
timestamp 1698431365
transform 1 0 46592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_408
timestamp 1698431365
transform 1 0 47040 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_440
timestamp 1698431365
transform 1 0 50624 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_448
timestamp 1698431365
transform 1 0 51520 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_452
timestamp 1698431365
transform 1 0 51968 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_454
timestamp 1698431365
transform 1 0 52192 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_521
timestamp 1698431365
transform 1 0 59696 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_527
timestamp 1698431365
transform 1 0 60368 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_591
timestamp 1698431365
transform 1 0 67536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_597
timestamp 1698431365
transform 1 0 68208 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_661
timestamp 1698431365
transform 1 0 75376 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_667
timestamp 1698431365
transform 1 0 76048 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_683
timestamp 1698431365
transform 1 0 77840 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_6
timestamp 1698431365
transform 1 0 2016 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_276
timestamp 1698431365
transform 1 0 32256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_346
timestamp 1698431365
transform 1 0 40096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_416
timestamp 1698431365
transform 1 0 47936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_486
timestamp 1698431365
transform 1 0 55776 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_556
timestamp 1698431365
transform 1 0 63616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_562
timestamp 1698431365
transform 1 0 64288 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_626
timestamp 1698431365
transform 1 0 71456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_632
timestamp 1698431365
transform 1 0 72128 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_664
timestamp 1698431365
transform 1 0 75712 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_680
timestamp 1698431365
transform 1 0 77504 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_6
timestamp 1698431365
transform 1 0 2016 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_22
timestamp 1698431365
transform 1 0 3808 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_30
timestamp 1698431365
transform 1 0 4704 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_279
timestamp 1698431365
transform 1 0 32592 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_287
timestamp 1698431365
transform 1 0 33488 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_291
timestamp 1698431365
transform 1 0 33936 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_302
timestamp 1698431365
transform 1 0 35168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_304
timestamp 1698431365
transform 1 0 35392 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_349
timestamp 1698431365
transform 1 0 40432 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_365
timestamp 1698431365
transform 1 0 42224 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_375
timestamp 1698431365
transform 1 0 43344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_379
timestamp 1698431365
transform 1 0 43792 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_383
timestamp 1698431365
transform 1 0 44240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_395
timestamp 1698431365
transform 1 0 45584 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_399
timestamp 1698431365
transform 1 0 46032 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_431
timestamp 1698431365
transform 1 0 49616 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_447
timestamp 1698431365
transform 1 0 51408 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_521
timestamp 1698431365
transform 1 0 59696 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_527
timestamp 1698431365
transform 1 0 60368 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_591
timestamp 1698431365
transform 1 0 67536 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_597
timestamp 1698431365
transform 1 0 68208 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_661
timestamp 1698431365
transform 1 0 75376 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_667
timestamp 1698431365
transform 1 0 76048 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_683
timestamp 1698431365
transform 1 0 77840 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_28
timestamp 1698431365
transform 1 0 4480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_32
timestamp 1698431365
transform 1 0 4928 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_64
timestamp 1698431365
transform 1 0 8512 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_276
timestamp 1698431365
transform 1 0 32256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_346
timestamp 1698431365
transform 1 0 40096 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_360
timestamp 1698431365
transform 1 0 41664 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_364
timestamp 1698431365
transform 1 0 42112 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_380
timestamp 1698431365
transform 1 0 43904 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_388
timestamp 1698431365
transform 1 0 44800 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_397
timestamp 1698431365
transform 1 0 45808 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_401
timestamp 1698431365
transform 1 0 46256 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_417
timestamp 1698431365
transform 1 0 48048 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698431365
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_486
timestamp 1698431365
transform 1 0 55776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_556
timestamp 1698431365
transform 1 0 63616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_562
timestamp 1698431365
transform 1 0 64288 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_626
timestamp 1698431365
transform 1 0 71456 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_632
timestamp 1698431365
transform 1 0 72128 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_664
timestamp 1698431365
transform 1 0 75712 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_680
timestamp 1698431365
transform 1 0 77504 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_10
timestamp 1698431365
transform 1 0 2464 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_26
timestamp 1698431365
transform 1 0 4256 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_101
timestamp 1698431365
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_241
timestamp 1698431365
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_311
timestamp 1698431365
transform 1 0 36176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_381
timestamp 1698431365
transform 1 0 44016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698431365
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_521
timestamp 1698431365
transform 1 0 59696 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_527
timestamp 1698431365
transform 1 0 60368 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_591
timestamp 1698431365
transform 1 0 67536 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_597
timestamp 1698431365
transform 1 0 68208 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_661
timestamp 1698431365
transform 1 0 75376 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_667
timestamp 1698431365
transform 1 0 76048 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_675
timestamp 1698431365
transform 1 0 76944 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_679
timestamp 1698431365
transform 1 0 77392 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_6
timestamp 1698431365
transform 1 0 2016 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_136
timestamp 1698431365
transform 1 0 16576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_206
timestamp 1698431365
transform 1 0 24416 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_276
timestamp 1698431365
transform 1 0 32256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_290
timestamp 1698431365
transform 1 0 33824 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_294
timestamp 1698431365
transform 1 0 34272 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_296
timestamp 1698431365
transform 1 0 34496 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_307
timestamp 1698431365
transform 1 0 35728 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_339
timestamp 1698431365
transform 1 0 39312 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_347
timestamp 1698431365
transform 1 0 40208 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_349
timestamp 1698431365
transform 1 0 40432 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_368
timestamp 1698431365
transform 1 0 42560 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_377
timestamp 1698431365
transform 1 0 43568 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_381
timestamp 1698431365
transform 1 0 44016 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_397
timestamp 1698431365
transform 1 0 45808 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_407
timestamp 1698431365
transform 1 0 46928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_411
timestamp 1698431365
transform 1 0 47376 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_419
timestamp 1698431365
transform 1 0 48272 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_422
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_486
timestamp 1698431365
transform 1 0 55776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_556
timestamp 1698431365
transform 1 0 63616 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_562
timestamp 1698431365
transform 1 0 64288 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_626
timestamp 1698431365
transform 1 0 71456 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_632
timestamp 1698431365
transform 1 0 72128 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_648
timestamp 1698431365
transform 1 0 73920 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_656
timestamp 1698431365
transform 1 0 74816 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_6
timestamp 1698431365
transform 1 0 2016 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_22
timestamp 1698431365
transform 1 0 3808 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_30
timestamp 1698431365
transform 1 0 4704 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_101
timestamp 1698431365
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_241
timestamp 1698431365
transform 1 0 28336 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_279
timestamp 1698431365
transform 1 0 32592 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_295
timestamp 1698431365
transform 1 0 34384 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_303
timestamp 1698431365
transform 1 0 35280 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_381
timestamp 1698431365
transform 1 0 44016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_451
timestamp 1698431365
transform 1 0 51856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_521
timestamp 1698431365
transform 1 0 59696 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_527
timestamp 1698431365
transform 1 0 60368 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_591
timestamp 1698431365
transform 1 0 67536 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_597
timestamp 1698431365
transform 1 0 68208 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_661
timestamp 1698431365
transform 1 0 75376 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_667
timestamp 1698431365
transform 1 0 76048 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_683
timestamp 1698431365
transform 1 0 77840 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_6
timestamp 1698431365
transform 1 0 2016 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698431365
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_206
timestamp 1698431365
transform 1 0 24416 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_276
timestamp 1698431365
transform 1 0 32256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_314
timestamp 1698431365
transform 1 0 36512 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_330
timestamp 1698431365
transform 1 0 38304 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_338
timestamp 1698431365
transform 1 0 39200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_368
timestamp 1698431365
transform 1 0 42560 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_372
timestamp 1698431365
transform 1 0 43008 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_381
timestamp 1698431365
transform 1 0 44016 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_385
timestamp 1698431365
transform 1 0 44464 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_417
timestamp 1698431365
transform 1 0 48048 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_419
timestamp 1698431365
transform 1 0 48272 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_486
timestamp 1698431365
transform 1 0 55776 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_556
timestamp 1698431365
transform 1 0 63616 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_562
timestamp 1698431365
transform 1 0 64288 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_626
timestamp 1698431365
transform 1 0 71456 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_632
timestamp 1698431365
transform 1 0 72128 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_664
timestamp 1698431365
transform 1 0 75712 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_680
timestamp 1698431365
transform 1 0 77504 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_6
timestamp 1698431365
transform 1 0 2016 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_22
timestamp 1698431365
transform 1 0 3808 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_30
timestamp 1698431365
transform 1 0 4704 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_171
timestamp 1698431365
transform 1 0 20496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_241
timestamp 1698431365
transform 1 0 28336 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_311
timestamp 1698431365
transform 1 0 36176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_381
timestamp 1698431365
transform 1 0 44016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_451
timestamp 1698431365
transform 1 0 51856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_521
timestamp 1698431365
transform 1 0 59696 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_527
timestamp 1698431365
transform 1 0 60368 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_591
timestamp 1698431365
transform 1 0 67536 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_597
timestamp 1698431365
transform 1 0 68208 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_661
timestamp 1698431365
transform 1 0 75376 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_667
timestamp 1698431365
transform 1 0 76048 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_683
timestamp 1698431365
transform 1 0 77840 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_6
timestamp 1698431365
transform 1 0 2016 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_276
timestamp 1698431365
transform 1 0 32256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_346
timestamp 1698431365
transform 1 0 40096 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_416
timestamp 1698431365
transform 1 0 47936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_422
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_486
timestamp 1698431365
transform 1 0 55776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_556
timestamp 1698431365
transform 1 0 63616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_562
timestamp 1698431365
transform 1 0 64288 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_626
timestamp 1698431365
transform 1 0 71456 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_632
timestamp 1698431365
transform 1 0 72128 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_664
timestamp 1698431365
transform 1 0 75712 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_680
timestamp 1698431365
transform 1 0 77504 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_10
timestamp 1698431365
transform 1 0 2464 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_26
timestamp 1698431365
transform 1 0 4256 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_171
timestamp 1698431365
transform 1 0 20496 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_241
timestamp 1698431365
transform 1 0 28336 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_311
timestamp 1698431365
transform 1 0 36176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_381
timestamp 1698431365
transform 1 0 44016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_451
timestamp 1698431365
transform 1 0 51856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_521
timestamp 1698431365
transform 1 0 59696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_527
timestamp 1698431365
transform 1 0 60368 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_591
timestamp 1698431365
transform 1 0 67536 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_597
timestamp 1698431365
transform 1 0 68208 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_661
timestamp 1698431365
transform 1 0 75376 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_667
timestamp 1698431365
transform 1 0 76048 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_675
timestamp 1698431365
transform 1 0 76944 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_679
timestamp 1698431365
transform 1 0 77392 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_6
timestamp 1698431365
transform 1 0 2016 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_136
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698431365
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_276
timestamp 1698431365
transform 1 0 32256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_346
timestamp 1698431365
transform 1 0 40096 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_416
timestamp 1698431365
transform 1 0 47936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_422
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_486
timestamp 1698431365
transform 1 0 55776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_556
timestamp 1698431365
transform 1 0 63616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_562
timestamp 1698431365
transform 1 0 64288 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_626
timestamp 1698431365
transform 1 0 71456 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_632
timestamp 1698431365
transform 1 0 72128 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_664
timestamp 1698431365
transform 1 0 75712 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_6
timestamp 1698431365
transform 1 0 2016 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_22
timestamp 1698431365
transform 1 0 3808 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_30
timestamp 1698431365
transform 1 0 4704 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_171
timestamp 1698431365
transform 1 0 20496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_241
timestamp 1698431365
transform 1 0 28336 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_311
timestamp 1698431365
transform 1 0 36176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_381
timestamp 1698431365
transform 1 0 44016 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_451
timestamp 1698431365
transform 1 0 51856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_521
timestamp 1698431365
transform 1 0 59696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_527
timestamp 1698431365
transform 1 0 60368 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_591
timestamp 1698431365
transform 1 0 67536 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_597
timestamp 1698431365
transform 1 0 68208 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_661
timestamp 1698431365
transform 1 0 75376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_667
timestamp 1698431365
transform 1 0 76048 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_683
timestamp 1698431365
transform 1 0 77840 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_6
timestamp 1698431365
transform 1 0 2016 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_136
timestamp 1698431365
transform 1 0 16576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_276
timestamp 1698431365
transform 1 0 32256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_346
timestamp 1698431365
transform 1 0 40096 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_416
timestamp 1698431365
transform 1 0 47936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_486
timestamp 1698431365
transform 1 0 55776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_556
timestamp 1698431365
transform 1 0 63616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_562
timestamp 1698431365
transform 1 0 64288 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_626
timestamp 1698431365
transform 1 0 71456 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_632
timestamp 1698431365
transform 1 0 72128 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_664
timestamp 1698431365
transform 1 0 75712 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_680
timestamp 1698431365
transform 1 0 77504 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_8
timestamp 1698431365
transform 1 0 2240 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_12
timestamp 1698431365
transform 1 0 2688 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_28
timestamp 1698431365
transform 1 0 4480 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_32
timestamp 1698431365
transform 1 0 4928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_171
timestamp 1698431365
transform 1 0 20496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_241
timestamp 1698431365
transform 1 0 28336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698431365
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_381
timestamp 1698431365
transform 1 0 44016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698431365
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_521
timestamp 1698431365
transform 1 0 59696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_527
timestamp 1698431365
transform 1 0 60368 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_591
timestamp 1698431365
transform 1 0 67536 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_597
timestamp 1698431365
transform 1 0 68208 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_661
timestamp 1698431365
transform 1 0 75376 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_667
timestamp 1698431365
transform 1 0 76048 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_683
timestamp 1698431365
transform 1 0 77840 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_6
timestamp 1698431365
transform 1 0 2016 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698431365
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_206
timestamp 1698431365
transform 1 0 24416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_276
timestamp 1698431365
transform 1 0 32256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_346
timestamp 1698431365
transform 1 0 40096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_416
timestamp 1698431365
transform 1 0 47936 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_556
timestamp 1698431365
transform 1 0 63616 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_562
timestamp 1698431365
transform 1 0 64288 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_626
timestamp 1698431365
transform 1 0 71456 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_632
timestamp 1698431365
transform 1 0 72128 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_648
timestamp 1698431365
transform 1 0 73920 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_656
timestamp 1698431365
transform 1 0 74816 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_10
timestamp 1698431365
transform 1 0 2464 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_26
timestamp 1698431365
transform 1 0 4256 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_171
timestamp 1698431365
transform 1 0 20496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_241
timestamp 1698431365
transform 1 0 28336 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_311
timestamp 1698431365
transform 1 0 36176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_381
timestamp 1698431365
transform 1 0 44016 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_451
timestamp 1698431365
transform 1 0 51856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_521
timestamp 1698431365
transform 1 0 59696 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_527
timestamp 1698431365
transform 1 0 60368 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_591
timestamp 1698431365
transform 1 0 67536 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_597
timestamp 1698431365
transform 1 0 68208 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_661
timestamp 1698431365
transform 1 0 75376 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_667
timestamp 1698431365
transform 1 0 76048 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_675
timestamp 1698431365
transform 1 0 76944 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_679
timestamp 1698431365
transform 1 0 77392 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_6
timestamp 1698431365
transform 1 0 2016 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_136
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_142
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_206
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_212
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_276
timestamp 1698431365
transform 1 0 32256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_282
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_346
timestamp 1698431365
transform 1 0 40096 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_416
timestamp 1698431365
transform 1 0 47936 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_422
timestamp 1698431365
transform 1 0 48608 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_486
timestamp 1698431365
transform 1 0 55776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_492
timestamp 1698431365
transform 1 0 56448 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_556
timestamp 1698431365
transform 1 0 63616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_562
timestamp 1698431365
transform 1 0 64288 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_626
timestamp 1698431365
transform 1 0 71456 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_632
timestamp 1698431365
transform 1 0 72128 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_664
timestamp 1698431365
transform 1 0 75712 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_680
timestamp 1698431365
transform 1 0 77504 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_6
timestamp 1698431365
transform 1 0 2016 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_22
timestamp 1698431365
transform 1 0 3808 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_30
timestamp 1698431365
transform 1 0 4704 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1698431365
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_37
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_101
timestamp 1698431365
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_107
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_171
timestamp 1698431365
transform 1 0 20496 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_177
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_241
timestamp 1698431365
transform 1 0 28336 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_247
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_311
timestamp 1698431365
transform 1 0 36176 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_317
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_381
timestamp 1698431365
transform 1 0 44016 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_387
timestamp 1698431365
transform 1 0 44688 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_451
timestamp 1698431365
transform 1 0 51856 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_457
timestamp 1698431365
transform 1 0 52528 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_521
timestamp 1698431365
transform 1 0 59696 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_527
timestamp 1698431365
transform 1 0 60368 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_591
timestamp 1698431365
transform 1 0 67536 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_597
timestamp 1698431365
transform 1 0 68208 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_661
timestamp 1698431365
transform 1 0 75376 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_667
timestamp 1698431365
transform 1 0 76048 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_675
timestamp 1698431365
transform 1 0 76944 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_679
timestamp 1698431365
transform 1 0 77392 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_6
timestamp 1698431365
transform 1 0 2016 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_72
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_136
timestamp 1698431365
transform 1 0 16576 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_206
timestamp 1698431365
transform 1 0 24416 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_212
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_276
timestamp 1698431365
transform 1 0 32256 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_346
timestamp 1698431365
transform 1 0 40096 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_352
timestamp 1698431365
transform 1 0 40768 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_416
timestamp 1698431365
transform 1 0 47936 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_422
timestamp 1698431365
transform 1 0 48608 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_486
timestamp 1698431365
transform 1 0 55776 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_492
timestamp 1698431365
transform 1 0 56448 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_556
timestamp 1698431365
transform 1 0 63616 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_562
timestamp 1698431365
transform 1 0 64288 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_626
timestamp 1698431365
transform 1 0 71456 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_632
timestamp 1698431365
transform 1 0 72128 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_648
timestamp 1698431365
transform 1 0 73920 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_656
timestamp 1698431365
transform 1 0 74816 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_6
timestamp 1698431365
transform 1 0 2016 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_22
timestamp 1698431365
transform 1 0 3808 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_30
timestamp 1698431365
transform 1 0 4704 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698431365
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_101
timestamp 1698431365
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_107
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_171
timestamp 1698431365
transform 1 0 20496 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_241
timestamp 1698431365
transform 1 0 28336 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_311
timestamp 1698431365
transform 1 0 36176 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_381
timestamp 1698431365
transform 1 0 44016 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_387
timestamp 1698431365
transform 1 0 44688 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_451
timestamp 1698431365
transform 1 0 51856 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_457
timestamp 1698431365
transform 1 0 52528 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_521
timestamp 1698431365
transform 1 0 59696 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_527
timestamp 1698431365
transform 1 0 60368 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_591
timestamp 1698431365
transform 1 0 67536 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_597
timestamp 1698431365
transform 1 0 68208 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_661
timestamp 1698431365
transform 1 0 75376 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_667
timestamp 1698431365
transform 1 0 76048 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_683
timestamp 1698431365
transform 1 0 77840 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_6
timestamp 1698431365
transform 1 0 2016 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_72
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_136
timestamp 1698431365
transform 1 0 16576 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_142
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_206
timestamp 1698431365
transform 1 0 24416 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_276
timestamp 1698431365
transform 1 0 32256 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_282
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_346
timestamp 1698431365
transform 1 0 40096 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_352
timestamp 1698431365
transform 1 0 40768 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_416
timestamp 1698431365
transform 1 0 47936 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_422
timestamp 1698431365
transform 1 0 48608 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_486
timestamp 1698431365
transform 1 0 55776 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_492
timestamp 1698431365
transform 1 0 56448 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_556
timestamp 1698431365
transform 1 0 63616 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_562
timestamp 1698431365
transform 1 0 64288 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_626
timestamp 1698431365
transform 1 0 71456 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_632
timestamp 1698431365
transform 1 0 72128 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_664
timestamp 1698431365
transform 1 0 75712 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_10
timestamp 1698431365
transform 1 0 2464 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_26
timestamp 1698431365
transform 1 0 4256 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_37
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_101
timestamp 1698431365
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_107
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_171
timestamp 1698431365
transform 1 0 20496 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_241
timestamp 1698431365
transform 1 0 28336 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_247
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_311
timestamp 1698431365
transform 1 0 36176 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_317
timestamp 1698431365
transform 1 0 36848 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_381
timestamp 1698431365
transform 1 0 44016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_387
timestamp 1698431365
transform 1 0 44688 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_451
timestamp 1698431365
transform 1 0 51856 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_457
timestamp 1698431365
transform 1 0 52528 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_521
timestamp 1698431365
transform 1 0 59696 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_527
timestamp 1698431365
transform 1 0 60368 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_591
timestamp 1698431365
transform 1 0 67536 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_597
timestamp 1698431365
transform 1 0 68208 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_661
timestamp 1698431365
transform 1 0 75376 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_667
timestamp 1698431365
transform 1 0 76048 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_683
timestamp 1698431365
transform 1 0 77840 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_687
timestamp 1698431365
transform 1 0 78288 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_8
timestamp 1698431365
transform 1 0 2240 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_12
timestamp 1698431365
transform 1 0 2688 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_44
timestamp 1698431365
transform 1 0 6272 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_60
timestamp 1698431365
transform 1 0 8064 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_68
timestamp 1698431365
transform 1 0 8960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_72
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_136
timestamp 1698431365
transform 1 0 16576 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_142
timestamp 1698431365
transform 1 0 17248 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_206
timestamp 1698431365
transform 1 0 24416 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_212
timestamp 1698431365
transform 1 0 25088 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_276
timestamp 1698431365
transform 1 0 32256 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_282
timestamp 1698431365
transform 1 0 32928 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_346
timestamp 1698431365
transform 1 0 40096 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_352
timestamp 1698431365
transform 1 0 40768 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_416
timestamp 1698431365
transform 1 0 47936 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_422
timestamp 1698431365
transform 1 0 48608 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_486
timestamp 1698431365
transform 1 0 55776 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_492
timestamp 1698431365
transform 1 0 56448 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_556
timestamp 1698431365
transform 1 0 63616 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_562
timestamp 1698431365
transform 1 0 64288 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_626
timestamp 1698431365
transform 1 0 71456 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_632
timestamp 1698431365
transform 1 0 72128 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_664
timestamp 1698431365
transform 1 0 75712 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_680
timestamp 1698431365
transform 1 0 77504 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_6
timestamp 1698431365
transform 1 0 2016 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_22
timestamp 1698431365
transform 1 0 3808 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_30
timestamp 1698431365
transform 1 0 4704 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_34
timestamp 1698431365
transform 1 0 5152 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_37
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_101
timestamp 1698431365
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_107
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_171
timestamp 1698431365
transform 1 0 20496 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_177
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_241
timestamp 1698431365
transform 1 0 28336 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_247
timestamp 1698431365
transform 1 0 29008 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_311
timestamp 1698431365
transform 1 0 36176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_317
timestamp 1698431365
transform 1 0 36848 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_381
timestamp 1698431365
transform 1 0 44016 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_387
timestamp 1698431365
transform 1 0 44688 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_451
timestamp 1698431365
transform 1 0 51856 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_457
timestamp 1698431365
transform 1 0 52528 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_521
timestamp 1698431365
transform 1 0 59696 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_527
timestamp 1698431365
transform 1 0 60368 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_591
timestamp 1698431365
transform 1 0 67536 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_597
timestamp 1698431365
transform 1 0 68208 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_661
timestamp 1698431365
transform 1 0 75376 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_667
timestamp 1698431365
transform 1 0 76048 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_683
timestamp 1698431365
transform 1 0 77840 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_687
timestamp 1698431365
transform 1 0 78288 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_6
timestamp 1698431365
transform 1 0 2016 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_72
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_136
timestamp 1698431365
transform 1 0 16576 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_142
timestamp 1698431365
transform 1 0 17248 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_206
timestamp 1698431365
transform 1 0 24416 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_212
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_276
timestamp 1698431365
transform 1 0 32256 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_282
timestamp 1698431365
transform 1 0 32928 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_346
timestamp 1698431365
transform 1 0 40096 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_352
timestamp 1698431365
transform 1 0 40768 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_416
timestamp 1698431365
transform 1 0 47936 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_422
timestamp 1698431365
transform 1 0 48608 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_486
timestamp 1698431365
transform 1 0 55776 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_492
timestamp 1698431365
transform 1 0 56448 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_556
timestamp 1698431365
transform 1 0 63616 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_562
timestamp 1698431365
transform 1 0 64288 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_626
timestamp 1698431365
transform 1 0 71456 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_632
timestamp 1698431365
transform 1 0 72128 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_664
timestamp 1698431365
transform 1 0 75712 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_680
timestamp 1698431365
transform 1 0 77504 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_6
timestamp 1698431365
transform 1 0 2016 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_22
timestamp 1698431365
transform 1 0 3808 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_30
timestamp 1698431365
transform 1 0 4704 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1698431365
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_101
timestamp 1698431365
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_107
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_171
timestamp 1698431365
transform 1 0 20496 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_241
timestamp 1698431365
transform 1 0 28336 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_247
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_311
timestamp 1698431365
transform 1 0 36176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_317
timestamp 1698431365
transform 1 0 36848 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_381
timestamp 1698431365
transform 1 0 44016 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_387
timestamp 1698431365
transform 1 0 44688 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_451
timestamp 1698431365
transform 1 0 51856 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_457
timestamp 1698431365
transform 1 0 52528 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_521
timestamp 1698431365
transform 1 0 59696 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_527
timestamp 1698431365
transform 1 0 60368 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_591
timestamp 1698431365
transform 1 0 67536 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_597
timestamp 1698431365
transform 1 0 68208 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_661
timestamp 1698431365
transform 1 0 75376 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_667
timestamp 1698431365
transform 1 0 76048 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_683
timestamp 1698431365
transform 1 0 77840 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_687
timestamp 1698431365
transform 1 0 78288 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_6
timestamp 1698431365
transform 1 0 2016 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_72
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_136
timestamp 1698431365
transform 1 0 16576 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_142
timestamp 1698431365
transform 1 0 17248 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_206
timestamp 1698431365
transform 1 0 24416 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_212
timestamp 1698431365
transform 1 0 25088 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_276
timestamp 1698431365
transform 1 0 32256 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_282
timestamp 1698431365
transform 1 0 32928 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_346
timestamp 1698431365
transform 1 0 40096 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_352
timestamp 1698431365
transform 1 0 40768 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_416
timestamp 1698431365
transform 1 0 47936 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_422
timestamp 1698431365
transform 1 0 48608 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_486
timestamp 1698431365
transform 1 0 55776 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_492
timestamp 1698431365
transform 1 0 56448 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_556
timestamp 1698431365
transform 1 0 63616 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_562
timestamp 1698431365
transform 1 0 64288 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_626
timestamp 1698431365
transform 1 0 71456 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_632
timestamp 1698431365
transform 1 0 72128 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_664
timestamp 1698431365
transform 1 0 75712 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_680
timestamp 1698431365
transform 1 0 77504 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_12
timestamp 1698431365
transform 1 0 2688 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_16
timestamp 1698431365
transform 1 0 3136 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_32
timestamp 1698431365
transform 1 0 4928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698431365
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_37
timestamp 1698431365
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_101
timestamp 1698431365
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_107
timestamp 1698431365
transform 1 0 13328 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_171
timestamp 1698431365
transform 1 0 20496 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_177
timestamp 1698431365
transform 1 0 21168 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_241
timestamp 1698431365
transform 1 0 28336 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_247
timestamp 1698431365
transform 1 0 29008 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_311
timestamp 1698431365
transform 1 0 36176 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_317
timestamp 1698431365
transform 1 0 36848 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_381
timestamp 1698431365
transform 1 0 44016 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_387
timestamp 1698431365
transform 1 0 44688 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_451
timestamp 1698431365
transform 1 0 51856 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_457
timestamp 1698431365
transform 1 0 52528 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_521
timestamp 1698431365
transform 1 0 59696 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_527
timestamp 1698431365
transform 1 0 60368 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_591
timestamp 1698431365
transform 1 0 67536 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_597
timestamp 1698431365
transform 1 0 68208 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_661
timestamp 1698431365
transform 1 0 75376 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_667
timestamp 1698431365
transform 1 0 76048 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_683
timestamp 1698431365
transform 1 0 77840 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_687
timestamp 1698431365
transform 1 0 78288 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_6
timestamp 1698431365
transform 1 0 2016 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_72
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_136
timestamp 1698431365
transform 1 0 16576 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_142
timestamp 1698431365
transform 1 0 17248 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_206
timestamp 1698431365
transform 1 0 24416 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_212
timestamp 1698431365
transform 1 0 25088 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_276
timestamp 1698431365
transform 1 0 32256 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_282
timestamp 1698431365
transform 1 0 32928 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_346
timestamp 1698431365
transform 1 0 40096 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_352
timestamp 1698431365
transform 1 0 40768 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_416
timestamp 1698431365
transform 1 0 47936 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_422
timestamp 1698431365
transform 1 0 48608 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_486
timestamp 1698431365
transform 1 0 55776 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_492
timestamp 1698431365
transform 1 0 56448 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_556
timestamp 1698431365
transform 1 0 63616 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_562
timestamp 1698431365
transform 1 0 64288 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_626
timestamp 1698431365
transform 1 0 71456 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_632
timestamp 1698431365
transform 1 0 72128 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_664
timestamp 1698431365
transform 1 0 75712 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_680
timestamp 1698431365
transform 1 0 77504 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_6
timestamp 1698431365
transform 1 0 2016 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_22
timestamp 1698431365
transform 1 0 3808 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_30
timestamp 1698431365
transform 1 0 4704 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_34
timestamp 1698431365
transform 1 0 5152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_37
timestamp 1698431365
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_101
timestamp 1698431365
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_107
timestamp 1698431365
transform 1 0 13328 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_171
timestamp 1698431365
transform 1 0 20496 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_177
timestamp 1698431365
transform 1 0 21168 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_241
timestamp 1698431365
transform 1 0 28336 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_247
timestamp 1698431365
transform 1 0 29008 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_311
timestamp 1698431365
transform 1 0 36176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_317
timestamp 1698431365
transform 1 0 36848 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_381
timestamp 1698431365
transform 1 0 44016 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_387
timestamp 1698431365
transform 1 0 44688 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_451
timestamp 1698431365
transform 1 0 51856 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_457
timestamp 1698431365
transform 1 0 52528 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_521
timestamp 1698431365
transform 1 0 59696 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_527
timestamp 1698431365
transform 1 0 60368 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_591
timestamp 1698431365
transform 1 0 67536 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_597
timestamp 1698431365
transform 1 0 68208 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_661
timestamp 1698431365
transform 1 0 75376 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_667
timestamp 1698431365
transform 1 0 76048 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_683
timestamp 1698431365
transform 1 0 77840 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_687
timestamp 1698431365
transform 1 0 78288 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_6
timestamp 1698431365
transform 1 0 2016 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_72
timestamp 1698431365
transform 1 0 9408 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_136
timestamp 1698431365
transform 1 0 16576 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_142
timestamp 1698431365
transform 1 0 17248 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_206
timestamp 1698431365
transform 1 0 24416 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_212
timestamp 1698431365
transform 1 0 25088 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_276
timestamp 1698431365
transform 1 0 32256 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_282
timestamp 1698431365
transform 1 0 32928 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_346
timestamp 1698431365
transform 1 0 40096 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_352
timestamp 1698431365
transform 1 0 40768 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_416
timestamp 1698431365
transform 1 0 47936 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_422
timestamp 1698431365
transform 1 0 48608 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_486
timestamp 1698431365
transform 1 0 55776 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_492
timestamp 1698431365
transform 1 0 56448 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_556
timestamp 1698431365
transform 1 0 63616 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_562
timestamp 1698431365
transform 1 0 64288 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_626
timestamp 1698431365
transform 1 0 71456 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_632
timestamp 1698431365
transform 1 0 72128 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_664
timestamp 1698431365
transform 1 0 75712 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_680
timestamp 1698431365
transform 1 0 77504 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_28
timestamp 1698431365
transform 1 0 4480 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_32
timestamp 1698431365
transform 1 0 4928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_34
timestamp 1698431365
transform 1 0 5152 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_37
timestamp 1698431365
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_101
timestamp 1698431365
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_107
timestamp 1698431365
transform 1 0 13328 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_171
timestamp 1698431365
transform 1 0 20496 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_177
timestamp 1698431365
transform 1 0 21168 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_241
timestamp 1698431365
transform 1 0 28336 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_247
timestamp 1698431365
transform 1 0 29008 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_311
timestamp 1698431365
transform 1 0 36176 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_317
timestamp 1698431365
transform 1 0 36848 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_381
timestamp 1698431365
transform 1 0 44016 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_387
timestamp 1698431365
transform 1 0 44688 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_451
timestamp 1698431365
transform 1 0 51856 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_457
timestamp 1698431365
transform 1 0 52528 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_521
timestamp 1698431365
transform 1 0 59696 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_527
timestamp 1698431365
transform 1 0 60368 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_591
timestamp 1698431365
transform 1 0 67536 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_597
timestamp 1698431365
transform 1 0 68208 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_661
timestamp 1698431365
transform 1 0 75376 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_667
timestamp 1698431365
transform 1 0 76048 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_683
timestamp 1698431365
transform 1 0 77840 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_687
timestamp 1698431365
transform 1 0 78288 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_2
timestamp 1698431365
transform 1 0 1568 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_66
timestamp 1698431365
transform 1 0 8736 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_72
timestamp 1698431365
transform 1 0 9408 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_136
timestamp 1698431365
transform 1 0 16576 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_142
timestamp 1698431365
transform 1 0 17248 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_206
timestamp 1698431365
transform 1 0 24416 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_212
timestamp 1698431365
transform 1 0 25088 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_276
timestamp 1698431365
transform 1 0 32256 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_282
timestamp 1698431365
transform 1 0 32928 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_346
timestamp 1698431365
transform 1 0 40096 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_352
timestamp 1698431365
transform 1 0 40768 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_416
timestamp 1698431365
transform 1 0 47936 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_422
timestamp 1698431365
transform 1 0 48608 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_486
timestamp 1698431365
transform 1 0 55776 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_492
timestamp 1698431365
transform 1 0 56448 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_556
timestamp 1698431365
transform 1 0 63616 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_562
timestamp 1698431365
transform 1 0 64288 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_626
timestamp 1698431365
transform 1 0 71456 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_632
timestamp 1698431365
transform 1 0 72128 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_664
timestamp 1698431365
transform 1 0 75712 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_680
timestamp 1698431365
transform 1 0 77504 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_2
timestamp 1698431365
transform 1 0 1568 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_34
timestamp 1698431365
transform 1 0 5152 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_37
timestamp 1698431365
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_101
timestamp 1698431365
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_107
timestamp 1698431365
transform 1 0 13328 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_171
timestamp 1698431365
transform 1 0 20496 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_177
timestamp 1698431365
transform 1 0 21168 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_241
timestamp 1698431365
transform 1 0 28336 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_247
timestamp 1698431365
transform 1 0 29008 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_311
timestamp 1698431365
transform 1 0 36176 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_317
timestamp 1698431365
transform 1 0 36848 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_381
timestamp 1698431365
transform 1 0 44016 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_387
timestamp 1698431365
transform 1 0 44688 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_451
timestamp 1698431365
transform 1 0 51856 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_457
timestamp 1698431365
transform 1 0 52528 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_521
timestamp 1698431365
transform 1 0 59696 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_527
timestamp 1698431365
transform 1 0 60368 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_591
timestamp 1698431365
transform 1 0 67536 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_597
timestamp 1698431365
transform 1 0 68208 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_661
timestamp 1698431365
transform 1 0 75376 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_667
timestamp 1698431365
transform 1 0 76048 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_683
timestamp 1698431365
transform 1 0 77840 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_687
timestamp 1698431365
transform 1 0 78288 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_2
timestamp 1698431365
transform 1 0 1568 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_66
timestamp 1698431365
transform 1 0 8736 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_72
timestamp 1698431365
transform 1 0 9408 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_136
timestamp 1698431365
transform 1 0 16576 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_142
timestamp 1698431365
transform 1 0 17248 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_206
timestamp 1698431365
transform 1 0 24416 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_212
timestamp 1698431365
transform 1 0 25088 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_276
timestamp 1698431365
transform 1 0 32256 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_282
timestamp 1698431365
transform 1 0 32928 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_346
timestamp 1698431365
transform 1 0 40096 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_352
timestamp 1698431365
transform 1 0 40768 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_416
timestamp 1698431365
transform 1 0 47936 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_422
timestamp 1698431365
transform 1 0 48608 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_486
timestamp 1698431365
transform 1 0 55776 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_492
timestamp 1698431365
transform 1 0 56448 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_556
timestamp 1698431365
transform 1 0 63616 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_562
timestamp 1698431365
transform 1 0 64288 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_626
timestamp 1698431365
transform 1 0 71456 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_632
timestamp 1698431365
transform 1 0 72128 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_664
timestamp 1698431365
transform 1 0 75712 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_680
timestamp 1698431365
transform 1 0 77504 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_2
timestamp 1698431365
transform 1 0 1568 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_34
timestamp 1698431365
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_37
timestamp 1698431365
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_101
timestamp 1698431365
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_107
timestamp 1698431365
transform 1 0 13328 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_171
timestamp 1698431365
transform 1 0 20496 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_177
timestamp 1698431365
transform 1 0 21168 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_241
timestamp 1698431365
transform 1 0 28336 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_247
timestamp 1698431365
transform 1 0 29008 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_311
timestamp 1698431365
transform 1 0 36176 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_317
timestamp 1698431365
transform 1 0 36848 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_381
timestamp 1698431365
transform 1 0 44016 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_387
timestamp 1698431365
transform 1 0 44688 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_451
timestamp 1698431365
transform 1 0 51856 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_457
timestamp 1698431365
transform 1 0 52528 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_521
timestamp 1698431365
transform 1 0 59696 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_527
timestamp 1698431365
transform 1 0 60368 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_591
timestamp 1698431365
transform 1 0 67536 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_597
timestamp 1698431365
transform 1 0 68208 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_661
timestamp 1698431365
transform 1 0 75376 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_667
timestamp 1698431365
transform 1 0 76048 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_683
timestamp 1698431365
transform 1 0 77840 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_687
timestamp 1698431365
transform 1 0 78288 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_2
timestamp 1698431365
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_66
timestamp 1698431365
transform 1 0 8736 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_72
timestamp 1698431365
transform 1 0 9408 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_136
timestamp 1698431365
transform 1 0 16576 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_142
timestamp 1698431365
transform 1 0 17248 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_206
timestamp 1698431365
transform 1 0 24416 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_212
timestamp 1698431365
transform 1 0 25088 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_276
timestamp 1698431365
transform 1 0 32256 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_282
timestamp 1698431365
transform 1 0 32928 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_346
timestamp 1698431365
transform 1 0 40096 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_352
timestamp 1698431365
transform 1 0 40768 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_416
timestamp 1698431365
transform 1 0 47936 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_422
timestamp 1698431365
transform 1 0 48608 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_486
timestamp 1698431365
transform 1 0 55776 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_492
timestamp 1698431365
transform 1 0 56448 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_556
timestamp 1698431365
transform 1 0 63616 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_562
timestamp 1698431365
transform 1 0 64288 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_626
timestamp 1698431365
transform 1 0 71456 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_632
timestamp 1698431365
transform 1 0 72128 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_664
timestamp 1698431365
transform 1 0 75712 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_87_680
timestamp 1698431365
transform 1 0 77504 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_2
timestamp 1698431365
transform 1 0 1568 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_34
timestamp 1698431365
transform 1 0 5152 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_37
timestamp 1698431365
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_101
timestamp 1698431365
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_107
timestamp 1698431365
transform 1 0 13328 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_171
timestamp 1698431365
transform 1 0 20496 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_177
timestamp 1698431365
transform 1 0 21168 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_241
timestamp 1698431365
transform 1 0 28336 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_247
timestamp 1698431365
transform 1 0 29008 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_311
timestamp 1698431365
transform 1 0 36176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_317
timestamp 1698431365
transform 1 0 36848 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_381
timestamp 1698431365
transform 1 0 44016 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_387
timestamp 1698431365
transform 1 0 44688 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_451
timestamp 1698431365
transform 1 0 51856 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_457
timestamp 1698431365
transform 1 0 52528 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_521
timestamp 1698431365
transform 1 0 59696 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_527
timestamp 1698431365
transform 1 0 60368 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_591
timestamp 1698431365
transform 1 0 67536 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_597
timestamp 1698431365
transform 1 0 68208 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_661
timestamp 1698431365
transform 1 0 75376 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_667
timestamp 1698431365
transform 1 0 76048 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_683
timestamp 1698431365
transform 1 0 77840 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_687
timestamp 1698431365
transform 1 0 78288 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_2
timestamp 1698431365
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_66
timestamp 1698431365
transform 1 0 8736 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_72
timestamp 1698431365
transform 1 0 9408 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_136
timestamp 1698431365
transform 1 0 16576 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_142
timestamp 1698431365
transform 1 0 17248 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_206
timestamp 1698431365
transform 1 0 24416 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_212
timestamp 1698431365
transform 1 0 25088 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_276
timestamp 1698431365
transform 1 0 32256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_282
timestamp 1698431365
transform 1 0 32928 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_346
timestamp 1698431365
transform 1 0 40096 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_352
timestamp 1698431365
transform 1 0 40768 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_416
timestamp 1698431365
transform 1 0 47936 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_422
timestamp 1698431365
transform 1 0 48608 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_486
timestamp 1698431365
transform 1 0 55776 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_492
timestamp 1698431365
transform 1 0 56448 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_556
timestamp 1698431365
transform 1 0 63616 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_562
timestamp 1698431365
transform 1 0 64288 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_626
timestamp 1698431365
transform 1 0 71456 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_632
timestamp 1698431365
transform 1 0 72128 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_664
timestamp 1698431365
transform 1 0 75712 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_680
timestamp 1698431365
transform 1 0 77504 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_2
timestamp 1698431365
transform 1 0 1568 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_34
timestamp 1698431365
transform 1 0 5152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_37
timestamp 1698431365
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_101
timestamp 1698431365
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_107
timestamp 1698431365
transform 1 0 13328 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_171
timestamp 1698431365
transform 1 0 20496 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_177
timestamp 1698431365
transform 1 0 21168 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_241
timestamp 1698431365
transform 1 0 28336 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_247
timestamp 1698431365
transform 1 0 29008 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_311
timestamp 1698431365
transform 1 0 36176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_317
timestamp 1698431365
transform 1 0 36848 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_381
timestamp 1698431365
transform 1 0 44016 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_387
timestamp 1698431365
transform 1 0 44688 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_451
timestamp 1698431365
transform 1 0 51856 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_457
timestamp 1698431365
transform 1 0 52528 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_521
timestamp 1698431365
transform 1 0 59696 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_527
timestamp 1698431365
transform 1 0 60368 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_591
timestamp 1698431365
transform 1 0 67536 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_597
timestamp 1698431365
transform 1 0 68208 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_661
timestamp 1698431365
transform 1 0 75376 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_667
timestamp 1698431365
transform 1 0 76048 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_683
timestamp 1698431365
transform 1 0 77840 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_687
timestamp 1698431365
transform 1 0 78288 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_2
timestamp 1698431365
transform 1 0 1568 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_66
timestamp 1698431365
transform 1 0 8736 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_72
timestamp 1698431365
transform 1 0 9408 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_136
timestamp 1698431365
transform 1 0 16576 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_142
timestamp 1698431365
transform 1 0 17248 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_206
timestamp 1698431365
transform 1 0 24416 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_212
timestamp 1698431365
transform 1 0 25088 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_276
timestamp 1698431365
transform 1 0 32256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_282
timestamp 1698431365
transform 1 0 32928 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_314
timestamp 1698431365
transform 1 0 36512 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_317
timestamp 1698431365
transform 1 0 36848 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_333
timestamp 1698431365
transform 1 0 38640 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_341
timestamp 1698431365
transform 1 0 39536 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_345
timestamp 1698431365
transform 1 0 39984 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_349
timestamp 1698431365
transform 1 0 40432 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_352
timestamp 1698431365
transform 1 0 40768 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_356
timestamp 1698431365
transform 1 0 41216 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_360
timestamp 1698431365
transform 1 0 41664 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_365
timestamp 1698431365
transform 1 0 42224 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_373
timestamp 1698431365
transform 1 0 43120 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_376
timestamp 1698431365
transform 1 0 43456 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_408
timestamp 1698431365
transform 1 0 47040 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_416
timestamp 1698431365
transform 1 0 47936 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_422
timestamp 1698431365
transform 1 0 48608 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_438
timestamp 1698431365
transform 1 0 50400 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_442
timestamp 1698431365
transform 1 0 50848 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_471
timestamp 1698431365
transform 1 0 54096 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_475
timestamp 1698431365
transform 1 0 54544 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_483
timestamp 1698431365
transform 1 0 55440 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_487
timestamp 1698431365
transform 1 0 55888 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_489
timestamp 1698431365
transform 1 0 56112 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_492
timestamp 1698431365
transform 1 0 56448 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_556
timestamp 1698431365
transform 1 0 63616 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_562
timestamp 1698431365
transform 1 0 64288 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_626
timestamp 1698431365
transform 1 0 71456 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_632
timestamp 1698431365
transform 1 0 72128 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_664
timestamp 1698431365
transform 1 0 75712 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_680
timestamp 1698431365
transform 1 0 77504 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_2
timestamp 1698431365
transform 1 0 1568 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_34
timestamp 1698431365
transform 1 0 5152 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_37
timestamp 1698431365
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_101
timestamp 1698431365
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_107
timestamp 1698431365
transform 1 0 13328 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_171
timestamp 1698431365
transform 1 0 20496 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_177
timestamp 1698431365
transform 1 0 21168 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_185
timestamp 1698431365
transform 1 0 22064 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_213
timestamp 1698431365
transform 1 0 25200 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_217
timestamp 1698431365
transform 1 0 25648 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_233
timestamp 1698431365
transform 1 0 27440 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_237
timestamp 1698431365
transform 1 0 27888 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_240
timestamp 1698431365
transform 1 0 28224 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_242
timestamp 1698431365
transform 1 0 28448 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_257
timestamp 1698431365
transform 1 0 30128 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_263
timestamp 1698431365
transform 1 0 30800 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_269
timestamp 1698431365
transform 1 0 31472 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_273
timestamp 1698431365
transform 1 0 31920 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_317
timestamp 1698431365
transform 1 0 36848 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_321
timestamp 1698431365
transform 1 0 37296 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_379
timestamp 1698431365
transform 1 0 43792 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_383
timestamp 1698431365
transform 1 0 44240 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_387
timestamp 1698431365
transform 1 0 44688 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_419
timestamp 1698431365
transform 1 0 48272 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_435
timestamp 1698431365
transform 1 0 50064 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_439
timestamp 1698431365
transform 1 0 50512 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_441
timestamp 1698431365
transform 1 0 50736 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_444
timestamp 1698431365
transform 1 0 51072 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_448
timestamp 1698431365
transform 1 0 51520 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_483
timestamp 1698431365
transform 1 0 55440 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_491
timestamp 1698431365
transform 1 0 56336 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_495
timestamp 1698431365
transform 1 0 56784 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_503
timestamp 1698431365
transform 1 0 57680 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_507
timestamp 1698431365
transform 1 0 58128 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_509
timestamp 1698431365
transform 1 0 58352 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_512
timestamp 1698431365
transform 1 0 58688 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_520
timestamp 1698431365
transform 1 0 59584 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_524
timestamp 1698431365
transform 1 0 60032 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_527
timestamp 1698431365
transform 1 0 60368 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_591
timestamp 1698431365
transform 1 0 67536 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_597
timestamp 1698431365
transform 1 0 68208 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_661
timestamp 1698431365
transform 1 0 75376 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_667
timestamp 1698431365
transform 1 0 76048 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_683
timestamp 1698431365
transform 1 0 77840 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_687
timestamp 1698431365
transform 1 0 78288 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_2
timestamp 1698431365
transform 1 0 1568 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_36
timestamp 1698431365
transform 1 0 5376 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_70
timestamp 1698431365
transform 1 0 9184 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_104
timestamp 1698431365
transform 1 0 12992 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_138
timestamp 1698431365
transform 1 0 16800 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_172
timestamp 1698431365
transform 1 0 20608 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_188
timestamp 1698431365
transform 1 0 22400 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_190
timestamp 1698431365
transform 1 0 22624 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_197
timestamp 1698431365
transform 1 0 23408 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_199
timestamp 1698431365
transform 1 0 23632 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_216
timestamp 1698431365
transform 1 0 25536 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_221
timestamp 1698431365
transform 1 0 26096 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_227
timestamp 1698431365
transform 1 0 26768 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_266
timestamp 1698431365
transform 1 0 31136 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_274
timestamp 1698431365
transform 1 0 32032 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_276
timestamp 1698431365
transform 1 0 32256 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_281
timestamp 1698431365
transform 1 0 32816 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_287
timestamp 1698431365
transform 1 0 33488 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_291
timestamp 1698431365
transform 1 0 33936 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_299
timestamp 1698431365
transform 1 0 34832 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_305
timestamp 1698431365
transform 1 0 35504 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_318
timestamp 1698431365
transform 1 0 36960 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_329
timestamp 1698431365
transform 1 0 38192 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_333
timestamp 1698431365
transform 1 0 38640 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_335
timestamp 1698431365
transform 1 0 38864 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_342
timestamp 1698431365
transform 1 0 39648 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_347
timestamp 1698431365
transform 1 0 40208 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_390
timestamp 1698431365
transform 1 0 45024 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_395
timestamp 1698431365
transform 1 0 45584 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_401
timestamp 1698431365
transform 1 0 46256 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_407
timestamp 1698431365
transform 1 0 46928 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_410
timestamp 1698431365
transform 1 0 47264 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_412
timestamp 1698431365
transform 1 0 47488 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_419
timestamp 1698431365
transform 1 0 48272 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_431
timestamp 1698431365
transform 1 0 49616 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_433
timestamp 1698431365
transform 1 0 49840 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_492
timestamp 1698431365
transform 1 0 56448 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_503
timestamp 1698431365
transform 1 0 57680 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_509
timestamp 1698431365
transform 1 0 58352 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_538
timestamp 1698431365
transform 1 0 61600 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_542
timestamp 1698431365
transform 1 0 62048 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_546
timestamp 1698431365
transform 1 0 62496 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_580
timestamp 1698431365
transform 1 0 66304 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_614
timestamp 1698431365
transform 1 0 70112 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_648
timestamp 1698431365
transform 1 0 73920 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_682
timestamp 1698431365
transform 1 0 77728 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_686
timestamp 1698431365
transform 1 0 78176 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42448 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 41104 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input3
timestamp 1698431365
transform -1 0 78400 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 37072 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 35840 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input6
timestamp 1698431365
transform -1 0 78400 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 78400 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input10
timestamp 1698431365
transform 1 0 1568 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 42560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 27328 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 47040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input15
timestamp 1698431365
transform 1 0 27328 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 49168 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 29008 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input18
timestamp 1698431365
transform -1 0 78400 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input19
timestamp 1698431365
transform 1 0 28336 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 78400 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input21
timestamp 1698431365
transform -1 0 55552 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input22
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 44128 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input25
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input26
timestamp 1698431365
transform -1 0 54656 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input28
timestamp 1698431365
transform -1 0 57232 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform -1 0 50848 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input30
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 24416 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input34
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output35
timestamp 1698431365
transform 1 0 77728 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output36 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 75488 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output37
timestamp 1698431365
transform 1 0 75488 0 -1 58016
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output38
timestamp 1698431365
transform -1 0 4480 0 1 67424
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output39
timestamp 1698431365
transform 1 0 51856 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output40
timestamp 1698431365
transform -1 0 25200 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output41
timestamp 1698431365
transform -1 0 4480 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output42
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output43
timestamp 1698431365
transform -1 0 29904 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output44
timestamp 1698431365
transform 1 0 58688 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output45
timestamp 1698431365
transform 1 0 52528 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output46
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output47
timestamp 1698431365
transform 1 0 43120 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output48
timestamp 1698431365
transform 1 0 75488 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output49
timestamp 1698431365
transform -1 0 40432 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output50
timestamp 1698431365
transform 1 0 40432 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51
timestamp 1698431365
transform 1 0 75488 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output52
timestamp 1698431365
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53
timestamp 1698431365
transform -1 0 4480 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698431365
transform 1 0 75488 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698431365
transform -1 0 4480 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698431365
transform 1 0 75488 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output57
timestamp 1698431365
transform -1 0 4480 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output58
timestamp 1698431365
transform -1 0 43232 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output59
timestamp 1698431365
transform 1 0 75488 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output60
timestamp 1698431365
transform -1 0 36624 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output61
timestamp 1698431365
transform -1 0 31136 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output62
timestamp 1698431365
transform 1 0 75488 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output63
timestamp 1698431365
transform 1 0 75488 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output64
timestamp 1698431365
transform 1 0 51072 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output65
timestamp 1698431365
transform -1 0 4480 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output66
timestamp 1698431365
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output67
timestamp 1698431365
transform -1 0 36624 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output68
timestamp 1698431365
transform 1 0 51184 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output69
timestamp 1698431365
transform -1 0 4480 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_94 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_136
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_137
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 78624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_138
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 78624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_139
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 78624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_140
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 78624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_141
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 78624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_142
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 78624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_143
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 78624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_144
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 78624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_145
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 78624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_146
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 78624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_147
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 78624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_148
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 78624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_149
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 78624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_150
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 78624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_151
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 78624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_152
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 78624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_153
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 78624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_154
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 78624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_155
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 78624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_156
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 78624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_157
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 78624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_158
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 78624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_159
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 78624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_160
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 78624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_161
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 78624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_162
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 78624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_163
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 78624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_164
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 78624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_165
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 78624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_166
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 78624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_167
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 78624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_168
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 78624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_169
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 78624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_170
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 78624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_171
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 78624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_172
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 78624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_173
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 78624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_174
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 78624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_175
timestamp 1698431365
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698431365
transform -1 0 78624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_176
timestamp 1698431365
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698431365
transform -1 0 78624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_177
timestamp 1698431365
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698431365
transform -1 0 78624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_178
timestamp 1698431365
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698431365
transform -1 0 78624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_179
timestamp 1698431365
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698431365
transform -1 0 78624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_180
timestamp 1698431365
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698431365
transform -1 0 78624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_181
timestamp 1698431365
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698431365
transform -1 0 78624 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_182
timestamp 1698431365
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698431365
transform -1 0 78624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_183
timestamp 1698431365
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698431365
transform -1 0 78624 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_184
timestamp 1698431365
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698431365
transform -1 0 78624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_185
timestamp 1698431365
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698431365
transform -1 0 78624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_186
timestamp 1698431365
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698431365
transform -1 0 78624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_187
timestamp 1698431365
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698431365
transform -1 0 78624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_188 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_189
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_190
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_191
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_192
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_193
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_194
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_195
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_196
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_197
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_198
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_199
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_200
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_201
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_202
timestamp 1698431365
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_203
timestamp 1698431365
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_204
timestamp 1698431365
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_205
timestamp 1698431365
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_206
timestamp 1698431365
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_207
timestamp 1698431365
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_208
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_209
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_210
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_211
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_212
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_213
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_214
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_215
timestamp 1698431365
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_216
timestamp 1698431365
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_217
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_218
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_219
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_220
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_221
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_222
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_223
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_224
timestamp 1698431365
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_225
timestamp 1698431365
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_226
timestamp 1698431365
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_227
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_228
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_229
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_230
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_231
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_232
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_233
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_234
timestamp 1698431365
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_235
timestamp 1698431365
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_236
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_237
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_238
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_239
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_240
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_241
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_242
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_243
timestamp 1698431365
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_244
timestamp 1698431365
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_245
timestamp 1698431365
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_246
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_247
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_248
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_249
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_250
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_251
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_252
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_253
timestamp 1698431365
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_254
timestamp 1698431365
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_255
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_256
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_257
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_258
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_259
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_260
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_261
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_262
timestamp 1698431365
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_263
timestamp 1698431365
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_264
timestamp 1698431365
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_265
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_266
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_267
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_268
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_269
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_270
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_271
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_272
timestamp 1698431365
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_273
timestamp 1698431365
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_274
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_275
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_276
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_277
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_278
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_279
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_280
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_281
timestamp 1698431365
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_282
timestamp 1698431365
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_283
timestamp 1698431365
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_284
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_285
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_286
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_287
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_288
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_289
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_290
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_291
timestamp 1698431365
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_292
timestamp 1698431365
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_293
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_294
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_295
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_296
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_297
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_298
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_299
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_300
timestamp 1698431365
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_301
timestamp 1698431365
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_302
timestamp 1698431365
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_303
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_304
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_305
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_306
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_307
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_308
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_309
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_310
timestamp 1698431365
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_311
timestamp 1698431365
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_312
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_313
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_314
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_315
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_316
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_317
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_318
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_319
timestamp 1698431365
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_320
timestamp 1698431365
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_321
timestamp 1698431365
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_322
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_323
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_324
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_325
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_326
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_327
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_328
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_329
timestamp 1698431365
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_330
timestamp 1698431365
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_331
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_332
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_333
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_334
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_335
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_336
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_337
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_338
timestamp 1698431365
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_339
timestamp 1698431365
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_340
timestamp 1698431365
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_341
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_342
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_343
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_344
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_345
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_346
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_347
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_348
timestamp 1698431365
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_349
timestamp 1698431365
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_350
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_351
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_352
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_353
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_354
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_355
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_356
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_357
timestamp 1698431365
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_358
timestamp 1698431365
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_359
timestamp 1698431365
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_360
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_361
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_362
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_363
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_364
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_365
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_366
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_367
timestamp 1698431365
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_368
timestamp 1698431365
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_369
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_370
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_371
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_372
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_373
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_374
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_375
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_376
timestamp 1698431365
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_377
timestamp 1698431365
transform 1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_378
timestamp 1698431365
transform 1 0 75824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_379
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_380
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_381
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_382
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_383
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_384
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_385
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_386
timestamp 1698431365
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_387
timestamp 1698431365
transform 1 0 71904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_388
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_389
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_390
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_391
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_392
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_393
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_394
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_395
timestamp 1698431365
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_396
timestamp 1698431365
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_397
timestamp 1698431365
transform 1 0 75824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_398
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_399
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_400
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_401
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_402
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_403
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_404
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_405
timestamp 1698431365
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_406
timestamp 1698431365
transform 1 0 71904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_407
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_408
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_409
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_410
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_411
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_412
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_413
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_414
timestamp 1698431365
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_415
timestamp 1698431365
transform 1 0 67984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_416
timestamp 1698431365
transform 1 0 75824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_417
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_418
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_419
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_420
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_421
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_422
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_423
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_424
timestamp 1698431365
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_425
timestamp 1698431365
transform 1 0 71904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_426
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_427
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_428
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_429
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_430
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_431
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_432
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_433
timestamp 1698431365
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_434
timestamp 1698431365
transform 1 0 67984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_435
timestamp 1698431365
transform 1 0 75824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_436
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_437
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_438
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_439
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_440
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_441
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_442
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_443
timestamp 1698431365
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_444
timestamp 1698431365
transform 1 0 71904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_445
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_446
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_447
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_448
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_449
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_450
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_451
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_452
timestamp 1698431365
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_453
timestamp 1698431365
transform 1 0 67984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_454
timestamp 1698431365
transform 1 0 75824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_455
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_456
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_457
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_458
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_459
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_460
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_461
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_462
timestamp 1698431365
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_463
timestamp 1698431365
transform 1 0 71904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_464
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_465
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_466
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_467
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_468
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_469
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_470
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_471
timestamp 1698431365
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_472
timestamp 1698431365
transform 1 0 67984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_473
timestamp 1698431365
transform 1 0 75824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_474
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_475
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_476
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_477
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_478
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_479
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_480
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_481
timestamp 1698431365
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_482
timestamp 1698431365
transform 1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_483
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_484
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_485
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_486
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_487
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_488
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_489
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_490
timestamp 1698431365
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_491
timestamp 1698431365
transform 1 0 67984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_492
timestamp 1698431365
transform 1 0 75824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_493
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_494
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_495
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_496
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_497
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_498
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_499
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_500
timestamp 1698431365
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_501
timestamp 1698431365
transform 1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_502
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_503
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_504
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_505
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_506
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_507
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_508
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_509
timestamp 1698431365
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_510
timestamp 1698431365
transform 1 0 67984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_511
timestamp 1698431365
transform 1 0 75824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_512
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_513
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_514
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_515
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_516
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_517
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_518
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_519
timestamp 1698431365
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_520
timestamp 1698431365
transform 1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_521
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_522
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_523
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_524
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_525
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_526
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_527
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_528
timestamp 1698431365
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_529
timestamp 1698431365
transform 1 0 67984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_530
timestamp 1698431365
transform 1 0 75824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_531
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_532
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_533
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_534
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_535
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_536
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_537
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_538
timestamp 1698431365
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_539
timestamp 1698431365
transform 1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_540
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_541
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_542
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_543
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_544
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_545
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_546
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_547
timestamp 1698431365
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_548
timestamp 1698431365
transform 1 0 67984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_549
timestamp 1698431365
transform 1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_550
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_551
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_552
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_553
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_554
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_555
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_556
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_557
timestamp 1698431365
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_558
timestamp 1698431365
transform 1 0 71904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_559
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_560
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_561
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_562
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_563
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_564
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_565
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_566
timestamp 1698431365
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_567
timestamp 1698431365
transform 1 0 67984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_568
timestamp 1698431365
transform 1 0 75824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_569
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_570
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_571
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_572
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_573
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_574
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_575
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_576
timestamp 1698431365
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_577
timestamp 1698431365
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_578
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_579
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_580
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_581
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_582
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_583
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_584
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_585
timestamp 1698431365
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_586
timestamp 1698431365
transform 1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_587
timestamp 1698431365
transform 1 0 75824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_588
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_589
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_590
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_591
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_592
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_593
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_594
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_595
timestamp 1698431365
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_596
timestamp 1698431365
transform 1 0 71904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_597
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_598
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_599
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_600
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_601
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_602
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_603
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_604
timestamp 1698431365
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_605
timestamp 1698431365
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_606
timestamp 1698431365
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_607
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_608
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_609
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_610
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_611
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_612
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_613
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_614
timestamp 1698431365
transform 1 0 64064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_615
timestamp 1698431365
transform 1 0 71904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_616
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_617
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_618
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_619
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_620
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_621
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_622
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_623
timestamp 1698431365
transform 1 0 60144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_624
timestamp 1698431365
transform 1 0 67984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_625
timestamp 1698431365
transform 1 0 75824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_626
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_627
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_628
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_629
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_630
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_631
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_632
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_633
timestamp 1698431365
transform 1 0 64064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_634
timestamp 1698431365
transform 1 0 71904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_635
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_636
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_637
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_638
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_639
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_640
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_641
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_642
timestamp 1698431365
transform 1 0 60144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_643
timestamp 1698431365
transform 1 0 67984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_644
timestamp 1698431365
transform 1 0 75824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_645
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_646
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_647
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_648
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_649
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_650
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_651
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_652
timestamp 1698431365
transform 1 0 64064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_653
timestamp 1698431365
transform 1 0 71904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_654
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_655
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_656
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_657
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_658
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_659
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_660
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_661
timestamp 1698431365
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_662
timestamp 1698431365
transform 1 0 67984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_663
timestamp 1698431365
transform 1 0 75824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_664
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_665
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_666
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_667
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_668
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_669
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_670
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_671
timestamp 1698431365
transform 1 0 64064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_672
timestamp 1698431365
transform 1 0 71904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_673
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_674
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_675
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_676
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_677
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_678
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_679
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_680
timestamp 1698431365
transform 1 0 60144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_681
timestamp 1698431365
transform 1 0 67984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_682
timestamp 1698431365
transform 1 0 75824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_683
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_684
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_685
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_686
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_687
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_688
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_689
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_690
timestamp 1698431365
transform 1 0 64064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_691
timestamp 1698431365
transform 1 0 71904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_692
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_693
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_694
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_695
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_696
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_697
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_698
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_699
timestamp 1698431365
transform 1 0 60144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_700
timestamp 1698431365
transform 1 0 67984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_701
timestamp 1698431365
transform 1 0 75824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_702
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_703
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_704
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_705
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_706
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_707
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_708
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_709
timestamp 1698431365
transform 1 0 64064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_710
timestamp 1698431365
transform 1 0 71904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_711
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_712
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_713
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_714
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_715
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_716
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_717
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_718
timestamp 1698431365
transform 1 0 60144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_719
timestamp 1698431365
transform 1 0 67984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_720
timestamp 1698431365
transform 1 0 75824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_721
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_722
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_723
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_724
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_725
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_726
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_727
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_728
timestamp 1698431365
transform 1 0 64064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_729
timestamp 1698431365
transform 1 0 71904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_730
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_731
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_732
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_733
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_734
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_735
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_736
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_737
timestamp 1698431365
transform 1 0 60144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_738
timestamp 1698431365
transform 1 0 67984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_739
timestamp 1698431365
transform 1 0 75824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_740
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_741
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_742
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_743
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_744
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_745
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_746
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_747
timestamp 1698431365
transform 1 0 64064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_748
timestamp 1698431365
transform 1 0 71904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_749
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_750
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_751
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_752
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_753
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_754
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_755
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_756
timestamp 1698431365
transform 1 0 60144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_757
timestamp 1698431365
transform 1 0 67984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_758
timestamp 1698431365
transform 1 0 75824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_759
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_760
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_761
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_762
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_763
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_764
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_765
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_766
timestamp 1698431365
transform 1 0 64064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_767
timestamp 1698431365
transform 1 0 71904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_768
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_769
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_770
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_771
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_772
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_773
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_774
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_775
timestamp 1698431365
transform 1 0 60144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_776
timestamp 1698431365
transform 1 0 67984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_777
timestamp 1698431365
transform 1 0 75824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_778
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_779
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_780
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_781
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_782
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_783
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_784
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_785
timestamp 1698431365
transform 1 0 64064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_786
timestamp 1698431365
transform 1 0 71904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_787
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_788
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_789
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_790
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_791
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_792
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_793
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_794
timestamp 1698431365
transform 1 0 60144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_795
timestamp 1698431365
transform 1 0 67984 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_796
timestamp 1698431365
transform 1 0 75824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_797
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_798
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_799
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_800
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_801
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_802
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_803
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_804
timestamp 1698431365
transform 1 0 64064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_805
timestamp 1698431365
transform 1 0 71904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_806
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_807
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_808
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_809
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_810
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_811
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_812
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_813
timestamp 1698431365
transform 1 0 60144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_814
timestamp 1698431365
transform 1 0 67984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_815
timestamp 1698431365
transform 1 0 75824 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_816
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_817
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_818
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_819
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_820
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_821
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_822
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_823
timestamp 1698431365
transform 1 0 64064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_824
timestamp 1698431365
transform 1 0 71904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_825
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_826
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_827
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_828
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_829
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_830
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_831
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_832
timestamp 1698431365
transform 1 0 60144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_833
timestamp 1698431365
transform 1 0 67984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_834
timestamp 1698431365
transform 1 0 75824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_835
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_836
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_837
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_838
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_839
timestamp 1698431365
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_840
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_841
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_842
timestamp 1698431365
transform 1 0 64064 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_843
timestamp 1698431365
transform 1 0 71904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_844
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_845
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_846
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_847
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_848
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_849
timestamp 1698431365
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_850
timestamp 1698431365
transform 1 0 52304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_851
timestamp 1698431365
transform 1 0 60144 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_852
timestamp 1698431365
transform 1 0 67984 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_853
timestamp 1698431365
transform 1 0 75824 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_854
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_855
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_856
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_857
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_858
timestamp 1698431365
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_859
timestamp 1698431365
transform 1 0 48384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_860
timestamp 1698431365
transform 1 0 56224 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_861
timestamp 1698431365
transform 1 0 64064 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_862
timestamp 1698431365
transform 1 0 71904 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_863
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_864
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_865
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_866
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_867
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_868
timestamp 1698431365
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_869
timestamp 1698431365
transform 1 0 52304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_870
timestamp 1698431365
transform 1 0 60144 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_871
timestamp 1698431365
transform 1 0 67984 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_872
timestamp 1698431365
transform 1 0 75824 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_873
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_874
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_875
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_876
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_877
timestamp 1698431365
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_878
timestamp 1698431365
transform 1 0 48384 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_879
timestamp 1698431365
transform 1 0 56224 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_880
timestamp 1698431365
transform 1 0 64064 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_881
timestamp 1698431365
transform 1 0 71904 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_882
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_883
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_884
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_885
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_886
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_887
timestamp 1698431365
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_888
timestamp 1698431365
transform 1 0 52304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_889
timestamp 1698431365
transform 1 0 60144 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_890
timestamp 1698431365
transform 1 0 67984 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_891
timestamp 1698431365
transform 1 0 75824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_892
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_893
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_894
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_895
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_896
timestamp 1698431365
transform 1 0 40544 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_897
timestamp 1698431365
transform 1 0 48384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_898
timestamp 1698431365
transform 1 0 56224 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_899
timestamp 1698431365
transform 1 0 64064 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_900
timestamp 1698431365
transform 1 0 71904 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_901
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_902
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_903
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_904
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_905
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_906
timestamp 1698431365
transform 1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_907
timestamp 1698431365
transform 1 0 52304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_908
timestamp 1698431365
transform 1 0 60144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_909
timestamp 1698431365
transform 1 0 67984 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_910
timestamp 1698431365
transform 1 0 75824 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_911
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_912
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_913
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_914
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_915
timestamp 1698431365
transform 1 0 40544 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_916
timestamp 1698431365
transform 1 0 48384 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_917
timestamp 1698431365
transform 1 0 56224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_918
timestamp 1698431365
transform 1 0 64064 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_919
timestamp 1698431365
transform 1 0 71904 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_920
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_921
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_922
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_923
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_924
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_925
timestamp 1698431365
transform 1 0 44464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_926
timestamp 1698431365
transform 1 0 52304 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_927
timestamp 1698431365
transform 1 0 60144 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_928
timestamp 1698431365
transform 1 0 67984 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_929
timestamp 1698431365
transform 1 0 75824 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_930
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_931
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_932
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_933
timestamp 1698431365
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_934
timestamp 1698431365
transform 1 0 40544 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_935
timestamp 1698431365
transform 1 0 48384 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_936
timestamp 1698431365
transform 1 0 56224 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_937
timestamp 1698431365
transform 1 0 64064 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_938
timestamp 1698431365
transform 1 0 71904 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_939
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_940
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_941
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_942
timestamp 1698431365
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_943
timestamp 1698431365
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_944
timestamp 1698431365
transform 1 0 44464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_945
timestamp 1698431365
transform 1 0 52304 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_946
timestamp 1698431365
transform 1 0 60144 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_947
timestamp 1698431365
transform 1 0 67984 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_948
timestamp 1698431365
transform 1 0 75824 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_949
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_950
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_951
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_952
timestamp 1698431365
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_953
timestamp 1698431365
transform 1 0 40544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_954
timestamp 1698431365
transform 1 0 48384 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_955
timestamp 1698431365
transform 1 0 56224 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_956
timestamp 1698431365
transform 1 0 64064 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_957
timestamp 1698431365
transform 1 0 71904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_958
timestamp 1698431365
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_959
timestamp 1698431365
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_960
timestamp 1698431365
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_961
timestamp 1698431365
transform 1 0 28784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_962
timestamp 1698431365
transform 1 0 36624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_963
timestamp 1698431365
transform 1 0 44464 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_964
timestamp 1698431365
transform 1 0 52304 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_965
timestamp 1698431365
transform 1 0 60144 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_966
timestamp 1698431365
transform 1 0 67984 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_967
timestamp 1698431365
transform 1 0 75824 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_968
timestamp 1698431365
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_969
timestamp 1698431365
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_970
timestamp 1698431365
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_971
timestamp 1698431365
transform 1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_972
timestamp 1698431365
transform 1 0 40544 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_973
timestamp 1698431365
transform 1 0 48384 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_974
timestamp 1698431365
transform 1 0 56224 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_975
timestamp 1698431365
transform 1 0 64064 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_976
timestamp 1698431365
transform 1 0 71904 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_977
timestamp 1698431365
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_978
timestamp 1698431365
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_979
timestamp 1698431365
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_980
timestamp 1698431365
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_981
timestamp 1698431365
transform 1 0 36624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_982
timestamp 1698431365
transform 1 0 44464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_983
timestamp 1698431365
transform 1 0 52304 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_984
timestamp 1698431365
transform 1 0 60144 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_985
timestamp 1698431365
transform 1 0 67984 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_986
timestamp 1698431365
transform 1 0 75824 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_987
timestamp 1698431365
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_988
timestamp 1698431365
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_989
timestamp 1698431365
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_990
timestamp 1698431365
transform 1 0 32704 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_991
timestamp 1698431365
transform 1 0 40544 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_992
timestamp 1698431365
transform 1 0 48384 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_993
timestamp 1698431365
transform 1 0 56224 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_994
timestamp 1698431365
transform 1 0 64064 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_995
timestamp 1698431365
transform 1 0 71904 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_996
timestamp 1698431365
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_997
timestamp 1698431365
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_998
timestamp 1698431365
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_999
timestamp 1698431365
transform 1 0 28784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1000
timestamp 1698431365
transform 1 0 36624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1001
timestamp 1698431365
transform 1 0 44464 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1002
timestamp 1698431365
transform 1 0 52304 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1003
timestamp 1698431365
transform 1 0 60144 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1004
timestamp 1698431365
transform 1 0 67984 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1005
timestamp 1698431365
transform 1 0 75824 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1006
timestamp 1698431365
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1007
timestamp 1698431365
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1008
timestamp 1698431365
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1009
timestamp 1698431365
transform 1 0 32704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1010
timestamp 1698431365
transform 1 0 40544 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1011
timestamp 1698431365
transform 1 0 48384 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1012
timestamp 1698431365
transform 1 0 56224 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1013
timestamp 1698431365
transform 1 0 64064 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1014
timestamp 1698431365
transform 1 0 71904 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1015
timestamp 1698431365
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1016
timestamp 1698431365
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1017
timestamp 1698431365
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1018
timestamp 1698431365
transform 1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1019
timestamp 1698431365
transform 1 0 36624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1020
timestamp 1698431365
transform 1 0 44464 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1021
timestamp 1698431365
transform 1 0 52304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1022
timestamp 1698431365
transform 1 0 60144 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1023
timestamp 1698431365
transform 1 0 67984 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1024
timestamp 1698431365
transform 1 0 75824 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1025
timestamp 1698431365
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1026
timestamp 1698431365
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1027
timestamp 1698431365
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1028
timestamp 1698431365
transform 1 0 32704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1029
timestamp 1698431365
transform 1 0 40544 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1030
timestamp 1698431365
transform 1 0 48384 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1031
timestamp 1698431365
transform 1 0 56224 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1032
timestamp 1698431365
transform 1 0 64064 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1033
timestamp 1698431365
transform 1 0 71904 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1034
timestamp 1698431365
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1035
timestamp 1698431365
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1036
timestamp 1698431365
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1037
timestamp 1698431365
transform 1 0 28784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1038
timestamp 1698431365
transform 1 0 36624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1039
timestamp 1698431365
transform 1 0 44464 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1040
timestamp 1698431365
transform 1 0 52304 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1041
timestamp 1698431365
transform 1 0 60144 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1042
timestamp 1698431365
transform 1 0 67984 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1043
timestamp 1698431365
transform 1 0 75824 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1044
timestamp 1698431365
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1045
timestamp 1698431365
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1046
timestamp 1698431365
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1047
timestamp 1698431365
transform 1 0 32704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1048
timestamp 1698431365
transform 1 0 40544 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1049
timestamp 1698431365
transform 1 0 48384 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1050
timestamp 1698431365
transform 1 0 56224 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1051
timestamp 1698431365
transform 1 0 64064 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1052
timestamp 1698431365
transform 1 0 71904 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1053
timestamp 1698431365
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1054
timestamp 1698431365
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1055
timestamp 1698431365
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1056
timestamp 1698431365
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1057
timestamp 1698431365
transform 1 0 36624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1058
timestamp 1698431365
transform 1 0 44464 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1059
timestamp 1698431365
transform 1 0 52304 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1060
timestamp 1698431365
transform 1 0 60144 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1061
timestamp 1698431365
transform 1 0 67984 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1062
timestamp 1698431365
transform 1 0 75824 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1063
timestamp 1698431365
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1064
timestamp 1698431365
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1065
timestamp 1698431365
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1066
timestamp 1698431365
transform 1 0 32704 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1067
timestamp 1698431365
transform 1 0 40544 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1068
timestamp 1698431365
transform 1 0 48384 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1069
timestamp 1698431365
transform 1 0 56224 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1070
timestamp 1698431365
transform 1 0 64064 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1071
timestamp 1698431365
transform 1 0 71904 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1072
timestamp 1698431365
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1073
timestamp 1698431365
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1074
timestamp 1698431365
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1075
timestamp 1698431365
transform 1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1076
timestamp 1698431365
transform 1 0 36624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1077
timestamp 1698431365
transform 1 0 44464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1078
timestamp 1698431365
transform 1 0 52304 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1079
timestamp 1698431365
transform 1 0 60144 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1080
timestamp 1698431365
transform 1 0 67984 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1081
timestamp 1698431365
transform 1 0 75824 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1082
timestamp 1698431365
transform 1 0 5152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1083
timestamp 1698431365
transform 1 0 8960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1084
timestamp 1698431365
transform 1 0 12768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1085
timestamp 1698431365
transform 1 0 16576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1086
timestamp 1698431365
transform 1 0 20384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1087
timestamp 1698431365
transform 1 0 24192 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1088
timestamp 1698431365
transform 1 0 28000 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1089
timestamp 1698431365
transform 1 0 31808 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1090
timestamp 1698431365
transform 1 0 35616 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1091
timestamp 1698431365
transform 1 0 39424 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1092
timestamp 1698431365
transform 1 0 43232 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1093
timestamp 1698431365
transform 1 0 47040 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1094
timestamp 1698431365
transform 1 0 50848 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1095
timestamp 1698431365
transform 1 0 54656 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1096
timestamp 1698431365
transform 1 0 58464 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1097
timestamp 1698431365
transform 1 0 62272 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1098
timestamp 1698431365
transform 1 0 66080 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1099
timestamp 1698431365
transform 1 0 69888 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1100
timestamp 1698431365
transform 1 0 73696 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1101
timestamp 1698431365
transform 1 0 77504 0 -1 76832
box -86 -86 310 870
<< labels >>
flabel metal3 s 79200 58464 80000 58576 0 FreeSans 448 0 0 0 clk
port 0 nsew signal tristate
flabel metal3 s 79200 20160 80000 20272 0 FreeSans 448 0 0 0 in[0]
port 1 nsew signal tristate
flabel metal3 s 79200 57792 80000 57904 0 FreeSans 448 0 0 0 in[10]
port 2 nsew signal tristate
flabel metal3 s 0 67200 800 67312 0 FreeSans 448 0 0 0 in[11]
port 3 nsew signal tristate
flabel metal2 s 51744 0 51856 800 0 FreeSans 448 90 0 0 in[12]
port 4 nsew signal tristate
flabel metal2 s 22176 79200 22288 80000 0 FreeSans 448 90 0 0 in[13]
port 5 nsew signal tristate
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 in[14]
port 6 nsew signal tristate
flabel metal2 s 50400 0 50512 800 0 FreeSans 448 90 0 0 in[15]
port 7 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 in[16]
port 8 nsew signal tristate
flabel metal2 s 58464 79200 58576 80000 0 FreeSans 448 90 0 0 in[17]
port 9 nsew signal tristate
flabel metal2 s 51744 79200 51856 80000 0 FreeSans 448 90 0 0 in[1]
port 10 nsew signal tristate
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 in[2]
port 11 nsew signal tristate
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 in[3]
port 12 nsew signal tristate
flabel metal3 s 79200 24864 80000 24976 0 FreeSans 448 0 0 0 in[4]
port 13 nsew signal tristate
flabel metal2 s 38304 79200 38416 80000 0 FreeSans 448 90 0 0 in[5]
port 14 nsew signal tristate
flabel metal2 s 40320 79200 40432 80000 0 FreeSans 448 90 0 0 in[6]
port 15 nsew signal tristate
flabel metal3 s 79200 21504 80000 21616 0 FreeSans 448 0 0 0 in[7]
port 16 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 in[8]
port 17 nsew signal tristate
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 in[9]
port 18 nsew signal tristate
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 io_in[0]
port 19 nsew signal input
flabel metal2 s 41664 0 41776 800 0 FreeSans 448 90 0 0 io_in[10]
port 20 nsew signal input
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 io_in[11]
port 21 nsew signal input
flabel metal3 s 79200 26208 80000 26320 0 FreeSans 448 0 0 0 io_in[12]
port 22 nsew signal input
flabel metal2 s 36960 79200 37072 80000 0 FreeSans 448 90 0 0 io_in[13]
port 23 nsew signal input
flabel metal2 s 35616 79200 35728 80000 0 FreeSans 448 90 0 0 io_in[14]
port 24 nsew signal input
flabel metal3 s 79200 20832 80000 20944 0 FreeSans 448 0 0 0 io_in[15]
port 25 nsew signal input
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 io_in[16]
port 26 nsew signal input
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 io_in[17]
port 27 nsew signal input
flabel metal3 s 79200 51072 80000 51184 0 FreeSans 448 0 0 0 io_in[18]
port 28 nsew signal input
flabel metal3 s 0 64512 800 64624 0 FreeSans 448 0 0 0 io_in[19]
port 29 nsew signal input
flabel metal2 s 65184 0 65296 800 0 FreeSans 448 90 0 0 io_in[1]
port 30 nsew signal input
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 io_in[20]
port 31 nsew signal input
flabel metal2 s 28224 79200 28336 80000 0 FreeSans 448 90 0 0 io_in[21]
port 32 nsew signal input
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 io_in[22]
port 33 nsew signal input
flabel metal2 s 44352 0 44464 800 0 FreeSans 448 90 0 0 io_in[23]
port 34 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 io_in[24]
port 35 nsew signal input
flabel metal2 s 48384 79200 48496 80000 0 FreeSans 448 90 0 0 io_in[25]
port 36 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 io_in[26]
port 37 nsew signal input
flabel metal2 s 67200 0 67312 800 0 FreeSans 448 90 0 0 io_in[27]
port 38 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 io_in[28]
port 39 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 io_in[29]
port 40 nsew signal input
flabel metal2 s 73248 0 73360 800 0 FreeSans 448 90 0 0 io_in[2]
port 41 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 io_in[30]
port 42 nsew signal input
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 io_in[31]
port 43 nsew signal input
flabel metal2 s 56448 0 56560 800 0 FreeSans 448 90 0 0 io_in[32]
port 44 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 io_in[33]
port 45 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 io_in[34]
port 46 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 io_in[35]
port 47 nsew signal input
flabel metal2 s 58464 0 58576 800 0 FreeSans 448 90 0 0 io_in[36]
port 48 nsew signal input
flabel metal2 s 59808 0 59920 800 0 FreeSans 448 90 0 0 io_in[37]
port 49 nsew signal input
flabel metal2 s 59136 0 59248 800 0 FreeSans 448 90 0 0 io_in[3]
port 50 nsew signal input
flabel metal2 s 77280 0 77392 800 0 FreeSans 448 90 0 0 io_in[4]
port 51 nsew signal input
flabel metal2 s 28896 79200 29008 80000 0 FreeSans 448 90 0 0 io_in[5]
port 52 nsew signal input
flabel metal3 s 79200 56448 80000 56560 0 FreeSans 448 0 0 0 io_in[6]
port 53 nsew signal input
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 io_in[7]
port 54 nsew signal input
flabel metal3 s 79200 33600 80000 33712 0 FreeSans 448 0 0 0 io_in[8]
port 55 nsew signal input
flabel metal2 s 54432 79200 54544 80000 0 FreeSans 448 90 0 0 io_in[9]
port 56 nsew signal input
flabel metal2 s 46368 79200 46480 80000 0 FreeSans 448 90 0 0 io_oeb[0]
port 57 nsew signal tristate
flabel metal2 s 31584 79200 31696 80000 0 FreeSans 448 90 0 0 io_oeb[10]
port 58 nsew signal tristate
flabel metal3 s 79200 57120 80000 57232 0 FreeSans 448 0 0 0 io_oeb[11]
port 59 nsew signal tristate
flabel metal3 s 79200 53088 80000 53200 0 FreeSans 448 0 0 0 io_oeb[12]
port 60 nsew signal tristate
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 io_oeb[13]
port 61 nsew signal tristate
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 io_oeb[14]
port 62 nsew signal tristate
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 io_oeb[15]
port 63 nsew signal tristate
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 io_oeb[16]
port 64 nsew signal tristate
flabel metal3 s 79200 34944 80000 35056 0 FreeSans 448 0 0 0 io_oeb[17]
port 65 nsew signal tristate
flabel metal3 s 79200 38976 80000 39088 0 FreeSans 448 0 0 0 io_oeb[18]
port 66 nsew signal tristate
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 io_oeb[19]
port 67 nsew signal tristate
flabel metal3 s 0 63840 800 63952 0 FreeSans 448 0 0 0 io_oeb[1]
port 68 nsew signal tristate
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 io_oeb[20]
port 69 nsew signal tristate
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 io_oeb[21]
port 70 nsew signal tristate
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 io_oeb[22]
port 71 nsew signal tristate
flabel metal3 s 79200 30912 80000 31024 0 FreeSans 448 0 0 0 io_oeb[23]
port 72 nsew signal tristate
flabel metal3 s 0 54432 800 54544 0 FreeSans 448 0 0 0 io_oeb[24]
port 73 nsew signal tristate
flabel metal3 s 79200 35616 80000 35728 0 FreeSans 448 0 0 0 io_oeb[25]
port 74 nsew signal tristate
flabel metal3 s 79200 40992 80000 41104 0 FreeSans 448 0 0 0 io_oeb[26]
port 75 nsew signal tristate
flabel metal3 s 79200 32256 80000 32368 0 FreeSans 448 0 0 0 io_oeb[27]
port 76 nsew signal tristate
flabel metal2 s 53088 79200 53200 80000 0 FreeSans 448 90 0 0 io_oeb[28]
port 77 nsew signal tristate
flabel metal2 s 24864 79200 24976 80000 0 FreeSans 448 90 0 0 io_oeb[29]
port 78 nsew signal tristate
flabel metal2 s 38976 79200 39088 80000 0 FreeSans 448 90 0 0 io_oeb[2]
port 79 nsew signal tristate
flabel metal3 s 79200 45696 80000 45808 0 FreeSans 448 0 0 0 io_oeb[30]
port 80 nsew signal tristate
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 io_oeb[31]
port 81 nsew signal tristate
flabel metal3 s 79200 24192 80000 24304 0 FreeSans 448 0 0 0 io_oeb[32]
port 82 nsew signal tristate
flabel metal3 s 79200 43680 80000 43792 0 FreeSans 448 0 0 0 io_oeb[33]
port 83 nsew signal tristate
flabel metal3 s 79200 43008 80000 43120 0 FreeSans 448 0 0 0 io_oeb[34]
port 84 nsew signal tristate
flabel metal2 s 32256 79200 32368 80000 0 FreeSans 448 90 0 0 io_oeb[35]
port 85 nsew signal tristate
flabel metal2 s 30912 79200 31024 80000 0 FreeSans 448 90 0 0 io_oeb[36]
port 86 nsew signal tristate
flabel metal3 s 0 61824 800 61936 0 FreeSans 448 0 0 0 io_oeb[37]
port 87 nsew signal tristate
flabel metal2 s 30240 79200 30352 80000 0 FreeSans 448 90 0 0 io_oeb[3]
port 88 nsew signal tristate
flabel metal3 s 79200 38304 80000 38416 0 FreeSans 448 0 0 0 io_oeb[4]
port 89 nsew signal tristate
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 io_oeb[5]
port 90 nsew signal tristate
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 io_oeb[6]
port 91 nsew signal tristate
flabel metal2 s 34272 79200 34384 80000 0 FreeSans 448 90 0 0 io_oeb[7]
port 92 nsew signal tristate
flabel metal3 s 79200 52416 80000 52528 0 FreeSans 448 0 0 0 io_oeb[8]
port 93 nsew signal tristate
flabel metal2 s 49056 79200 49168 80000 0 FreeSans 448 90 0 0 io_oeb[9]
port 94 nsew signal tristate
flabel metal3 s 79200 36960 80000 37072 0 FreeSans 448 0 0 0 io_out[0]
port 95 nsew signal tristate
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 io_out[10]
port 96 nsew signal tristate
flabel metal3 s 0 45024 800 45136 0 FreeSans 448 0 0 0 io_out[11]
port 97 nsew signal tristate
flabel metal3 s 0 62496 800 62608 0 FreeSans 448 0 0 0 io_out[12]
port 98 nsew signal tristate
flabel metal3 s 79200 49056 80000 49168 0 FreeSans 448 0 0 0 io_out[13]
port 99 nsew signal tristate
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 io_out[14]
port 100 nsew signal tristate
flabel metal3 s 0 38976 800 39088 0 FreeSans 448 0 0 0 io_out[15]
port 101 nsew signal tristate
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 io_out[16]
port 102 nsew signal tristate
flabel metal3 s 79200 36288 80000 36400 0 FreeSans 448 0 0 0 io_out[17]
port 103 nsew signal tristate
flabel metal2 s 55104 79200 55216 80000 0 FreeSans 448 90 0 0 io_out[18]
port 104 nsew signal tristate
flabel metal3 s 0 42336 800 42448 0 FreeSans 448 0 0 0 io_out[19]
port 105 nsew signal tristate
flabel metal3 s 79200 37632 80000 37744 0 FreeSans 448 0 0 0 io_out[1]
port 106 nsew signal tristate
flabel metal2 s 25536 79200 25648 80000 0 FreeSans 448 90 0 0 io_out[20]
port 107 nsew signal tristate
flabel metal2 s 22848 79200 22960 80000 0 FreeSans 448 90 0 0 io_out[21]
port 108 nsew signal tristate
flabel metal2 s 26880 79200 26992 80000 0 FreeSans 448 90 0 0 io_out[22]
port 109 nsew signal tristate
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 io_out[23]
port 110 nsew signal tristate
flabel metal3 s 79200 32928 80000 33040 0 FreeSans 448 0 0 0 io_out[24]
port 111 nsew signal tristate
flabel metal2 s 46368 0 46480 800 0 FreeSans 448 90 0 0 io_out[25]
port 112 nsew signal tristate
flabel metal3 s 79200 30240 80000 30352 0 FreeSans 448 0 0 0 io_out[26]
port 113 nsew signal tristate
flabel metal3 s 0 41664 800 41776 0 FreeSans 448 0 0 0 io_out[27]
port 114 nsew signal tristate
flabel metal3 s 79200 53760 80000 53872 0 FreeSans 448 0 0 0 io_out[28]
port 115 nsew signal tristate
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 io_out[29]
port 116 nsew signal tristate
flabel metal3 s 79200 40320 80000 40432 0 FreeSans 448 0 0 0 io_out[2]
port 117 nsew signal tristate
flabel metal2 s 40992 79200 41104 80000 0 FreeSans 448 90 0 0 io_out[30]
port 118 nsew signal tristate
flabel metal3 s 79200 47040 80000 47152 0 FreeSans 448 0 0 0 io_out[31]
port 119 nsew signal tristate
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 io_out[32]
port 120 nsew signal tristate
flabel metal2 s 27552 79200 27664 80000 0 FreeSans 448 90 0 0 io_out[33]
port 121 nsew signal tristate
flabel metal3 s 79200 25536 80000 25648 0 FreeSans 448 0 0 0 io_out[34]
port 122 nsew signal tristate
flabel metal3 s 79200 22848 80000 22960 0 FreeSans 448 0 0 0 io_out[35]
port 123 nsew signal tristate
flabel metal2 s 49728 79200 49840 80000 0 FreeSans 448 90 0 0 io_out[36]
port 124 nsew signal tristate
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 io_out[37]
port 125 nsew signal tristate
flabel metal3 s 79200 55776 80000 55888 0 FreeSans 448 0 0 0 io_out[3]
port 126 nsew signal tristate
flabel metal3 s 79200 55104 80000 55216 0 FreeSans 448 0 0 0 io_out[4]
port 127 nsew signal tristate
flabel metal3 s 79200 44352 80000 44464 0 FreeSans 448 0 0 0 io_out[5]
port 128 nsew signal tristate
flabel metal2 s 51072 0 51184 800 0 FreeSans 448 90 0 0 io_out[6]
port 129 nsew signal tristate
flabel metal3 s 79200 49728 80000 49840 0 FreeSans 448 0 0 0 io_out[7]
port 130 nsew signal tristate
flabel metal2 s 45696 79200 45808 80000 0 FreeSans 448 90 0 0 io_out[8]
port 131 nsew signal tristate
flabel metal3 s 79200 39648 80000 39760 0 FreeSans 448 0 0 0 io_out[9]
port 132 nsew signal tristate
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 la_data_in[0]
port 133 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 la_data_in[10]
port 134 nsew signal input
flabel metal2 s 60480 0 60592 800 0 FreeSans 448 90 0 0 la_data_in[11]
port 135 nsew signal input
flabel metal2 s 55104 0 55216 800 0 FreeSans 448 90 0 0 la_data_in[12]
port 136 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 la_data_in[13]
port 137 nsew signal input
flabel metal2 s 67872 0 67984 800 0 FreeSans 448 90 0 0 la_data_in[14]
port 138 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 la_data_in[15]
port 139 nsew signal input
flabel metal2 s 74592 0 74704 800 0 FreeSans 448 90 0 0 la_data_in[16]
port 140 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 la_data_in[17]
port 141 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 la_data_in[18]
port 142 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 la_data_in[19]
port 143 nsew signal input
flabel metal2 s 78624 0 78736 800 0 FreeSans 448 90 0 0 la_data_in[1]
port 144 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 la_data_in[20]
port 145 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 la_data_in[21]
port 146 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 la_data_in[22]
port 147 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 la_data_in[23]
port 148 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 la_data_in[24]
port 149 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 la_data_in[25]
port 150 nsew signal input
flabel metal2 s 65856 0 65968 800 0 FreeSans 448 90 0 0 la_data_in[26]
port 151 nsew signal input
flabel metal2 s 79296 0 79408 800 0 FreeSans 448 90 0 0 la_data_in[27]
port 152 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 la_data_in[28]
port 153 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 la_data_in[29]
port 154 nsew signal input
flabel metal2 s 57120 0 57232 800 0 FreeSans 448 90 0 0 la_data_in[2]
port 155 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 la_data_in[30]
port 156 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 la_data_in[31]
port 157 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 la_data_in[32]
port 158 nsew signal input
flabel metal2 s 53760 0 53872 800 0 FreeSans 448 90 0 0 la_data_in[33]
port 159 nsew signal input
flabel metal2 s 71904 0 72016 800 0 FreeSans 448 90 0 0 la_data_in[34]
port 160 nsew signal input
flabel metal2 s 62496 0 62608 800 0 FreeSans 448 90 0 0 la_data_in[35]
port 161 nsew signal input
flabel metal2 s 57792 0 57904 800 0 FreeSans 448 90 0 0 la_data_in[36]
port 162 nsew signal input
flabel metal2 s 52416 0 52528 800 0 FreeSans 448 90 0 0 la_data_in[37]
port 163 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 la_data_in[38]
port 164 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 la_data_in[39]
port 165 nsew signal input
flabel metal2 s 64512 0 64624 800 0 FreeSans 448 90 0 0 la_data_in[3]
port 166 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 la_data_in[40]
port 167 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 la_data_in[41]
port 168 nsew signal input
flabel metal2 s 72576 0 72688 800 0 FreeSans 448 90 0 0 la_data_in[42]
port 169 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 la_data_in[43]
port 170 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 la_data_in[44]
port 171 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 la_data_in[45]
port 172 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 la_data_in[46]
port 173 nsew signal input
flabel metal2 s 63840 0 63952 800 0 FreeSans 448 90 0 0 la_data_in[47]
port 174 nsew signal input
flabel metal2 s 76608 0 76720 800 0 FreeSans 448 90 0 0 la_data_in[48]
port 175 nsew signal input
flabel metal2 s 63168 0 63280 800 0 FreeSans 448 90 0 0 la_data_in[49]
port 176 nsew signal input
flabel metal2 s 69888 0 70000 800 0 FreeSans 448 90 0 0 la_data_in[4]
port 177 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 la_data_in[50]
port 178 nsew signal input
flabel metal2 s 66528 0 66640 800 0 FreeSans 448 90 0 0 la_data_in[51]
port 179 nsew signal input
flabel metal2 s 73920 0 74032 800 0 FreeSans 448 90 0 0 la_data_in[52]
port 180 nsew signal input
flabel metal2 s 75264 0 75376 800 0 FreeSans 448 90 0 0 la_data_in[53]
port 181 nsew signal input
flabel metal2 s 68544 0 68656 800 0 FreeSans 448 90 0 0 la_data_in[54]
port 182 nsew signal input
flabel metal2 s 53088 0 53200 800 0 FreeSans 448 90 0 0 la_data_in[55]
port 183 nsew signal input
flabel metal2 s 71232 0 71344 800 0 FreeSans 448 90 0 0 la_data_in[56]
port 184 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 la_data_in[57]
port 185 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 la_data_in[58]
port 186 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 la_data_in[59]
port 187 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 la_data_in[5]
port 188 nsew signal input
flabel metal2 s 75936 0 76048 800 0 FreeSans 448 90 0 0 la_data_in[60]
port 189 nsew signal input
flabel metal2 s 61824 0 61936 800 0 FreeSans 448 90 0 0 la_data_in[61]
port 190 nsew signal input
flabel metal2 s 70560 0 70672 800 0 FreeSans 448 90 0 0 la_data_in[62]
port 191 nsew signal input
flabel metal2 s 55776 0 55888 800 0 FreeSans 448 90 0 0 la_data_in[63]
port 192 nsew signal input
flabel metal2 s 54432 0 54544 800 0 FreeSans 448 90 0 0 la_data_in[6]
port 193 nsew signal input
flabel metal2 s 69216 0 69328 800 0 FreeSans 448 90 0 0 la_data_in[7]
port 194 nsew signal input
flabel metal2 s 61152 0 61264 800 0 FreeSans 448 90 0 0 la_data_in[8]
port 195 nsew signal input
flabel metal2 s 77952 0 78064 800 0 FreeSans 448 90 0 0 la_data_in[9]
port 196 nsew signal input
flabel metal3 s 79200 46368 80000 46480 0 FreeSans 448 0 0 0 la_data_out[0]
port 197 nsew signal tristate
flabel metal3 s 79200 23520 80000 23632 0 FreeSans 448 0 0 0 la_data_out[10]
port 198 nsew signal tristate
flabel metal3 s 0 53760 800 53872 0 FreeSans 448 0 0 0 la_data_out[11]
port 199 nsew signal tristate
flabel metal2 s 57120 79200 57232 80000 0 FreeSans 448 90 0 0 la_data_out[12]
port 200 nsew signal tristate
flabel metal3 s 79200 27552 80000 27664 0 FreeSans 448 0 0 0 la_data_out[13]
port 201 nsew signal tristate
flabel metal3 s 79200 29568 80000 29680 0 FreeSans 448 0 0 0 la_data_out[14]
port 202 nsew signal tristate
flabel metal2 s 39648 79200 39760 80000 0 FreeSans 448 90 0 0 la_data_out[15]
port 203 nsew signal tristate
flabel metal3 s 79200 54432 80000 54544 0 FreeSans 448 0 0 0 la_data_out[16]
port 204 nsew signal tristate
flabel metal2 s 49728 0 49840 800 0 FreeSans 448 90 0 0 la_data_out[17]
port 205 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 la_data_out[18]
port 206 nsew signal tristate
flabel metal2 s 47712 0 47824 800 0 FreeSans 448 90 0 0 la_data_out[19]
port 207 nsew signal tristate
flabel metal2 s 47712 79200 47824 80000 0 FreeSans 448 90 0 0 la_data_out[1]
port 208 nsew signal tristate
flabel metal2 s 45024 79200 45136 80000 0 FreeSans 448 90 0 0 la_data_out[20]
port 209 nsew signal tristate
flabel metal3 s 0 59808 800 59920 0 FreeSans 448 0 0 0 la_data_out[21]
port 210 nsew signal tristate
flabel metal2 s 29568 79200 29680 80000 0 FreeSans 448 90 0 0 la_data_out[22]
port 211 nsew signal tristate
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 la_data_out[23]
port 212 nsew signal tristate
flabel metal2 s 49056 0 49168 800 0 FreeSans 448 90 0 0 la_data_out[24]
port 213 nsew signal tristate
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 la_data_out[25]
port 214 nsew signal tristate
flabel metal3 s 79200 22176 80000 22288 0 FreeSans 448 0 0 0 la_data_out[26]
port 215 nsew signal tristate
flabel metal3 s 79200 34272 80000 34384 0 FreeSans 448 0 0 0 la_data_out[27]
port 216 nsew signal tristate
flabel metal3 s 0 43008 800 43120 0 FreeSans 448 0 0 0 la_data_out[28]
port 217 nsew signal tristate
flabel metal2 s 42336 79200 42448 80000 0 FreeSans 448 90 0 0 la_data_out[29]
port 218 nsew signal tristate
flabel metal3 s 0 56448 800 56560 0 FreeSans 448 0 0 0 la_data_out[2]
port 219 nsew signal tristate
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 la_data_out[30]
port 220 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 la_data_out[31]
port 221 nsew signal tristate
flabel metal2 s 48384 0 48496 800 0 FreeSans 448 90 0 0 la_data_out[32]
port 222 nsew signal tristate
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 la_data_out[33]
port 223 nsew signal tristate
flabel metal2 s 32928 79200 33040 80000 0 FreeSans 448 90 0 0 la_data_out[34]
port 224 nsew signal tristate
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 la_data_out[35]
port 225 nsew signal tristate
flabel metal3 s 79200 51744 80000 51856 0 FreeSans 448 0 0 0 la_data_out[36]
port 226 nsew signal tristate
flabel metal2 s 45024 0 45136 800 0 FreeSans 448 90 0 0 la_data_out[37]
port 227 nsew signal tristate
flabel metal2 s 55776 79200 55888 80000 0 FreeSans 448 90 0 0 la_data_out[38]
port 228 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 la_data_out[39]
port 229 nsew signal tristate
flabel metal2 s 41664 79200 41776 80000 0 FreeSans 448 90 0 0 la_data_out[3]
port 230 nsew signal tristate
flabel metal3 s 79200 47712 80000 47824 0 FreeSans 448 0 0 0 la_data_out[40]
port 231 nsew signal tristate
flabel metal3 s 0 65856 800 65968 0 FreeSans 448 0 0 0 la_data_out[41]
port 232 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 la_data_out[42]
port 233 nsew signal tristate
flabel metal3 s 79200 26880 80000 26992 0 FreeSans 448 0 0 0 la_data_out[43]
port 234 nsew signal tristate
flabel metal3 s 79200 28224 80000 28336 0 FreeSans 448 0 0 0 la_data_out[44]
port 235 nsew signal tristate
flabel metal2 s 24192 79200 24304 80000 0 FreeSans 448 90 0 0 la_data_out[45]
port 236 nsew signal tristate
flabel metal2 s 52416 79200 52528 80000 0 FreeSans 448 90 0 0 la_data_out[46]
port 237 nsew signal tristate
flabel metal3 s 79200 41664 80000 41776 0 FreeSans 448 0 0 0 la_data_out[47]
port 238 nsew signal tristate
flabel metal2 s 45696 0 45808 800 0 FreeSans 448 90 0 0 la_data_out[48]
port 239 nsew signal tristate
flabel metal2 s 47040 0 47152 800 0 FreeSans 448 90 0 0 la_data_out[49]
port 240 nsew signal tristate
flabel metal3 s 79200 50400 80000 50512 0 FreeSans 448 0 0 0 la_data_out[4]
port 241 nsew signal tristate
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 la_data_out[50]
port 242 nsew signal tristate
flabel metal2 s 26208 79200 26320 80000 0 FreeSans 448 90 0 0 la_data_out[51]
port 243 nsew signal tristate
flabel metal2 s 44352 79200 44464 80000 0 FreeSans 448 90 0 0 la_data_out[52]
port 244 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 la_data_out[53]
port 245 nsew signal tristate
flabel metal3 s 79200 45024 80000 45136 0 FreeSans 448 0 0 0 la_data_out[54]
port 246 nsew signal tristate
flabel metal2 s 37632 79200 37744 80000 0 FreeSans 448 90 0 0 la_data_out[55]
port 247 nsew signal tristate
flabel metal3 s 0 57120 800 57232 0 FreeSans 448 0 0 0 la_data_out[56]
port 248 nsew signal tristate
flabel metal3 s 0 65184 800 65296 0 FreeSans 448 0 0 0 la_data_out[57]
port 249 nsew signal tristate
flabel metal2 s 43680 79200 43792 80000 0 FreeSans 448 90 0 0 la_data_out[58]
port 250 nsew signal tristate
flabel metal3 s 79200 42336 80000 42448 0 FreeSans 448 0 0 0 la_data_out[59]
port 251 nsew signal tristate
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 la_data_out[5]
port 252 nsew signal tristate
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 la_data_out[60]
port 253 nsew signal tristate
flabel metal2 s 57792 79200 57904 80000 0 FreeSans 448 90 0 0 la_data_out[61]
port 254 nsew signal tristate
flabel metal3 s 79200 28896 80000 29008 0 FreeSans 448 0 0 0 la_data_out[62]
port 255 nsew signal tristate
flabel metal2 s 34944 79200 35056 80000 0 FreeSans 448 90 0 0 la_data_out[63]
port 256 nsew signal tristate
flabel metal3 s 79200 31584 80000 31696 0 FreeSans 448 0 0 0 la_data_out[6]
port 257 nsew signal tristate
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 la_data_out[7]
port 258 nsew signal tristate
flabel metal3 s 79200 48384 80000 48496 0 FreeSans 448 0 0 0 la_data_out[8]
port 259 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 la_data_out[9]
port 260 nsew signal tristate
flabel metal3 s 79200 3360 80000 3472 0 FreeSans 448 0 0 0 la_oenb[0]
port 261 nsew signal input
flabel metal3 s 79200 73920 80000 74032 0 FreeSans 448 0 0 0 la_oenb[10]
port 262 nsew signal input
flabel metal3 s 79200 61152 80000 61264 0 FreeSans 448 0 0 0 la_oenb[11]
port 263 nsew signal input
flabel metal3 s 79200 16128 80000 16240 0 FreeSans 448 0 0 0 la_oenb[12]
port 264 nsew signal input
flabel metal3 s 79200 9408 80000 9520 0 FreeSans 448 0 0 0 la_oenb[13]
port 265 nsew signal input
flabel metal3 s 79200 63168 80000 63280 0 FreeSans 448 0 0 0 la_oenb[14]
port 266 nsew signal input
flabel metal3 s 79200 17472 80000 17584 0 FreeSans 448 0 0 0 la_oenb[15]
port 267 nsew signal input
flabel metal3 s 79200 10080 80000 10192 0 FreeSans 448 0 0 0 la_oenb[16]
port 268 nsew signal input
flabel metal3 s 79200 69216 80000 69328 0 FreeSans 448 0 0 0 la_oenb[17]
port 269 nsew signal input
flabel metal3 s 79200 12096 80000 12208 0 FreeSans 448 0 0 0 la_oenb[18]
port 270 nsew signal input
flabel metal3 s 79200 8064 80000 8176 0 FreeSans 448 0 0 0 la_oenb[19]
port 271 nsew signal input
flabel metal3 s 79200 6720 80000 6832 0 FreeSans 448 0 0 0 la_oenb[1]
port 272 nsew signal input
flabel metal3 s 79200 77952 80000 78064 0 FreeSans 448 0 0 0 la_oenb[20]
port 273 nsew signal input
flabel metal3 s 79200 14784 80000 14896 0 FreeSans 448 0 0 0 la_oenb[21]
port 274 nsew signal input
flabel metal3 s 79200 11424 80000 11536 0 FreeSans 448 0 0 0 la_oenb[22]
port 275 nsew signal input
flabel metal3 s 79200 7392 80000 7504 0 FreeSans 448 0 0 0 la_oenb[23]
port 276 nsew signal input
flabel metal3 s 79200 1344 80000 1456 0 FreeSans 448 0 0 0 la_oenb[24]
port 277 nsew signal input
flabel metal3 s 79200 75264 80000 75376 0 FreeSans 448 0 0 0 la_oenb[25]
port 278 nsew signal input
flabel metal3 s 79200 0 80000 112 0 FreeSans 448 0 0 0 la_oenb[26]
port 279 nsew signal input
flabel metal3 s 79200 79296 80000 79408 0 FreeSans 448 0 0 0 la_oenb[27]
port 280 nsew signal input
flabel metal3 s 79200 18144 80000 18256 0 FreeSans 448 0 0 0 la_oenb[28]
port 281 nsew signal input
flabel metal3 s 79200 5376 80000 5488 0 FreeSans 448 0 0 0 la_oenb[29]
port 282 nsew signal input
flabel metal3 s 79200 73248 80000 73360 0 FreeSans 448 0 0 0 la_oenb[2]
port 283 nsew signal input
flabel metal3 s 79200 19488 80000 19600 0 FreeSans 448 0 0 0 la_oenb[30]
port 284 nsew signal input
flabel metal3 s 79200 75936 80000 76048 0 FreeSans 448 0 0 0 la_oenb[31]
port 285 nsew signal input
flabel metal3 s 79200 2016 80000 2128 0 FreeSans 448 0 0 0 la_oenb[32]
port 286 nsew signal input
flabel metal3 s 79200 18816 80000 18928 0 FreeSans 448 0 0 0 la_oenb[33]
port 287 nsew signal input
flabel metal3 s 79200 6048 80000 6160 0 FreeSans 448 0 0 0 la_oenb[34]
port 288 nsew signal input
flabel metal3 s 79200 59808 80000 59920 0 FreeSans 448 0 0 0 la_oenb[35]
port 289 nsew signal input
flabel metal3 s 79200 77280 80000 77392 0 FreeSans 448 0 0 0 la_oenb[36]
port 290 nsew signal input
flabel metal3 s 79200 76608 80000 76720 0 FreeSans 448 0 0 0 la_oenb[37]
port 291 nsew signal input
flabel metal3 s 79200 72576 80000 72688 0 FreeSans 448 0 0 0 la_oenb[38]
port 292 nsew signal input
flabel metal3 s 79200 2688 80000 2800 0 FreeSans 448 0 0 0 la_oenb[39]
port 293 nsew signal input
flabel metal3 s 79200 65856 80000 65968 0 FreeSans 448 0 0 0 la_oenb[3]
port 294 nsew signal input
flabel metal3 s 79200 71904 80000 72016 0 FreeSans 448 0 0 0 la_oenb[40]
port 295 nsew signal input
flabel metal3 s 79200 66528 80000 66640 0 FreeSans 448 0 0 0 la_oenb[41]
port 296 nsew signal input
flabel metal3 s 79200 15456 80000 15568 0 FreeSans 448 0 0 0 la_oenb[42]
port 297 nsew signal input
flabel metal3 s 79200 61824 80000 61936 0 FreeSans 448 0 0 0 la_oenb[43]
port 298 nsew signal input
flabel metal3 s 79200 67872 80000 67984 0 FreeSans 448 0 0 0 la_oenb[44]
port 299 nsew signal input
flabel metal3 s 79200 78624 80000 78736 0 FreeSans 448 0 0 0 la_oenb[45]
port 300 nsew signal input
flabel metal3 s 79200 4032 80000 4144 0 FreeSans 448 0 0 0 la_oenb[46]
port 301 nsew signal input
flabel metal3 s 79200 63840 80000 63952 0 FreeSans 448 0 0 0 la_oenb[47]
port 302 nsew signal input
flabel metal3 s 79200 64512 80000 64624 0 FreeSans 448 0 0 0 la_oenb[48]
port 303 nsew signal input
flabel metal3 s 79200 10752 80000 10864 0 FreeSans 448 0 0 0 la_oenb[49]
port 304 nsew signal input
flabel metal3 s 79200 60480 80000 60592 0 FreeSans 448 0 0 0 la_oenb[4]
port 305 nsew signal input
flabel metal3 s 79200 70560 80000 70672 0 FreeSans 448 0 0 0 la_oenb[50]
port 306 nsew signal input
flabel metal3 s 79200 4704 80000 4816 0 FreeSans 448 0 0 0 la_oenb[51]
port 307 nsew signal input
flabel metal3 s 79200 16800 80000 16912 0 FreeSans 448 0 0 0 la_oenb[52]
port 308 nsew signal input
flabel metal3 s 79200 69888 80000 70000 0 FreeSans 448 0 0 0 la_oenb[53]
port 309 nsew signal input
flabel metal3 s 79200 62496 80000 62608 0 FreeSans 448 0 0 0 la_oenb[54]
port 310 nsew signal input
flabel metal3 s 79200 74592 80000 74704 0 FreeSans 448 0 0 0 la_oenb[55]
port 311 nsew signal input
flabel metal3 s 79200 12768 80000 12880 0 FreeSans 448 0 0 0 la_oenb[56]
port 312 nsew signal input
flabel metal3 s 79200 14112 80000 14224 0 FreeSans 448 0 0 0 la_oenb[57]
port 313 nsew signal input
flabel metal3 s 79200 59136 80000 59248 0 FreeSans 448 0 0 0 la_oenb[58]
port 314 nsew signal input
flabel metal3 s 79200 13440 80000 13552 0 FreeSans 448 0 0 0 la_oenb[59]
port 315 nsew signal input
flabel metal3 s 79200 68544 80000 68656 0 FreeSans 448 0 0 0 la_oenb[5]
port 316 nsew signal input
flabel metal3 s 79200 8736 80000 8848 0 FreeSans 448 0 0 0 la_oenb[60]
port 317 nsew signal input
flabel metal3 s 79200 71232 80000 71344 0 FreeSans 448 0 0 0 la_oenb[61]
port 318 nsew signal input
flabel metal3 s 79200 65184 80000 65296 0 FreeSans 448 0 0 0 la_oenb[62]
port 319 nsew signal input
flabel metal3 s 79200 672 80000 784 0 FreeSans 448 0 0 0 la_oenb[63]
port 320 nsew signal input
flabel metal3 s 79200 67200 80000 67312 0 FreeSans 448 0 0 0 la_oenb[6]
port 321 nsew signal input
flabel metal2 s 73248 79200 73360 80000 0 FreeSans 448 90 0 0 la_oenb[7]
port 322 nsew signal input
flabel metal2 s 73920 79200 74032 80000 0 FreeSans 448 90 0 0 la_oenb[8]
port 323 nsew signal input
flabel metal2 s 10080 79200 10192 80000 0 FreeSans 448 90 0 0 la_oenb[9]
port 324 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 out[0]
port 325 nsew signal input
flabel metal2 s 43008 79200 43120 80000 0 FreeSans 448 90 0 0 out[10]
port 326 nsew signal input
flabel metal3 s 0 53088 800 53200 0 FreeSans 448 0 0 0 out[11]
port 327 nsew signal input
flabel metal3 s 0 60480 800 60592 0 FreeSans 448 0 0 0 out[1]
port 328 nsew signal input
flabel metal2 s 53760 79200 53872 80000 0 FreeSans 448 90 0 0 out[2]
port 329 nsew signal input
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 out[3]
port 330 nsew signal input
flabel metal2 s 56448 79200 56560 80000 0 FreeSans 448 90 0 0 out[4]
port 331 nsew signal input
flabel metal2 s 50400 79200 50512 80000 0 FreeSans 448 90 0 0 out[5]
port 332 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 out[6]
port 333 nsew signal input
flabel metal2 s 23520 79200 23632 80000 0 FreeSans 448 90 0 0 out[7]
port 334 nsew signal input
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 out[8]
port 335 nsew signal input
flabel metal3 s 0 38304 800 38416 0 FreeSans 448 0 0 0 out[9]
port 336 nsew signal input
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 rst_n
port 337 nsew signal tristate
flabel metal2 s 33600 79200 33712 80000 0 FreeSans 448 90 0 0 sel[0]
port 338 nsew signal tristate
flabel metal2 s 51072 79200 51184 80000 0 FreeSans 448 90 0 0 sel[1]
port 339 nsew signal tristate
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 sel[2]
port 340 nsew signal tristate
flabel metal2 s 64512 79200 64624 80000 0 FreeSans 448 90 0 0 user_clock2
port 341 nsew signal input
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 user_irq[0]
port 342 nsew signal tristate
flabel metal3 s 0 66528 800 66640 0 FreeSans 448 0 0 0 user_irq[1]
port 343 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 user_irq[2]
port 344 nsew signal tristate
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 345 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 345 nsew power bidirectional
flabel metal4 s 65888 3076 66208 76892 0 FreeSans 1280 90 0 0 vdd
port 345 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 346 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 76892 0 FreeSans 1280 90 0 0 vss
port 346 nsew ground bidirectional
flabel metal2 s 47040 79200 47152 80000 0 FreeSans 448 90 0 0 wb_clk_i
port 347 nsew signal input
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 wb_rst_i
port 348 nsew signal input
flabel metal2 s 36288 79200 36400 80000 0 FreeSans 448 90 0 0 wbs_ack_o
port 349 nsew signal tristate
flabel metal2 s 72576 79200 72688 80000 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 350 nsew signal input
flabel metal2 s 14784 79200 14896 80000 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 351 nsew signal input
flabel metal2 s 16800 79200 16912 80000 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 352 nsew signal input
flabel metal2 s 8736 79200 8848 80000 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 353 nsew signal input
flabel metal2 s 67872 79200 67984 80000 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 354 nsew signal input
flabel metal2 s 12768 79200 12880 80000 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 355 nsew signal input
flabel metal2 s 59136 79200 59248 80000 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 356 nsew signal input
flabel metal2 s 61824 79200 61936 80000 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 357 nsew signal input
flabel metal2 s 79296 79200 79408 80000 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 358 nsew signal input
flabel metal2 s 1344 79200 1456 80000 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 359 nsew signal input
flabel metal2 s 76608 79200 76720 80000 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 360 nsew signal input
flabel metal2 s 60480 79200 60592 80000 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 361 nsew signal input
flabel metal2 s 63840 79200 63952 80000 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 362 nsew signal input
flabel metal2 s 65184 79200 65296 80000 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 363 nsew signal input
flabel metal2 s 66528 79200 66640 80000 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 364 nsew signal input
flabel metal2 s 65856 79200 65968 80000 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 365 nsew signal input
flabel metal2 s 18144 79200 18256 80000 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 366 nsew signal input
flabel metal2 s 78624 79200 78736 80000 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 367 nsew signal input
flabel metal2 s 59808 79200 59920 80000 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 368 nsew signal input
flabel metal2 s 63168 79200 63280 80000 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 369 nsew signal input
flabel metal2 s 62496 79200 62608 80000 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 370 nsew signal input
flabel metal2 s 74592 79200 74704 80000 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 371 nsew signal input
flabel metal2 s 61152 79200 61264 80000 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 372 nsew signal input
flabel metal2 s 21504 79200 21616 80000 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 373 nsew signal input
flabel metal2 s 75264 79200 75376 80000 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 374 nsew signal input
flabel metal2 s 67200 79200 67312 80000 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 375 nsew signal input
flabel metal2 s 18816 79200 18928 80000 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 376 nsew signal input
flabel metal2 s 77952 79200 78064 80000 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 377 nsew signal input
flabel metal2 s 77280 79200 77392 80000 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 378 nsew signal input
flabel metal2 s 71904 79200 72016 80000 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 379 nsew signal input
flabel metal2 s 4704 79200 4816 80000 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 380 nsew signal input
flabel metal2 s 70560 79200 70672 80000 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 381 nsew signal input
flabel metal2 s 3360 79200 3472 80000 0 FreeSans 448 90 0 0 wbs_cyc_i
port 382 nsew signal input
flabel metal2 s 20160 79200 20272 80000 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 383 nsew signal input
flabel metal2 s 2016 79200 2128 80000 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 384 nsew signal input
flabel metal2 s 672 79200 784 80000 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 385 nsew signal input
flabel metal2 s 68544 79200 68656 80000 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 386 nsew signal input
flabel metal2 s 7392 79200 7504 80000 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 387 nsew signal input
flabel metal2 s 2688 79200 2800 80000 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 388 nsew signal input
flabel metal2 s 10752 79200 10864 80000 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 389 nsew signal input
flabel metal2 s 4032 79200 4144 80000 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 390 nsew signal input
flabel metal2 s 17472 79200 17584 80000 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 391 nsew signal input
flabel metal2 s 8064 79200 8176 80000 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 392 nsew signal input
flabel metal2 s 14112 79200 14224 80000 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 393 nsew signal input
flabel metal2 s 13440 79200 13552 80000 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 394 nsew signal input
flabel metal2 s 9408 79200 9520 80000 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 395 nsew signal input
flabel metal2 s 11424 79200 11536 80000 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 396 nsew signal input
flabel metal2 s 0 79200 112 80000 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 397 nsew signal input
flabel metal2 s 75936 79200 76048 80000 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 398 nsew signal input
flabel metal2 s 16128 79200 16240 80000 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 399 nsew signal input
flabel metal2 s 15456 79200 15568 80000 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 400 nsew signal input
flabel metal2 s 6048 79200 6160 80000 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 401 nsew signal input
flabel metal2 s 5376 79200 5488 80000 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 402 nsew signal input
flabel metal2 s 71232 79200 71344 80000 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 403 nsew signal input
flabel metal2 s 12096 79200 12208 80000 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 404 nsew signal input
flabel metal2 s 6720 79200 6832 80000 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 405 nsew signal input
flabel metal2 s 20832 79200 20944 80000 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 406 nsew signal input
flabel metal2 s 19488 79200 19600 80000 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 407 nsew signal input
flabel metal2 s 69216 79200 69328 80000 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 408 nsew signal input
flabel metal2 s 69888 79200 70000 80000 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 409 nsew signal input
flabel metal3 s 0 79296 800 79408 0 FreeSans 448 0 0 0 wbs_dat_i[5]
port 410 nsew signal input
flabel metal3 s 0 78624 800 78736 0 FreeSans 448 0 0 0 wbs_dat_i[6]
port 411 nsew signal input
flabel metal3 s 0 77952 800 78064 0 FreeSans 448 0 0 0 wbs_dat_i[7]
port 412 nsew signal input
flabel metal3 s 0 77280 800 77392 0 FreeSans 448 0 0 0 wbs_dat_i[8]
port 413 nsew signal input
flabel metal3 s 0 76608 800 76720 0 FreeSans 448 0 0 0 wbs_dat_i[9]
port 414 nsew signal input
flabel metal3 s 0 55104 800 55216 0 FreeSans 448 0 0 0 wbs_dat_o[0]
port 415 nsew signal tristate
flabel metal3 s 0 57792 800 57904 0 FreeSans 448 0 0 0 wbs_dat_o[10]
port 416 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 wbs_dat_o[11]
port 417 nsew signal tristate
flabel metal3 s 0 58464 800 58576 0 FreeSans 448 0 0 0 wbs_dat_o[12]
port 418 nsew signal tristate
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 wbs_dat_o[13]
port 419 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 wbs_dat_o[14]
port 420 nsew signal tristate
flabel metal3 s 0 51744 800 51856 0 FreeSans 448 0 0 0 wbs_dat_o[15]
port 421 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 wbs_dat_o[16]
port 422 nsew signal tristate
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 wbs_dat_o[17]
port 423 nsew signal tristate
flabel metal3 s 0 59136 800 59248 0 FreeSans 448 0 0 0 wbs_dat_o[18]
port 424 nsew signal tristate
flabel metal3 s 0 37632 800 37744 0 FreeSans 448 0 0 0 wbs_dat_o[19]
port 425 nsew signal tristate
flabel metal3 s 0 51072 800 51184 0 FreeSans 448 0 0 0 wbs_dat_o[1]
port 426 nsew signal tristate
flabel metal3 s 0 50400 800 50512 0 FreeSans 448 0 0 0 wbs_dat_o[20]
port 427 nsew signal tristate
flabel metal3 s 0 63168 800 63280 0 FreeSans 448 0 0 0 wbs_dat_o[21]
port 428 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 wbs_dat_o[22]
port 429 nsew signal tristate
flabel metal3 s 0 47712 800 47824 0 FreeSans 448 0 0 0 wbs_dat_o[23]
port 430 nsew signal tristate
flabel metal3 s 0 48384 800 48496 0 FreeSans 448 0 0 0 wbs_dat_o[24]
port 431 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 wbs_dat_o[25]
port 432 nsew signal tristate
flabel metal3 s 0 52416 800 52528 0 FreeSans 448 0 0 0 wbs_dat_o[26]
port 433 nsew signal tristate
flabel metal3 s 0 40992 800 41104 0 FreeSans 448 0 0 0 wbs_dat_o[27]
port 434 nsew signal tristate
flabel metal3 s 0 46368 800 46480 0 FreeSans 448 0 0 0 wbs_dat_o[28]
port 435 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 wbs_dat_o[29]
port 436 nsew signal tristate
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 wbs_dat_o[2]
port 437 nsew signal tristate
flabel metal3 s 0 55776 800 55888 0 FreeSans 448 0 0 0 wbs_dat_o[30]
port 438 nsew signal tristate
flabel metal3 s 0 45696 800 45808 0 FreeSans 448 0 0 0 wbs_dat_o[31]
port 439 nsew signal tristate
flabel metal3 s 0 61152 800 61264 0 FreeSans 448 0 0 0 wbs_dat_o[3]
port 440 nsew signal tristate
flabel metal3 s 0 47040 800 47152 0 FreeSans 448 0 0 0 wbs_dat_o[4]
port 441 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 wbs_dat_o[5]
port 442 nsew signal tristate
flabel metal3 s 0 49056 800 49168 0 FreeSans 448 0 0 0 wbs_dat_o[6]
port 443 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 wbs_dat_o[7]
port 444 nsew signal tristate
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 wbs_dat_o[8]
port 445 nsew signal tristate
flabel metal3 s 0 49728 800 49840 0 FreeSans 448 0 0 0 wbs_dat_o[9]
port 446 nsew signal tristate
flabel metal3 s 0 75936 800 76048 0 FreeSans 448 0 0 0 wbs_sel_i[0]
port 447 nsew signal input
flabel metal3 s 0 75264 800 75376 0 FreeSans 448 0 0 0 wbs_sel_i[1]
port 448 nsew signal input
flabel metal3 s 0 74592 800 74704 0 FreeSans 448 0 0 0 wbs_sel_i[2]
port 449 nsew signal input
flabel metal3 s 0 73920 800 74032 0 FreeSans 448 0 0 0 wbs_sel_i[3]
port 450 nsew signal input
flabel metal3 s 0 73248 800 73360 0 FreeSans 448 0 0 0 wbs_stb_i
port 451 nsew signal input
flabel metal3 s 0 72576 800 72688 0 FreeSans 448 0 0 0 wbs_we_i
port 452 nsew signal input
rlabel metal1 39984 76048 39984 76048 0 vdd
rlabel metal1 39984 76832 39984 76832 0 vss
rlabel metal2 78232 59080 78232 59080 0 clk
rlabel metal3 78610 20216 78610 20216 0 in[0]
rlabel metal2 77896 57680 77896 57680 0 in[10]
rlabel metal3 1358 67256 1358 67256 0 in[11]
rlabel metal2 51800 2422 51800 2422 0 in[12]
rlabel metal2 22680 76608 22680 76608 0 in[13]
rlabel metal3 1358 12152 1358 12152 0 in[14]
rlabel metal2 50456 2198 50456 2198 0 in[15]
rlabel metal2 26936 2422 26936 2422 0 in[16]
rlabel metal2 58520 77938 58520 77938 0 in[17]
rlabel metal2 51800 77490 51800 77490 0 in[1]
rlabel metal2 42392 2198 42392 2198 0 in[2]
rlabel metal2 43064 1414 43064 1414 0 in[3]
rlabel metal2 78008 24752 78008 24752 0 in[4]
rlabel metal2 38360 77546 38360 77546 0 in[5]
rlabel metal2 40376 77546 40376 77546 0 in[6]
rlabel metal2 78008 21504 78008 21504 0 in[7]
rlabel metal3 1358 16856 1358 16856 0 in[8]
rlabel metal3 1638 29624 1638 29624 0 in[9]
rlabel metal3 41944 3528 41944 3528 0 io_in[10]
rlabel metal2 41160 3416 41160 3416 0 io_in[11]
rlabel metal2 78232 26600 78232 26600 0 io_in[12]
rlabel metal2 37128 76552 37128 76552 0 io_in[13]
rlabel metal2 36008 77000 36008 77000 0 io_in[14]
rlabel metal2 78232 20832 78232 20832 0 io_in[15]
rlabel metal3 1246 36344 1246 36344 0 io_in[16]
rlabel metal2 1736 32424 1736 32424 0 io_in[17]
rlabel metal2 78232 51240 78232 51240 0 io_in[18]
rlabel metal3 1246 64568 1246 64568 0 io_in[19]
rlabel metal2 43736 1022 43736 1022 0 io_in[20]
rlabel metal2 27496 76776 27496 76776 0 io_in[21]
rlabel metal2 1848 34608 1848 34608 0 io_in[22]
rlabel metal2 46760 3472 46760 3472 0 io_in[23]
rlabel metal2 27608 2142 27608 2142 0 io_in[24]
rlabel metal3 48104 76440 48104 76440 0 io_in[25]
rlabel metal2 28840 75768 28840 75768 0 io_in[5]
rlabel metal2 78232 56560 78232 56560 0 io_in[6]
rlabel metal2 28392 3416 28392 3416 0 io_in[7]
rlabel metal2 78232 33880 78232 33880 0 io_in[8]
rlabel metal2 55272 76944 55272 76944 0 io_in[9]
rlabel metal2 78008 30520 78008 30520 0 io_out[26]
rlabel metal3 1358 41720 1358 41720 0 io_out[27]
rlabel metal2 77896 54096 77896 54096 0 io_out[28]
rlabel metal3 1358 30968 1358 30968 0 io_out[29]
rlabel metal2 41048 77770 41048 77770 0 io_out[30]
rlabel metal2 77896 46760 77896 46760 0 io_out[31]
rlabel metal2 33656 2422 33656 2422 0 io_out[32]
rlabel metal2 27608 77770 27608 77770 0 io_out[33]
rlabel metal2 78008 25816 78008 25816 0 io_out[34]
rlabel metal3 78610 22904 78610 22904 0 io_out[35]
rlabel metal2 49784 77938 49784 77938 0 io_out[36]
rlabel metal3 1358 44408 1358 44408 0 io_out[37]
rlabel metal3 41496 35560 41496 35560 0 net1
rlabel metal2 2016 49672 2016 49672 0 net10
rlabel metal2 55160 77938 55160 77938 0 net100
rlabel metal3 1246 42392 1246 42392 0 net101
rlabel metal2 25704 76664 25704 76664 0 net102
rlabel metal2 23016 76664 23016 76664 0 net103
rlabel metal2 26992 76664 26992 76664 0 net104
rlabel metal2 30968 2030 30968 2030 0 net105
rlabel metal2 78232 33040 78232 33040 0 net106
rlabel metal2 46424 2030 46424 2030 0 net107
rlabel metal2 78232 46816 78232 46816 0 net108
rlabel metal2 47880 76664 47880 76664 0 net109
rlabel metal2 43008 3416 43008 3416 0 net11
rlabel metal3 1246 56504 1246 56504 0 net110
rlabel metal2 41832 75096 41832 75096 0 net111
rlabel metal3 77784 50400 77784 50400 0 net112
rlabel metal3 854 15512 854 15512 0 net113
rlabel metal3 78722 31640 78722 31640 0 net114
rlabel metal3 1246 33656 1246 33656 0 net115
rlabel metal3 78232 48608 78232 48608 0 net116
rlabel metal3 1246 22904 1246 22904 0 net117
rlabel metal2 77784 23632 77784 23632 0 net118
rlabel metal3 1246 53816 1246 53816 0 net119
rlabel metal2 27832 60312 27832 60312 0 net12
rlabel metal2 57288 76664 57288 76664 0 net120
rlabel metal2 78232 27776 78232 27776 0 net121
rlabel metal2 78288 29960 78288 29960 0 net122
rlabel metal2 39816 76664 39816 76664 0 net123
rlabel metal2 78232 54768 78232 54768 0 net124
rlabel metal2 49784 2030 49784 2030 0 net125
rlabel metal2 32312 2030 32312 2030 0 net126
rlabel metal2 47768 1190 47768 1190 0 net127
rlabel metal2 45192 76664 45192 76664 0 net128
rlabel metal3 1470 59864 1470 59864 0 net129
rlabel metal2 32648 36232 32648 36232 0 net13
rlabel metal2 29736 75544 29736 75544 0 net130
rlabel metal2 1736 12600 1736 12600 0 net131
rlabel metal2 49112 2030 49112 2030 0 net132
rlabel metal2 37688 2030 37688 2030 0 net133
rlabel metal3 78722 22232 78722 22232 0 net134
rlabel metal2 78232 34496 78232 34496 0 net135
rlabel metal3 1246 43064 1246 43064 0 net136
rlabel metal2 43456 75544 43456 75544 0 net137
rlabel metal3 1246 35000 1246 35000 0 net138
rlabel metal2 39032 2030 39032 2030 0 net139
rlabel metal2 46536 3864 46536 3864 0 net14
rlabel metal2 48440 2030 48440 2030 0 net140
rlabel metal2 35000 2030 35000 2030 0 net141
rlabel metal2 33096 76664 33096 76664 0 net142
rlabel metal2 36344 2030 36344 2030 0 net143
rlabel metal2 78232 51856 78232 51856 0 net144
rlabel metal2 45080 2590 45080 2590 0 net145
rlabel metal2 55944 75544 55944 75544 0 net146
rlabel metal2 37016 2030 37016 2030 0 net147
rlabel metal2 78232 48048 78232 48048 0 net148
rlabel metal3 1246 65912 1246 65912 0 net149
rlabel metal3 33376 3416 33376 3416 0 net15
rlabel metal2 35672 2030 35672 2030 0 net150
rlabel metal3 77560 26880 77560 26880 0 net151
rlabel metal2 78232 28336 78232 28336 0 net152
rlabel metal2 24136 76664 24136 76664 0 net153
rlabel metal2 52304 75544 52304 75544 0 net154
rlabel metal2 78232 41888 78232 41888 0 net155
rlabel metal2 45752 854 45752 854 0 net156
rlabel metal2 47096 1302 47096 1302 0 net157
rlabel metal2 34328 2030 34328 2030 0 net158
rlabel metal2 26376 76664 26376 76664 0 net159
rlabel metal2 44128 48440 44128 48440 0 net16
rlabel metal2 44744 77280 44744 77280 0 net160
rlabel metal2 1736 26880 1736 26880 0 net161
rlabel metal2 78232 45528 78232 45528 0 net162
rlabel metal2 37800 76664 37800 76664 0 net163
rlabel metal3 1246 57176 1246 57176 0 net164
rlabel metal3 1246 65240 1246 65240 0 net165
rlabel metal2 44296 76944 44296 76944 0 net166
rlabel metal2 78232 42448 78232 42448 0 net167
rlabel metal3 1246 14168 1246 14168 0 net168
rlabel metal2 57960 76664 57960 76664 0 net169
rlabel metal2 29512 61320 29512 61320 0 net17
rlabel metal2 78232 29232 78232 29232 0 net170
rlabel metal2 35112 76664 35112 76664 0 net171
rlabel metal3 1246 24920 1246 24920 0 net172
rlabel metal3 1246 66584 1246 66584 0 net173
rlabel metal3 1246 24248 1246 24248 0 net174
rlabel metal2 36680 77280 36680 77280 0 net175
rlabel metal3 1470 55160 1470 55160 0 net176
rlabel metal3 1246 51128 1246 51128 0 net177
rlabel metal3 854 43736 854 43736 0 net178
rlabel metal3 1246 61208 1246 61208 0 net179
rlabel metal3 45640 44072 45640 44072 0 net18
rlabel metal3 1246 47096 1246 47096 0 net180
rlabel metal3 1246 23576 1246 23576 0 net181
rlabel metal3 1246 49112 1246 49112 0 net182
rlabel metal3 1582 16184 1582 16184 0 net183
rlabel metal3 1582 35672 1582 35672 0 net184
rlabel metal3 1302 49784 1302 49784 0 net185
rlabel metal3 854 57848 854 57848 0 net186
rlabel metal3 1246 25592 1246 25592 0 net187
rlabel metal3 1246 58520 1246 58520 0 net188
rlabel metal3 1246 27608 1246 27608 0 net189
rlabel metal2 28840 3472 28840 3472 0 net19
rlabel metal3 1246 18872 1246 18872 0 net190
rlabel metal3 1246 51800 1246 51800 0 net191
rlabel metal3 1470 26264 1470 26264 0 net192
rlabel metal3 1246 14840 1246 14840 0 net193
rlabel metal3 1302 59192 1302 59192 0 net194
rlabel metal3 1246 37688 1246 37688 0 net195
rlabel metal2 2184 50400 2184 50400 0 net196
rlabel metal3 1246 63224 1246 63224 0 net197
rlabel metal3 1246 20216 1246 20216 0 net198
rlabel metal3 1246 47768 1246 47768 0 net199
rlabel metal2 41328 33096 41328 33096 0 net2
rlabel metal2 46648 34048 46648 34048 0 net20
rlabel metal3 1246 48440 1246 48440 0 net200
rlabel metal3 1246 18200 1246 18200 0 net201
rlabel metal3 1246 52472 1246 52472 0 net202
rlabel metal3 1246 41048 1246 41048 0 net203
rlabel metal3 1246 46424 1246 46424 0 net204
rlabel metal3 1582 20888 1582 20888 0 net205
rlabel metal3 1246 55832 1246 55832 0 net206
rlabel metal3 1470 45752 1470 45752 0 net207
rlabel metal2 34552 76440 34552 76440 0 net208
rlabel metal2 78232 52584 78232 52584 0 net209
rlabel metal2 55048 60368 55048 60368 0 net21
rlabel metal2 49224 76328 49224 76328 0 net210
rlabel metal2 31640 77770 31640 77770 0 net211
rlabel metal2 78232 57848 78232 57848 0 net212
rlabel metal2 78232 53480 78232 53480 0 net213
rlabel metal3 1582 30296 1582 30296 0 net214
rlabel metal2 28952 2198 28952 2198 0 net215
rlabel metal3 1246 32984 1246 32984 0 net216
rlabel metal2 39704 2198 39704 2198 0 net217
rlabel metal2 78232 35224 78232 35224 0 net218
rlabel metal2 78232 39368 78232 39368 0 net219
rlabel metal2 2072 16856 2072 16856 0 net22
rlabel metal2 30296 2198 30296 2198 0 net220
rlabel metal3 1246 13496 1246 13496 0 net221
rlabel metal2 31640 2198 31640 2198 0 net222
rlabel metal3 1246 28952 1246 28952 0 net223
rlabel metal3 78498 30968 78498 30968 0 net224
rlabel metal3 854 54488 854 54488 0 net225
rlabel metal2 77784 36120 77784 36120 0 net226
rlabel metal2 46536 76328 46536 76328 0 net227
rlabel metal3 1582 63896 1582 63896 0 net228
rlabel metal2 39088 76328 39088 76328 0 net229
rlabel metal2 43456 46872 43456 46872 0 net23
rlabel metal2 30408 75880 30408 75880 0 net230
rlabel metal2 78232 38472 78232 38472 0 net231
rlabel metal3 1246 39704 1246 39704 0 net232
rlabel metal2 29624 2198 29624 2198 0 net233
rlabel metal2 2408 48832 2408 48832 0 net24
rlabel metal2 2632 48188 2632 48188 0 net25
rlabel metal3 50064 41944 50064 41944 0 net26
rlabel metal3 18032 31080 18032 31080 0 net27
rlabel metal3 41776 45080 41776 45080 0 net28
rlabel metal3 48272 45304 48272 45304 0 net29
rlabel metal2 77896 26992 77896 26992 0 net3
rlabel metal3 18312 20104 18312 20104 0 net30
rlabel metal2 24920 71876 24920 71876 0 net31
rlabel metal2 43736 38024 43736 38024 0 net32
rlabel metal2 40040 39144 40040 39144 0 net33
rlabel metal3 17864 21672 17864 21672 0 net34
rlabel metal2 77784 59080 77784 59080 0 net35
rlabel metal2 46088 26936 46088 26936 0 net36
rlabel metal2 75096 49084 75096 49084 0 net37
rlabel metal2 4536 67816 4536 67816 0 net38
rlabel metal2 51856 4312 51856 4312 0 net39
rlabel metal2 38248 41944 38248 41944 0 net4
rlabel metal2 25256 75656 25256 75656 0 net40
rlabel metal2 4312 12824 4312 12824 0 net41
rlabel metal2 50904 3864 50904 3864 0 net42
rlabel metal2 29624 4256 29624 4256 0 net43
rlabel metal3 50960 48104 50960 48104 0 net44
rlabel metal2 51632 75656 51632 75656 0 net45
rlabel metal2 43736 4368 43736 4368 0 net46
rlabel via2 42504 5096 42504 5096 0 net47
rlabel metal2 75768 24640 75768 24640 0 net48
rlabel metal2 39816 74816 39816 74816 0 net49
rlabel metal3 37968 48440 37968 48440 0 net5
rlabel metal2 40320 74760 40320 74760 0 net50
rlabel metal2 75488 21560 75488 21560 0 net51
rlabel metal2 4312 17528 4312 17528 0 net52
rlabel metal2 4312 30072 4312 30072 0 net53
rlabel metal2 75656 30912 75656 30912 0 net54
rlabel metal2 4312 41888 4312 41888 0 net55
rlabel metal2 75376 54376 75376 54376 0 net56
rlabel metal3 4592 31752 4592 31752 0 net57
rlabel metal3 42280 74760 42280 74760 0 net58
rlabel metal2 45192 45752 45192 45752 0 net59
rlabel metal3 59416 20552 59416 20552 0 net6
rlabel metal2 36008 5544 36008 5544 0 net60
rlabel metal2 30856 76720 30856 76720 0 net61
rlabel metal2 75656 26208 75656 26208 0 net62
rlabel metal2 75768 23072 75768 23072 0 net63
rlabel metal2 51240 76384 51240 76384 0 net64
rlabel metal3 4592 45080 4592 45080 0 net65
rlabel metal3 4592 22344 4592 22344 0 net66
rlabel metal2 36456 75208 36456 75208 0 net67
rlabel metal3 48160 44408 48160 44408 0 net68
rlabel metal3 4592 28616 4592 28616 0 net69
rlabel metal2 2072 36736 2072 36736 0 net7
rlabel metal3 78722 41048 78722 41048 0 net70
rlabel metal2 78232 32480 78232 32480 0 net71
rlabel metal2 53144 78218 53144 78218 0 net72
rlabel metal2 25200 76664 25200 76664 0 net73
rlabel metal3 78498 45752 78498 45752 0 net74
rlabel metal2 32984 2030 32984 2030 0 net75
rlabel metal2 78232 24024 78232 24024 0 net76
rlabel metal2 78288 44072 78288 44072 0 net77
rlabel metal3 78722 43064 78722 43064 0 net78
rlabel metal2 32424 76664 32424 76664 0 net79
rlabel metal2 34944 38696 34944 38696 0 net8
rlabel metal2 31080 75544 31080 75544 0 net80
rlabel metal3 1246 61880 1246 61880 0 net81
rlabel metal2 78232 37184 78232 37184 0 net82
rlabel metal2 78232 37744 78232 37744 0 net83
rlabel metal2 77784 40656 77784 40656 0 net84
rlabel metal2 78232 56000 78232 56000 0 net85
rlabel metal3 78498 55160 78498 55160 0 net86
rlabel metal2 78232 44800 78232 44800 0 net87
rlabel metal2 51128 2030 51128 2030 0 net88
rlabel metal2 78288 50344 78288 50344 0 net89
rlabel metal2 77784 47544 77784 47544 0 net9
rlabel metal2 45864 76664 45864 76664 0 net90
rlabel metal2 78232 40208 78232 40208 0 net91
rlabel metal3 1470 40376 1470 40376 0 net92
rlabel metal3 1246 45080 1246 45080 0 net93
rlabel metal3 1246 62552 1246 62552 0 net94
rlabel metal2 78232 49504 78232 49504 0 net95
rlabel metal2 40376 2030 40376 2030 0 net96
rlabel metal3 1246 39032 1246 39032 0 net97
rlabel metal2 38360 2030 38360 2030 0 net98
rlabel metal3 78722 36344 78722 36344 0 net99
rlabel metal2 1736 17304 1736 17304 0 out[0]
rlabel metal2 43848 76720 43848 76720 0 out[10]
rlabel metal2 1848 53424 1848 53424 0 out[11]
rlabel metal2 1736 60648 1736 60648 0 out[1]
rlabel metal2 54488 76832 54488 76832 0 out[2]
rlabel metal2 1736 31360 1736 31360 0 out[3]
rlabel metal2 57064 76832 57064 76832 0 out[4]
rlabel metal2 50512 76440 50512 76440 0 out[5]
rlabel metal2 1736 19768 1736 19768 0 out[6]
rlabel metal3 23240 76440 23240 76440 0 out[7]
rlabel metal2 1736 37128 1736 37128 0 out[8]
rlabel metal2 1736 38584 1736 38584 0 out[9]
rlabel metal3 1358 21560 1358 21560 0 rst_n
rlabel metal2 34104 76608 34104 76608 0 sel[0]
rlabel metal2 51128 77154 51128 77154 0 sel[1]
rlabel metal3 1358 28280 1358 28280 0 sel[2]
rlabel metal2 46536 46760 46536 46760 0 wb_clk_i
rlabel metal2 1736 22008 1736 22008 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>
