* NGSPICE file created from totp.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

.subckt totp clk in[0] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18]
+ in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] out[0] out[10] out[11] out[1]
+ out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] rst_n vdd vss
X_3155_ hotp.block.mixer.msg\[127\] hotp.block.mixer.msg\[128\] _1330_ _1331_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2106_ _0555_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3086_ _1291_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2037_ _0514_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold522_I hotp.block.sha1.mixer.w\[427\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3988_ net465 clknet_leaf_114_clk hotp.block.sha1.mixer.w\[215\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2939_ _1207_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold351 stream.key_buf\[21\] net371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold362 hotp.block.sha1.mixer.b\[3\] net382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold340 hotp.block.sha1.mixer.e\[4\] net360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold395 stream.key_buf\[139\] net415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold373 hotp.block.sha1.mixer.w\[319\] net393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold384 hotp.block.sha1.mixer.d\[1\] net404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3911_ net596 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[138\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3842_ net368 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[69\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3773_ net300 clknet_leaf_96_clk hotp.block.debug\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2724_ _1030_ _1055_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold103_I hotp.block.sha1.mixer.w\[461\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2655_ hotp.digest\[17\] _0993_ _0994_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2586_ hotp.digest\[9\] _0932_ _0933_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4325_ _0226_ clknet_leaf_89_clk hotp.block.mixer.msg\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold472_I hotp.block.sha1.mixer.w\[184\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3272__C _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4256_ net454 clknet_leaf_99_clk hotp.block.sha1.mixer.w\[483\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3207_ hotp.block.mixer.msg\[150\] hotp.block.mixer.msg\[151\] _1356_ _1360_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4187_ net331 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[414\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3138_ hotp.block.mixer.msg\[120\] hotp.block.mixer.msg\[121\] _1319_ _1321_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3069_ _1281_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold170 stream.key_buf\[59\] net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2858__I _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold181 hotp.block.sha1.mixer.w\[12\] net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold192 hotp.block.sha1.mixer.w\[432\] net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__1711__B _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ _0610_ _0632_ _0613_ _0798_ _0752_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_75_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2371_ _1421_ _0643_ _0741_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4110_ net277 clknet_leaf_19_clk hotp.block.sha1.mixer.w\[337\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4041_ net174 clknet_leaf_14_clk hotp.block.sha1.mixer.w\[268\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold220_I hotp.block.sha1.mixer.w\[379\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold318_I hotp.block.sha1.mixer.w\[458\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3825_ net151 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3756_ net500 clknet_leaf_81_clk hotp.block.sha1.mixer.e\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2707_ hotp.digest\[23\] _1040_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3687_ net761 clknet_leaf_82_clk hotp.block.sha1.mixer.c\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2638_ _0840_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2569_ _0918_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4308_ _0209_ clknet_leaf_105_clk hotp.block.mixer.msg\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2932__I1 hotp.block.mixer.msg\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3940__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4239_ net573 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[466\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1648__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1940_ hotp.block.sha1.mixer.c\[30\] _0421_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1871_ _1521_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3610_ _0183_ clknet_leaf_45_clk hotp.digest\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4190__D net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3541_ _0118_ clknet_leaf_17_clk stream.digest\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3472_ net572 clknet_leaf_32_clk stream.key_buf\[124\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_23_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2423_ stream.counter\[8\] _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2354_ _0729_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2285_ _0689_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_84_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4024_ net764 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[251\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_32_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_hold435_I hotp.block.sha1.mixer.w\[128\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_99_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold602_I hotp.block.sha1.mixer.w\[365\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3493__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_22_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3808_ net769 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3739_ net737 clknet_leaf_86_clk hotp.block.sha1.mixer.d\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_37_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3836__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2070_ _0529_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4185__D net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2972_ _1226_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1923_ _0407_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1854_ _1508_ _1504_ _1531_ _1607_ _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_53_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1785_ hotp.block.magic.step\[0\] _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold703 hotp.block.sha1.mixer.c\[25\] net723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold725 stream.key_buf\[14\] net745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold736 hotp.block.sha1.mixer.w\[272\] net756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3524_ _0101_ clknet_leaf_15_clk stream.digest\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold714 hotp.block.sha1.mixer.w\[18\] net734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3455_ net607 clknet_leaf_34_clk stream.key_buf\[107\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold747 hotp.block.sha1.mixer.e\[12\] net767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold758 hotp.block.sha1.mixer.d\[5\] net778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold769 hotp.block.sha1.mixer.d\[26\] net789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2406_ _1426_ _0769_ _0771_ _0746_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_hold385_I hotp.block.sha1.mixer.w\[251\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4141__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3386_ net517 clknet_leaf_54_clk stream.key_buf\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2337_ stream.digest\[22\] stream.digest\[23\] _0717_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2268_ _1439_ _0650_ _0634_ _0509_ _1448_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_46_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2276__A1 hotp.block.main_in vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4007_ net530 clknet_leaf_1_clk hotp.block.sha1.mixer.w\[234\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2199_ _0602_ _0603_ _0609_ _0612_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold30 hotp.block.sha1.mixer.w\[295\] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold41 hotp.block.sha1.mixer.w\[337\] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1770__I _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold74 stream.key_buf\[135\] net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold63 stream.key_buf\[147\] net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold52 hotp.block.sha1.mixer.w\[460\] net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold96 hotp.block.sha1.mixer.w\[335\] net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold85 hotp.block.sha1.mixer.w\[96\] net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_58_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_5 net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3240_ _1380_ _1381_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3171_ _1339_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3812__D net595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2122_ _0564_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2053_ _0525_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ _1216_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1906_ stream.ready _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2886_ _1177_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_20_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1837_ seg.digit\[3\] _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold511 hotp.block.sha1.mixer.w\[311\] net531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_96_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold500 hotp.block.sha1.mixer.w\[227\] net520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold533 hotp.block.sha1.mixer.w\[104\] net553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3507_ _0013_ clknet_leaf_42_clk stream.key_buf\[159\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold522 hotp.block.sha1.mixer.w\[427\] net542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold544 hotp.block.sha1.mixer.w\[469\] net564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1768_ _1510_ _1528_ _1512_ _1529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1699_ _1422_ _1464_ _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold588 hotp.block.sha1.mixer.w\[245\] net608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold555 hotp.block.sha1.mixer.w\[499\] net575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold566 hotp.block.sha1.mixer.w\[5\] net586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold577 hotp.block.sha1.mixer.e\[3\] net597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3438_ net82 clknet_leaf_35_clk stream.key_buf\[90\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold767_I hotp.block.sha1.mixer.w\[147\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold599 hotp.block.sha1.mixer.w\[59\] net619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3369_ net814 clknet_leaf_55_clk stream.key_buf\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4187__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_114_clk clknet_4_0_0_clk clknet_leaf_114_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 net20 out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_52_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3404__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2740_ hotp.digest\[30\] _1068_ _1069_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_105_clk clknet_4_2_0_clk clknet_leaf_105_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2671_ _0365_ _0429_ _1008_ hotp.digest\[22\] _0846_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_5_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4410_ _0311_ clknet_leaf_62_clk hotp.block.mixer.msg\[122\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3807__D net584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4341_ _0242_ clknet_leaf_86_clk hotp.block.mixer.msg\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4272_ net92 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[499\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3223_ hotp.block.mixer.msg\[157\] hotp.block.mixer.msg\[158\] _1366_ _1369_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3154_ _1329_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2105_ stream.msg_buf\[28\] stream.msg_buf\[29\] _0551_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3085_ hotp.block.mixer.msg\[97\] hotp.block.mixer.msg\[98\] _1288_ _1291_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_6_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2036_ _1439_ _1463_ _0513_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_hold348_I hotp.block.sha1.mixer.w\[70\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold515_I hotp.block.sha1.mixer.w\[167\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3987_ net397 clknet_leaf_114_clk hotp.block.sha1.mixer.w\[214\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2938_ hotp.block.mixer.msg\[34\] hotp.block.mixer.msg\[35\] _1203_ _1207_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2869_ hotp.block.mixer.msg\[4\] hotp.block.mixer.msg\[5\] _1166_ _1168_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold330 hotp.block.sha1.mixer.w\[353\] net350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold341 hotp.block.sha1.mixer.w\[430\] net361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold352 hotp.block.sha1.mixer.w\[15\] net372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold396 hotp.block.sha1.mixer.w\[133\] net416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold374 hotp.block.sha1.mixer.w\[407\] net394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold385 hotp.block.sha1.mixer.w\[251\] net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold363 hotp.block.sha1.mixer.a\[29\] net383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_5_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4202__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4193__D net797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3910_ net507 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[137\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3841_ net547 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[68\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3772_ hotp.block.sha1.mixer.d\[0\] clknet_leaf_85_clk hotp.block.sha1.mixer.e\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2723_ hotp.digest\[25\] _1053_ _1054_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2654_ _0975_ _0978_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_30_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2585_ _0918_ _0920_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4324_ _0225_ clknet_leaf_90_clk hotp.block.mixer.msg\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4255_ net700 clknet_leaf_99_clk hotp.block.sha1.mixer.w\[482\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold465_I hotp.block.sha1.mixer.w\[99\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3206_ _1359_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4186_ net77 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[413\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3137_ _1320_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3068_ hotp.block.mixer.msg\[90\] hotp.block.mixer.msg\[91\] _1277_ _1281_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2019_ hotp.block.sha1.mixer.a_carry\[0\] _1590_ _0497_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_9_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2140__S _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold171 hotp.block.sha1.mixer.w\[508\] net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold160 hotp.block.sha1.mixer.w\[240\] net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold182 stream.key_buf\[13\] net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold193 hotp.block.sha1.mixer.w\[418\] net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3910__D net507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_87_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2370_ _1463_ _0740_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4040_ net614 clknet_leaf_14_clk hotp.block.sha1.mixer.w\[267\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_96_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3824_ net260 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3755_ net661 clknet_leaf_81_clk hotp.block.sha1.mixer.e\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2706_ _0901_ _1039_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3686_ net444 clknet_leaf_82_clk hotp.block.sha1.mixer.c\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2637_ hotp.digest\[15\] _0978_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2568_ hotp.digest\[7\] hotp.digest\[8\] hotp.digest\[9\] _0918_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2499_ _0856_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4307_ _0208_ clknet_leaf_105_clk hotp.block.mixer.msg\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2895__S _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ net803 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[465\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1648__A2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4169_ net48 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[396\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_94_clk clknet_4_9_0_clk clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_85_clk clknet_4_8_0_clk clknet_leaf_85_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_61_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1870_ _1618_ _1605_ _1628_ _1524_ _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_12_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3540_ _0117_ clknet_leaf_14_clk stream.digest\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3471_ net722 clknet_leaf_32_clk stream.key_buf\[123\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2422_ _0646_ _0785_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2353_ stream.digest\[29\] stream.digest\[30\] _0727_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2284_ _0688_ _0625_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4023_ net405 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[250\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_88_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_76_clk clknet_4_11_0_clk clknet_leaf_76_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold428_I hotp.block.sha1.mixer.w\[234\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1858__I _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3638__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3807_ net584 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1999_ _0383_ _0466_ _0477_ _1575_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3738_ net721 clknet_leaf_86_clk hotp.block.sha1.mixer.d\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3669_ net552 clknet_leaf_93_clk hotp.block.sha1.mixer.b\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_67_clk clknet_4_12_0_clk clknet_leaf_67_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output12_I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2599__I _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold37_I hotp.block.sha1.mixer.w\[456\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_58_clk clknet_4_14_0_clk clknet_leaf_58_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4093__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2971_ hotp.block.mixer.msg\[48\] hotp.block.mixer.msg\[49\] _1224_ _1226_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1922_ _0406_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1853_ _1610_ _1588_ _1611_ _1612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1784_ hotp.block.magic.step\[1\] _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold737 stream.key_buf\[68\] net757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold704 stream.key_buf\[159\] net724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3523_ _0100_ clknet_leaf_15_clk stream.digest\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold726 hotp.block.sha1.mixer.w\[202\] net746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold715 hotp.block.sha1.mixer.w\[387\] net735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3454_ net428 clknet_leaf_34_clk stream.key_buf\[106\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold759 hotp.block.sha1.mixer.w\[280\] net779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold748 hotp.block.sha1.mixer.w\[239\] net768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2405_ _0676_ _0745_ _0770_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3385_ net687 clknet_leaf_54_clk stream.key_buf\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2336_ _0719_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_49_clk clknet_4_13_0_clk clknet_leaf_49_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2267_ _0672_ _0674_ _0662_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4006_ net448 clknet_leaf_1_clk hotp.block.sha1.mixer.w\[233\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2198_ _0610_ _0611_ stream.counter\[8\] _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_95_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold31 stream.key_buf\[54\] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold20 hotp.block.sha1.mixer.b\[1\] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold64 stream.key_buf\[103\] net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold53 hotp.block.sha1.mixer.w\[140\] net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold42 hotp.block.sha1.mixer.d\[10\] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold97 stream.key_buf\[11\] net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold75 hotp.block.sha1.mixer.w\[358\] net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold86 hotp.block.sha1.mixer.w\[29\] net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_109_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_83_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_6 net499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_98_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3170_ hotp.block.mixer.msg\[134\] hotp.block.mixer.msg\[135\] _1335_ _1339_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2121_ stream.msg_buf\[35\] stream.msg_buf\[36\] _0561_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_21_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2993__S _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__D net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2052_ stream.msg_buf\[5\] stream.msg_buf\[6\] _0524_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_36_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2954_ hotp.block.mixer.msg\[41\] hotp.block.mixer.msg\[42\] _1213_ _1216_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1905_ _1490_ _0393_ _0395_ _1489_ net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_2885_ hotp.block.mixer.msg\[11\] hotp.block.mixer.msg\[12\] _1176_ _1177_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1836_ seg.digit\[3\] _1487_ _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold501 hotp.block.sha1.mixer.w\[320\] net521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1767_ _1511_ _1528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold512 stream.key_buf\[90\] net532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold523 hotp.block.sha1.mixer.w\[137\] net543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold545 stream.key_buf\[153\] net565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3506_ net724 clknet_leaf_42_clk stream.key_buf\[158\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold534 hotp.block.sha1.mixer.w\[217\] net554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1698_ _1427_ _1445_ _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold556 hotp.block.sha1.mixer.w\[287\] net576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold567 hotp.block.sha1.mixer.w\[116\] net587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_60_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold578 hotp.block.sha1.mixer.w\[81\] net598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__2967__I _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3437_ net532 clknet_leaf_35_clk stream.key_buf\[89\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold589 hotp.block.sha1.mixer.w\[203\] net609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_109_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3368_ net371 clknet_leaf_55_clk stream.key_buf\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2319_ _0709_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3299_ _0040_ clknet_leaf_40_clk stream.msg_buf\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput10 net10 out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3913__D net407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1999__A1 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4131__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2670_ _1007_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_35_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3849__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4340_ _0241_ clknet_leaf_86_clk hotp.block.mixer.msg\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4271_ net575 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[498\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3222_ _1368_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input3_I in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3153_ _1159_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2104_ _0554_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3084_ _1290_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2035_ _0512_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold243_I hotp.block.sha1.mixer.w\[83\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_hold410_I hotp.block.sha1.mixer.w\[205\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3986_ net411 clknet_leaf_114_clk hotp.block.sha1.mixer.w\[213\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold508_I hotp.block.sha1.mixer.w\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2937_ _1206_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2868_ _1167_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_107_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold320 stream.key_buf\[132\] net340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2799_ _0807_ _1110_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1819_ _1495_ _1532_ _1579_ _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_5_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold331 stream.key_buf\[63\] net351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold353 hotp.block.sha1.mixer.w\[343\] net373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold342 hotp.block.sha1.mixer.w\[420\] net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold386 stream.key_buf\[72\] net406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold375 hotp.block.sha1.mixer.w\[17\] net395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold364 hotp.block.sha1.mixer.b\[21\] net384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold397 hotp.block.sha1.mixer.w\[233\] net417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_5_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_116_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_107_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2138__S _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3840_ net621 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[67\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3771_ net765 clknet_leaf_85_clk hotp.block.sha1.mixer.e\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2722_ _1037_ _1040_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_70_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3671__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2653_ _0992_ _0978_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_93_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2584_ _0931_ _0920_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4027__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4323_ _0224_ clknet_leaf_90_clk hotp.block.mixer.msg\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold193_I hotp.block.sha1.mixer.w\[418\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4254_ net292 clknet_leaf_96_clk hotp.block.sha1.mixer.w\[481\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3205_ hotp.block.mixer.msg\[149\] hotp.block.mixer.msg\[150\] _1356_ _1359_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4177__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4185_ net30 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[412\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold458_I hotp.block.sha1.mixer.w\[105\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3136_ hotp.block.mixer.msg\[119\] hotp.block.mixer.msg\[120\] _1319_ _1320_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3067_ _1280_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2018_ _1559_ _0479_ _0488_ _0496_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XTAP_TAPCELL_ROW_102_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3969_ net238 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[196\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold161 hotp.block.sha1.mixer.w\[112\] net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold150 hotp.block.sha1.mixer.w\[271\] net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold183 hotp.block.sha1.mixer.w\[208\] net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_0_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold172 hotp.block.sha1.mixer.w\[176\] net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold194 hotp.block.sha1.mixer.w\[26\] net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_69_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2606__A2 _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3823_ net445 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_15_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3754_ net791 clknet_leaf_81_clk hotp.block.sha1.mixer.e\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _1617_ _1036_ _1037_ _1038_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3685_ net810 clknet_leaf_82_clk hotp.block.sha1.mixer.c\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2636_ _0901_ _0977_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2567_ _1617_ _0378_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2498_ _0855_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold575_I hotp.block.sha1.mixer.w\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4306_ _0207_ clknet_leaf_105_clk hotp.block.mixer.msg\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4237_ net339 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[464\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold742_I hotp.block.sha1.mixer.w\[373\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ net327 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[395\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4099_ net80 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[326\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3119_ _1310_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3921__D net766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3470_ net175 clknet_leaf_33_clk stream.key_buf\[122\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4199__D net542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2421_ _0677_ _0776_ _0780_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2352_ _0728_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2283_ _0633_ _0687_ _0688_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4022_ net355 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[249\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_88_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4215__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold156_I hotp.block.sha1.mixer.w\[391\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold323_I hotp.block.sha1.mixer.w\[376\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3806_ net646 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1998_ _0449_ _0461_ _1620_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3737_ net216 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_99_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3668_ net27 clknet_leaf_69_clk hotp.block.sha1.mixer.b\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2619_ hotp.digest\[13\] _0961_ _0962_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3599_ _0172_ clknet_leaf_46_clk stream.key_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_110_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3732__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3916__D net499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3882__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2357__I1 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4238__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2970_ _1225_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1921_ _1418_ _1419_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1852_ _1515_ _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1783_ _1541_ _1542_ _1543_ _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold716 stream.key_buf\[41\] net736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold727 hotp.block.sha1.mixer.w\[143\] net747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3522_ _0099_ clknet_leaf_15_clk stream.digest\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold705 hotp.block.sha1.mixer.b\[27\] net725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3453_ net413 clknet_leaf_34_clk stream.key_buf\[105\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold749 hotp.block.sha1.mixer.w\[36\] net769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold738 hotp.block.sha1.mixer.b\[18\] net758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2404_ _0739_ _0767_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3384_ net248 clknet_leaf_55_clk stream.key_buf\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2335_ stream.digest\[21\] stream.digest\[22\] _0717_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2266_ _0657_ _0673_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold273_I hotp.block.sha1.mixer.w\[90\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2197_ stream.counter\[9\] _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4005_ net417 clknet_leaf_1_clk hotp.block.sha1.mixer.w\[232\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold538_I hotp.block.sha1.mixer.w\[266\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1787__A2 _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold21 hotp.block.sha1.mixer.w\[259\] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold32 hotp.block.sha1.mixer.w\[270\] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold10 hotp.block.sha1.mixer.w\[413\] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold54 stream.key_buf\[109\] net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold65 hotp.block.sha1.mixer.w\[502\] net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold43 hotp.block.sha1.mixer.c\[29\] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold87 stream.key_buf\[104\] net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold98 stream.key_buf\[7\] net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold76 hotp.block.sha1.mixer.d\[11\] net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2019__A3 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__A2 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3646__D net816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_7 net696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2120_ _0563_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2051_ _0516_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_107_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2953_ _1215_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1904_ _1581_ _1582_ _1597_ _0394_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_17_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2884_ _1161_ _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_44_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1835_ _1589_ _1578_ _1594_ _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_96_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1766_ _1517_ _1518_ _1522_ _1526_ _1527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xhold502 hotp.block.sha1.mixer.w\[180\] net522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold524 stream.key_buf\[64\] net544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3505_ net344 clknet_leaf_42_clk stream.key_buf\[157\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold513 hotp.block.sha1.mixer.w\[249\] net533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold535 hotp.block.sha1.mixer.w\[229\] net555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold579 hotp.block.sha1.mixer.w\[360\] net599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1697_ _1451_ _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold557 hotp.block.sha1.mixer.w\[497\] net577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_hold390_I hotp.block.sha1.mixer.w\[179\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold546 hotp.block.sha1.mixer.a\[25\] net566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold568 hotp.block.sha1.mixer.w\[503\] net588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3436_ net550 clknet_leaf_35_clk stream.key_buf\[88\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3367_ net187 clknet_leaf_49_clk stream.key_buf\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2318_ stream.digest\[14\] stream.digest\[15\] _0706_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3298_ _0039_ clknet_leaf_40_clk stream.msg_buf\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2249_ stream.digest\[0\] stream.digest\[4\] stream.digest\[8\] stream.digest\[12\]
+ _0658_ _0659_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_0_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xoutput11 net11 out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 net9 out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_32_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2893__I _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3920__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4270_ net112 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[497\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3221_ hotp.block.mixer.msg\[156\] hotp.block.mixer.msg\[157\] _1366_ _1368_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3152_ _1328_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4000__D net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2103_ stream.msg_buf\[27\] stream.msg_buf\[28\] _0551_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3083_ hotp.block.mixer.msg\[96\] hotp.block.mixer.msg\[97\] _1288_ _1290_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2034_ _1452_ _0507_ _0511_ _0406_ _1441_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_9_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3985_ net537 clknet_leaf_114_clk hotp.block.sha1.mixer.w\[212\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2936_ hotp.block.mixer.msg\[33\] hotp.block.mixer.msg\[34\] _1203_ _1206_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold403_I hotp.block.sha1.mixer.w\[153\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2867_ hotp.block.mixer.msg\[3\] hotp.block.mixer.msg\[4\] _1166_ _1167_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1818_ _1495_ _1578_ _1579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2798_ _1113_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold310 hotp.block.sha1.mixer.w\[55\] net330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold332 hotp.block.sha1.mixer.w\[117\] net352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold321 hotp.block.sha1.mixer.w\[178\] net341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1749_ hotp.block.mixer.round\[5\] _1510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold343 hotp.block.sha1.mixer.w\[257\] net363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold387 hotp.block.sha1.mixer.w\[141\] net407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold376 hotp.block.sha1.mixer.e\[2\] net396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold354 hotp.block.sha1.mixer.w\[219\] net374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold365 hotp.block.sha1.mixer.w\[485\] net385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold398 stream.key_buf\[92\] net418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3419_ net406 clknet_leaf_52_clk stream.key_buf\[71\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4399_ _0300_ clknet_leaf_61_clk hotp.block.mixer.msg\[111\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_82_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_97_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_62_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_20_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3924__D net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_35_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold12_I hotp.block.sha1.mixer.w\[82\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_108_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3770_ net128 clknet_leaf_84_clk hotp.block.sha1.mixer.e\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2721_ _1052_ _1040_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2652_ _0959_ _0968_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2583_ _0897_ _0908_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3834__D net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4322_ _0223_ clknet_leaf_90_clk hotp.block.mixer.msg\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4253_ _0011_ clknet_leaf_99_clk hotp.block.sha1.mixer.w\[480\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3204_ _1358_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4184_ net526 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[411\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold186_I hotp.block.sha1.mixer.w\[65\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3135_ _1308_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3066_ hotp.block.mixer.msg\[89\] hotp.block.mixer.msg\[90\] _1277_ _1280_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2017_ _1536_ _0491_ _0495_ _1559_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3968_ net739 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[195\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2919_ hotp.block.mixer.msg\[26\] hotp.block.mixer.msg\[27\] _1192_ _1196_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3899_ net697 clknet_leaf_25_clk hotp.block.sha1.mixer.w\[126\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold151 stream.key_buf\[120\] net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold162 hotp.block.sha1.mixer.w\[434\] net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold140 hotp.block.sha1.mixer.c\[1\] net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold184 hotp.block.sha1.mixer.w\[350\] net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold173 hotp.block.sha1.mixer.w\[345\] net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold195 hotp.block.sha1.mixer.w\[392\] net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3839__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3919__D net787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3822_ net288 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_15_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3753_ net281 clknet_leaf_80_clk hotp.block.sha1.mixer.e\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2704_ hotp.digest\[26\] _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3684_ net122 clknet_leaf_84_clk hotp.block.sha1.mixer.c\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2635_ _1617_ _0974_ _0975_ _0976_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2566_ _0380_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_10_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4305_ _0206_ clknet_leaf_105_clk hotp.block.mixer.msg\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2497_ _0837_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4236_ net290 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[463\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4167_ net560 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[394\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3118_ hotp.block.mixer.msg\[111\] hotp.block.mixer.msg\[112\] _1309_ _1310_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4098_ net398 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[325\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3049_ _1270_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2342__S _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2420_ _0781_ _0783_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2351_ stream.digest\[28\] stream.digest\[29\] _0727_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2282_ _1424_ _0406_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4021_ net533 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[248\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_88_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold149_I hotp.block.sha1.mixer.w\[443\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1997_ _1621_ _0473_ _0474_ _0475_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3805_ net632 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold316_I hotp.block.sha1.mixer.w\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3736_ net196 clknet_leaf_86_clk hotp.block.sha1.mixer.d\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3667_ net665 clknet_leaf_93_clk hotp.block.sha1.mixer.b\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3598_ _0171_ clknet_leaf_47_clk stream.key_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2618_ _0901_ _0917_ _0947_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2549_ _0846_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2986__I _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4219_ net322 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[446\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3932__D net641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2337__S _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1920_ _1490_ _1593_ _0405_ net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1851_ hotp.block.mixer.stage\[1\] _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1782_ hotp.block.magic.step\[2\] _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3521_ _0098_ clknet_leaf_15_clk stream.digest\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold706 stream.key_buf\[40\] net726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_52_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold728 hotp.block.sha1.mixer.w\[209\] net748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4003__D net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold717 hotp.block.sha1.mixer.d\[31\] net737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3452_ net610 clknet_leaf_34_clk stream.key_buf\[104\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold739 hotp.block.sha1.mixer.w\[110\] net759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3383_ net224 clknet_leaf_54_clk stream.key_buf\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2403_ _0509_ _0609_ _0736_ _0768_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3842__D net368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2334_ _0718_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2265_ stream.digest\[3\] stream.digest\[7\] stream.digest\[11\] stream.digest\[15\]
+ _0658_ _0659_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_34_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2196_ stream.counter\[10\] _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4004_ net613 clknet_leaf_1_clk hotp.block.sha1.mixer.w\[231\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold600_I hotp.block.sha1.mixer.w\[150\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3719_ net96 clknet_leaf_83_clk hotp.block.sha1.mixer.d\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold22 hotp.block.sha1.mixer.w\[278\] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold11 hotp.block.sha1.mixer.w\[84\] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold44 stream.key_buf\[157\] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold33 hotp.block.sha1.mixer.w\[282\] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold55 hotp.block.sha1.mixer.w\[510\] net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold66 stream.key_buf\[141\] net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold77 hotp.block.sha1.mixer.w\[309\] net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold99 hotp.block.sha1.mixer.w\[428\] net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold88 hotp.block.sha1.mixer.w\[370\] net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_79_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1795__I _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3927__D net475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4205__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2050_ _0523_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2952_ hotp.block.mixer.msg\[40\] hotp.block.mixer.msg\[41\] _1213_ _1215_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_108_clk clknet_4_2_0_clk clknet_leaf_108_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1903_ _1479_ _1481_ _1601_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_84_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2883_ _1175_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3837__D net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1834_ _1589_ _1593_ _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1765_ hotp.block.mixer.msg\[32\] _1525_ _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold536 stream.key_buf\[137\] net556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3504_ net64 clknet_leaf_20_clk stream.key_buf\[156\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold503 hotp.block.sha1.mixer.d\[25\] net523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold525 hotp.block.sha1.mixer.w\[195\] net545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold514 hotp.block.sha1.mixer.w\[419\] net534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3435_ net728 clknet_leaf_35_clk stream.key_buf\[87\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold558 hotp.block.sha1.mixer.w\[317\] net578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1696_ _1461_ _1462_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold569 hotp.block.sha1.mixer.w\[56\] net589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold547 hotp.block.sha1.mixer.e\[21\] net567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3366_ net262 clknet_leaf_54_clk stream.key_buf\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3297_ _0038_ clknet_leaf_40_clk stream.msg_buf\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2317_ _0708_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2248_ net5 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_hold648_I hotp.block.sha1.mixer.w\[173\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2179_ _0596_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold815_I hotp.block.sha1.mixer.w\[375\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3872__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput12 net12 out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_9_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3220_ _1367_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3151_ hotp.block.mixer.msg\[126\] hotp.block.mixer.msg\[127\] _1324_ _1328_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2102_ _0553_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3082_ _1289_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2033_ _1444_ _0510_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3984_ net688 clknet_leaf_114_clk hotp.block.sha1.mixer.w\[211\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold229_I hotp.block.sha1.mixer.w\[241\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2935_ _1205_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2866_ _1161_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1817_ _1544_ _1548_ _1577_ _1578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xhold300 stream.key_buf\[8\] net320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2797_ _0814_ _0807_ _1109_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold311 hotp.block.sha1.mixer.w\[415\] net331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_102_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold333 hotp.block.sha1.mixer.w\[325\] net353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold344 hotp.block.sha1.mixer.w\[285\] net364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1748_ _1497_ _1508_ _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold322 hotp.block.sha1.mixer.e\[1\] net342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold366 stream.key_buf\[17\] net386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1679_ _1420_ _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_68_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold377 hotp.block.sha1.mixer.w\[215\] net397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold355 hotp.block.sha1.mixer.a\[20\] net375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3418_ net470 clknet_leaf_52_clk stream.key_buf\[70\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold399 hotp.block.sha1.mixer.w\[318\] net419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4398_ _0299_ clknet_leaf_58_clk hotp.block.mixer.msg\[110\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold765_I hotp.block.sha1.mixer.w\[221\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold388 hotp.block.sha1.mixer.w\[476\] net408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3349_ net391 clknet_leaf_47_clk stream.key_buf\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3940__D net830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2720_ _1019_ _1029_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2651_ _0850_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1983__I _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2582_ hotp.digest\[11\] _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4321_ _0222_ clknet_leaf_90_clk hotp.block.mixer.msg\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4011__D net768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4252_ net811 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[479\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3203_ hotp.block.mixer.msg\[148\] hotp.block.mixer.msg\[149\] _1356_ _1358_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4183_ net695 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[410\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3850__D net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3134_ _1318_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_66_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3065_ _1279_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2016_ _0492_ _0493_ _0494_ _1554_ hotp.block.magic.step\[2\] _0495_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_49_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold513_I hotp.block.sha1.mixer.w\[249\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3967_ net545 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[194\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2918_ _1195_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_30_clk clknet_4_5_0_clk clknet_leaf_30_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_75_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3898_ net655 clknet_leaf_25_clk hotp.block.sha1.mixer.w\[125\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3910__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2849_ _1152_ _1153_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold130 stream.key_buf\[129\] net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold152 hotp.block.sha1.mixer.w\[457\] net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold141 hotp.block.sha1.mixer.w\[231\] net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold174 hotp.block.sha1.mixer.w\[331\] net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold163 hotp.block.sha1.mixer.a\[13\] net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold185 hotp.block.sha1.mixer.w\[390\] net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold196 hotp.block.sha1.mixer.d\[29\] net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_97_clk clknet_4_9_0_clk clknet_leaf_97_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_21_clk clknet_4_4_0_clk clknet_leaf_21_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3935__D net829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_88_clk clknet_4_8_0_clk clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4096__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3264__A1 _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1814__A2 _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3821_ net156 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4006__D net448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3933__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3752_ net767 clknet_leaf_80_clk hotp.block.sha1.mixer.e\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_clk clknet_4_1_0_clk clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2703_ hotp.digest\[23\] hotp.digest\[24\] hotp.digest\[25\] _1037_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3683_ net298 clknet_leaf_81_clk hotp.block.sha1.mixer.c\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3845__D net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2634_ hotp.digest\[18\] _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_81_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2565_ _0841_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4304_ _0205_ clknet_leaf_103_clk hotp.block.mixer.msg\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2496_ hotp.digest\[1\] _0842_ _0849_ _0853_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_10_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_96_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4235_ net104 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[462\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_79_clk clknet_4_10_0_clk clknet_leaf_79_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4166_ net743 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[393\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3117_ _1308_ _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4097_ net353 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[324\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3048_ hotp.block.mixer.msg\[81\] hotp.block.mixer.msg\[82\] _1267_ _1270_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold728_I hotp.block.sha1.mixer.w\[209\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_49_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_92_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_107_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold72_I hotp.block.sha1.mixer.w\[500\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_6_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1980__A1 _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2350_ _0711_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2281_ _0685_ _0686_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_1_clk clknet_4_0_0_clk clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4020_ net252 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[247\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_88_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3804_ net488 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1996_ _0458_ _0452_ _0454_ _1620_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3735_ net279 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3666_ net66 clknet_leaf_78_clk hotp.block.sha1.mixer.b\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4261__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3597_ _0170_ clknet_leaf_49_clk stream.key_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2617_ _0960_ _0948_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_hold580_I hotp.block.sha1.mixer.w\[446\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3829__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2548_ _0899_ _0887_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_hold678_I hotp.block.sha1.mixer.w\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3163__I _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2479_ hotp.rst_n _0821_ _0832_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4218_ net600 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[445\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4149_ net593 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[376\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2242__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4134__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2353__S _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1850_ _1532_ _1607_ _1608_ _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1781_ _1507_ _1501_ _1502_ _1530_ _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_4_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3520_ _0097_ clknet_leaf_15_clk stream.digest\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold718 hotp.block.sha1.mixer.w\[100\] net738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold707 hotp.block.sha1.mixer.w\[393\] net727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3451_ net107 clknet_leaf_31_clk stream.key_buf\[103\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold729 hotp.block.sha1.mixer.w\[400\] net749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3382_ net562 clknet_leaf_54_clk stream.key_buf\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2402_ _0613_ _0767_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2333_ stream.digest\[20\] stream.digest\[21\] _0717_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2264_ _0652_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2195_ stream.counter\[7\] _0605_ _0399_ _0608_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4003_ net161 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[230\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold426_I hotp.block.sha1.mixer.w\[171\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ _1546_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3718_ net62 clknet_leaf_86_clk hotp.block.sha1.mixer.d\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1944__A1 hotp.block.sha1.mixer.w\[64\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3649_ net210 clknet_leaf_80_clk hotp.block.sha1.mixer.b\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold23 hotp.block.sha1.mixer.w\[386\] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold12 hotp.block.sha1.mixer.w\[82\] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__2011__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold56 stream.key_buf\[111\] net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold34 hotp.block.sha1.mixer.w\[330\] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold45 hotp.block.sha1.mixer.e\[29\] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold89 hotp.block.sha1.mixer.w\[46\] net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold78 hotp.block.sha1.mixer.c\[17\] net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold67 hotp.block.sha1.mixer.c\[2\] net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output10_I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2901__S _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3943__D net446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2348__S _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2951_ _1214_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1902_ _1578_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3674__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2882_ hotp.block.mixer.msg\[10\] hotp.block.mixer.msg\[11\] _1171_ _1175_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1833_ _1592_ _1593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4014__D net711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1764_ _1509_ _1524_ _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3503_ net804 clknet_leaf_20_clk stream.key_buf\[155\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold526 hotp.block.sha1.mixer.w\[289\] net546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold515 hotp.block.sha1.mixer.w\[167\] net535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold504 hotp.block.sha1.mixer.w\[41\] net524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3853__D net598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3434_ net514 clknet_leaf_35_clk stream.key_buf\[86\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold548 hotp.block.sha1.mixer.w\[125\] net568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1695_ _1405_ _1422_ _1404_ _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold559 hotp.block.sha1.mixer.e\[19\] net579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold537 hotp.block.sha1.mixer.w\[7\] net557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3365_ net251 clknet_leaf_49_clk stream.key_buf\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3296_ _0037_ clknet_leaf_38_clk stream.msg_buf\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2316_ stream.digest\[13\] stream.digest\[14\] _0706_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2247_ net4 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2178_ stream.msg_buf\[60\] stream.msg_buf\[61\] _0592_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold808_I hotp.block.sha1.mixer.w\[334\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_14_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2006__B _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput13 net13 out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold5_I hotp.block.sha1.mixer.w\[410\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_67_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__D net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1908__A1 _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_91_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3150_ _1327_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2101_ stream.msg_buf\[26\] stream.msg_buf\[27\] _0551_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3081_ hotp.block.mixer.msg\[95\] hotp.block.mixer.msg\[96\] _1288_ _1289_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2032_ _1415_ _0509_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4009__D net527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3983_ net179 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[210\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3848__D net635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold124_I hotp.block.sha1.mixer.w\[384\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2934_ hotp.block.mixer.msg\[32\] hotp.block.mixer.msg\[33\] _1203_ _1205_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2865_ _1165_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1816_ _1561_ _1567_ _1570_ _1564_ _1576_ _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2796_ _1112_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold301 hotp.block.sha1.mixer.w\[61\] net321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold312 hotp.block.sha1.mixer.w\[368\] net332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold334 hotp.block.sha1.mixer.w\[369\] net354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold323 hotp.block.sha1.mixer.w\[376\] net343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1747_ _1507_ _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold378 hotp.block.sha1.mixer.w\[326\] net398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold367 hotp.block.sha1.mixer.w\[134\] net387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1678_ _1434_ _1446_ _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold345 hotp.block.sha1.mixer.w\[357\] net365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold356 hotp.block.sha1.mixer.a\[26\] net376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3417_ net751 clknet_leaf_52_clk stream.key_buf\[69\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4397_ _0298_ clknet_leaf_58_clk hotp.block.mixer.msg\[109\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold389 hotp.block.sha1.mixer.w\[188\] net409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3348_ net335 clknet_leaf_47_clk stream.key_buf\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3279_ _0020_ clknet_leaf_50_clk stream.msg_buf\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_107_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_103_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2650_ hotp.digest\[19\] _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3712__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2003__B1 _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_112_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_93_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2581_ _0914_ _0928_ _0929_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4320_ _0221_ clknet_leaf_92_clk hotp.block.mixer.msg\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4251_ net357 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[478\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3202_ _1357_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4182_ net25 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[409\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3133_ hotp.block.mixer.msg\[118\] hotp.block.mixer.msg\[119\] _1314_ _1318_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3064_ hotp.block.mixer.msg\[88\] hotp.block.mixer.msg\[89\] _1277_ _1279_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4218__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2015_ _1556_ _0470_ _0453_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_93_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2490__B1 _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3966_ net424 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[193\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold506_I hotp.block.sha1.mixer.w\[412\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2917_ hotp.block.mixer.msg\[25\] hotp.block.mixer.msg\[26\] _1192_ _1195_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3897_ net568 clknet_leaf_25_clk hotp.block.sha1.mixer.w\[124\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3392__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2848_ hotp.block.sha1.mixer.a_carry\[1\] _1142_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2779_ _1467_ _1456_ _0640_ _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4202__D net361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold131 hotp.block.sha1.mixer.w\[53\] net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold120 hotp.block.sha1.mixer.w\[422\] net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold153 hotp.block.sha1.mixer.c\[21\] net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold142 hotp.block.sha1.mixer.a\[2\] net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold175 stream.key_buf\[45\] net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold164 stream.key_buf\[116\] net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4449_ _0349_ clknet_leaf_68_clk hotp.block.mixer.round\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold186 hotp.block.sha1.mixer.w\[65\] net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold197 hotp.block.sha1.mixer.c\[5\] net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_8_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3735__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2784__A1 _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3951__D net410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_2_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3820_ net153 clknet_leaf_105_clk hotp.block.sha1.mixer.w\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_15_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3751_ net833 clknet_leaf_80_clk hotp.block.sha1.mixer.e\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2702_ _0374_ _0429_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3682_ net135 clknet_leaf_79_clk hotp.block.sha1.mixer.c\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2633_ hotp.digest\[15\] hotp.digest\[16\] hotp.digest\[17\] _0975_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2564_ _0883_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4022__D net355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4303_ _0204_ clknet_leaf_104_clk hotp.block.mixer.msg\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2495_ _0851_ _0852_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3861__D net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4234_ net69 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[461\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4165_ net727 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[392\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3116_ _1244_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4096_ net753 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[323\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3047_ _1269_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1805__A3 _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2766__A1 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3949_ net137 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[176\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2904__S _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3946__D net626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold65_I hotp.block.sha1.mixer.w\[502\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1980__A2 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2280_ _0676_ _1439_ _1416_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__D net608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3803_ net460 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3856__D net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1995_ _1574_ _0449_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3734_ net789 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3665_ net384 clknet_leaf_78_clk hotp.block.sha1.mixer.b\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2616_ _0930_ _0939_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1971__A2 hotp.block.sha1.mixer.c\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3596_ _0169_ clknet_leaf_50_clk stream.key_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2547_ _0867_ _0878_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2478_ _0816_ _0835_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_hold573_I hotp.block.sha1.mixer.w\[377\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4217_ net633 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[444\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold740_I hotp.block.sha1.mixer.w\[98\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4148_ net343 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[375\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4079_ net88 clknet_leaf_33_clk hotp.block.sha1.mixer.w\[306\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3923__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_80_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_95_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__D hotp.block.debug\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1780_ _1535_ _1540_ _1541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold708 stream.key_buf\[88\] net728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold719 hotp.block.sha1.mixer.w\[196\] net739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3450_ net84 clknet_leaf_35_clk stream.key_buf\[102\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3381_ net650 clknet_leaf_54_clk stream.key_buf\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2401_ _0400_ _0608_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2332_ _0711_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_33_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2263_ stream.digest\[19\] stream.digest\[23\] stream.digest\[27\] stream.digest\[31\]
+ _0653_ _0654_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4002_ net501 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[229\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2194_ stream.counter\[4\] _0607_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_48_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold321_I hotp.block.sha1.mixer.w\[178\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_106_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3717_ net259 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1978_ _0437_ _0451_ _0456_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1944__A2 hotp.block.sha1.mixer.w\[256\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold788_I hotp.block.sha1.mixer.w\[470\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3648_ net235 clknet_leaf_79_clk hotp.block.sha1.mixer.b\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3579_ _0152_ clknet_leaf_62_clk hotp.digest\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4210__D net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold13 hotp.block.sha1.mixer.a\[18\] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold35 stream.key_buf\[74\] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_4_10_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold24 hotp.block.sha1.mixer.b\[16\] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold46 hotp.block.sha1.mixer.b\[22\] net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold68 hotp.block.sha1.mixer.w\[307\] net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold57 hotp.block.sha1.mixer.w\[414\] net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold79 hotp.block.sha1.mixer.c\[27\] net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1880__B2 _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold28_I hotp.block.sha1.mixer.w\[397\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4101__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2950_ hotp.block.mixer.msg\[39\] hotp.block.mixer.msg\[40\] _1213_ _1214_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1901_ _1490_ _0390_ _0392_ _1489_ net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_8_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2881_ _1174_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1832_ _1590_ _1591_ _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1763_ _1523_ _1503_ _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3502_ net590 clknet_leaf_20_clk stream.key_buf\[154\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1694_ _1404_ _1449_ _1460_ _1410_ _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold527 hotp.block.sha1.mixer.w\[69\] net547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold516 hotp.block.sha1.mixer.w\[20\] net536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold505 hotp.block.sha1.mixer.w\[423\] net525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3433_ net689 clknet_leaf_35_clk stream.key_buf\[85\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold549 hotp.block.sha1.mixer.w\[336\] net569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold538 hotp.block.sha1.mixer.w\[266\] net558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4030__D net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3364_ net386 clknet_leaf_49_clk stream.key_buf\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3295_ _0036_ clknet_leaf_38_clk stream.msg_buf\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2315_ _0707_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2246_ net6 _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2177_ _0595_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_49_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_105_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4205__D net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput14 net14 out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2248__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4274__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3954__D net302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_78_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2100_ _0552_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3080_ _1287_ _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_27_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2031_ _1414_ _0508_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3641__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3982_ net601 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[209\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2933_ _1204_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4025__D net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2864_ hotp.block.mixer.msg\[2\] hotp.block.mixer.msg\[3\] _1162_ _1165_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2795_ _0809_ _0814_ _1110_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1815_ _1563_ _1549_ _1571_ _1573_ _1575_ _1576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_53_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold117_I hotp.block.sha1.mixer.w\[177\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3864__D net696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold302 hotp.block.sha1.mixer.w\[447\] net322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1746_ hotp.block.mixer.round\[1\] _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold313 stream.key_buf\[152\] net333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold324 stream.key_buf\[158\] net344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold335 hotp.block.sha1.mixer.w\[250\] net355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold357 stream.key_buf\[50\] net377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold368 hotp.block.sha1.mixer.w\[300\] net388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1677_ _1441_ _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold346 hotp.block.sha1.mixer.w\[263\] net366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_7_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3416_ net462 clknet_leaf_52_clk stream.key_buf\[68\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold379 hotp.block.sha1.mixer.w\[115\] net399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4396_ _0297_ clknet_leaf_58_clk hotp.block.mixer.msg\[108\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold486_I hotp.block.sha1.mixer.w\[374\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3347_ _0084_ clknet_leaf_16_clk seg.digit\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_51_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3278_ _0019_ clknet_leaf_39_clk stream.msg_buf\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_107_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2229_ _0642_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2012__B2 _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3949__D net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2003__A1 _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2580_ hotp.digest\[9\] _0906_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2003__B2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4250_ net752 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[477\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3201_ hotp.block.mixer.msg\[147\] hotp.block.mixer.msg\[148\] _1356_ _1357_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4181_ net574 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[408\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3132_ _1317_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3063_ _1278_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2014_ _0382_ _0463_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_89_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3859__D net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2490__B2 _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3965_ net149 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[192\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3896_ net692 clknet_leaf_25_clk hotp.block.sha1.mixer.w\[123\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2916_ _1194_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2847_ hotp.block.sha1.mixer.a_carry\[2\] _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2778_ _1098_ _1095_ _1099_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold110 hotp.block.sha1.mixer.w\[451\] net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold143 stream.key_buf\[97\] net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold132 hotp.block.sha1.mixer.w\[152\] net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_14_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold121 hotp.block.sha1.mixer.w\[225\] net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1729_ hotp.block.debug\[1\] _1491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold154 hotp.block.sha1.mixer.w\[269\] net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold165 hotp.block.sha1.mixer.w\[166\] net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold176 hotp.block.sha1.mixer.d\[28\] net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4448_ hotp.block.sha1.mixer.w_fb clknet_leaf_97_clk hotp.block.sha1.mixer.t vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold187 stream.key_buf\[55\] net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold198 hotp.block.sha1.mixer.a\[1\] net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4379_ _0280_ clknet_leaf_73_clk hotp.block.mixer.msg\[91\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1808__A1 hotp.block.magic.step\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold10_I hotp.block.sha1.mixer.w\[413\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3750_ net670 clknet_leaf_80_clk hotp.block.sha1.mixer.e\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2701_ _1005_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3681_ net217 clknet_leaf_84_clk hotp.block.sha1.mixer.c\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2632_ _0376_ _0374_ _0369_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2563_ _0884_ _0912_ _0913_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4302_ _0203_ clknet_leaf_104_clk hotp.block.mixer.msg\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2494_ hotp.digest\[39\] _0848_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4233_ net123 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[460\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4164_ net215 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[391\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4095_ net425 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[322\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3115_ _1307_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3046_ hotp.block.mixer.msg\[80\] hotp.block.mixer.msg\[81\] _1267_ _1269_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4335__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3948_ net192 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[175\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4213__D net718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3879_ net93 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[106\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_115_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4208__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3962__D net836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3802_ net318 clknet_leaf_107_clk hotp.block.sha1.mixer.w\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ _1574_ _0454_ _0443_ _0472_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3733_ net523 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_7_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3664_ net704 clknet_leaf_78_clk hotp.block.sha1.mixer.b\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2615_ hotp.digest\[15\] _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1971__A3 _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3595_ _0168_ clknet_leaf_50_clk stream.key_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3872__D net738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2546_ _0859_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2477_ _0364_ _0814_ _0807_ _1499_ _0834_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_110_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4216_ net316 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[443\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4147_ net835 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[374\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4078_ net476 clknet_leaf_33_clk hotp.block.sha1.mixer.w\[305\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4208__D net435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3029_ hotp.block.mixer.msg\[73\] hotp.block.mixer.msg\[74\] _1256_ _1259_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3875__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2009__C hotp.block.magic.step\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2739__A2 _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3957__D net549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold709 hotp.block.sha1.mixer.b\[19\] net729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _0764_ _0766_ _0759_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3380_ stream.key_buf\[33\] clknet_leaf_56_clk stream.key_buf\[32\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2331_ _0716_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2262_ _0668_ _0670_ _0662_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4001_ net555 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[228\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2193_ stream.counter\[3\] stream.counter\[2\] _0606_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4028__D net834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3867__D net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3716_ net167 clknet_leaf_86_clk hotp.block.sha1.mixer.d\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ _0453_ _0455_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3647_ net382 clknet_leaf_79_clk hotp.block.sha1.mixer.b\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3578_ _0151_ clknet_leaf_63_clk hotp.digest\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2529_ _0855_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_54_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold14 hotp.block.sha1.mixer.b\[14\] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold47 hotp.block.sha1.mixer.w\[501\] net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold25 hotp.block.sha1.mixer.d\[3\] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold36 hotp.block.sha1.mixer.w\[471\] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold58 hotp.block.sha1.mixer.w\[328\] net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold69 stream.key_buf\[149\] net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3190__I _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2409__A1 _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1900_ _1581_ _0391_ _1492_ _1597_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2880_ hotp.block.mixer.msg\[9\] hotp.block.mixer.msg\[10\] _1171_ _1174_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1831_ hotp.block.sha1.mixer.h_carry _1580_ _1591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_41_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1762_ _1500_ _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3501_ net684 clknet_leaf_20_clk stream.key_buf\[153\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1693_ _1402_ _1446_ _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold517 hotp.block.sha1.mixer.w\[213\] net537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold506 hotp.block.sha1.mixer.w\[412\] net526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3432_ net693 clknet_leaf_35_clk stream.key_buf\[84\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold528 hotp.block.sha1.mixer.w\[79\] net548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold539 hotp.block.sha1.mixer.w\[67\] net559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3363_ net790 clknet_leaf_49_clk stream.key_buf\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3294_ _0035_ clknet_leaf_38_clk stream.msg_buf\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2314_ stream.digest\[12\] stream.digest\[13\] _0706_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2245_ _0652_ _0655_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2176_ stream.msg_buf\[59\] stream.msg_buf\[60\] _0592_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold264_I hotp.block.sha1.mixer.w\[72\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold431_I hotp.block.sha1.mixer.w\[94\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold529_I hotp.block.sha1.mixer.w\[185\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60_clk clknet_4_14_0_clk clknet_leaf_60_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput15 net15 out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__4221__D net583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_94_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1853__A2 _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_51_clk clknet_4_13_0_clk clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_32_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_47_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4131__D net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold40_I hotp.block.sha1.mixer.w\[474\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3970__D net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4099__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2030_ stream.state\[1\] _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_105_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3981_ net748 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[208\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3936__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2932_ hotp.block.mixer.msg\[31\] hotp.block.mixer.msg\[32\] _1203_ _1204_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_42_clk clknet_4_6_0_clk clknet_leaf_42_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2863_ _1164_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2794_ _1111_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1814_ hotp.block.magic.step\[1\] _1574_ _1575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1745_ _1505_ _1506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold314 stream.key_buf\[83\] net334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold325 hotp.block.sha1.mixer.w\[340\] net345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold303 hotp.block.sha1.mixer.w\[206\] net323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold347 hotp.block.sha1.mixer.w\[288\] net367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold358 hotp.block.sha1.mixer.w\[351\] net378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1676_ _1444_ _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold336 hotp.block.sha1.mixer.e\[18\] net356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_22_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold369 hotp.block.sha1.mixer.b\[11\] net389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3415_ net757 clknet_leaf_52_clk stream.key_buf\[67\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4395_ _0296_ clknet_leaf_59_clk hotp.block.mixer.msg\[107\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3880__D net706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold479_I hotp.block.sha1.mixer.w\[144\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold381_I hotp.block.sha1.mixer.w\[362\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3346_ _0083_ clknet_leaf_98_clk seg.digit\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3277_ _0018_ clknet_leaf_39_clk stream.msg_buf\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_107_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2228_ stream.key_state\[0\] stream.msg_state\[0\] _1419_ _0641_ _0642_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2159_ _0585_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1835__A2 _1578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4216__D net316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33_clk clknet_4_5_0_clk clknet_leaf_33_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2012__A2 _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4241__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1771__B2 _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_24_clk clknet_4_4_0_clk clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_17_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold88_I hotp.block.sha1.mixer.w\[370\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3965__D net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_26_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4180_ net603 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[407\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3200_ _1350_ _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3131_ hotp.block.mixer.msg\[117\] hotp.block.mixer.msg\[118\] _1314_ _1317_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3062_ hotp.block.mixer.msg\[87\] hotp.block.mixer.msg\[88\] _1277_ _1278_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1817__A2 _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2013_ _1556_ _0444_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_35_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_102_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_15_clk clknet_4_3_0_clk clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3964_ net242 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[191\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3895_ net777 clknet_leaf_25_clk hotp.block.sha1.mixer.w\[122\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3875__D net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2915_ hotp.block.mixer.msg\[24\] hotp.block.mixer.msg\[25\] _1192_ _1194_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2846_ _0502_ _1146_ _1150_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2777_ stream.key_counter\[4\] _0638_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold100 hotp.block.sha1.mixer.w\[491\] net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_112_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold144 hotp.block.sha1.mixer.w\[131\] net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1728_ _1488_ _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold122 hotp.block.sha1.mixer.w\[506\] net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold133 hotp.block.sha1.mixer.w\[48\] net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold111 hotp.block.sha1.mixer.w\[11\] net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_44_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold155 stream.key_buf\[123\] net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold166 hotp.block.sha1.mixer.w\[118\] net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1659_ _1418_ _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4447_ _0348_ clknet_leaf_97_clk hotp.block.mixer.msg\[159\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold177 hotp.block.sha1.mixer.w\[363\] net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold188 hotp.block.sha1.mixer.w\[352\] net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold199 hotp.block.sha1.mixer.c\[3\] net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4378_ _0279_ clknet_leaf_60_clk hotp.block.mixer.msg\[90\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3329_ _0070_ clknet_leaf_40_clk stream.msg_buf\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_53_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_37_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1992__A1 _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_62_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1744__A1 _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_71_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4137__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2700_ _1006_ _1033_ _1034_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3680_ net683 clknet_leaf_84_clk hotp.block.sha1.mixer.c\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2631_ _0883_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2562_ _0897_ _0906_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4301_ _0202_ clknet_leaf_104_clk hotp.block.mixer.msg\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2493_ _0850_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4232_ net72 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[459\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4_clk clknet_4_0_0_clk clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_4_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ net176 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[390\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4094_ net516 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[321\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3114_ hotp.block.mixer.msg\[110\] hotp.block.mixer.msg\[111\] _1303_ _1307_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold177_I hotp.block.sha1.mixer.w\[363\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3045_ _1268_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold609_I hotp.block.sha1.mixer.w\[440\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3947_ net198 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[174\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3878_ net634 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[105\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2829_ _1136_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_115_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3801_ net106 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1993_ _0442_ _0439_ _1513_ _1550_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_15_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3732_ net458 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3663_ net729 clknet_leaf_78_clk hotp.block.sha1.mixer.b\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_99_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2614_ _0945_ _0957_ _0958_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3594_ _0167_ clknet_leaf_50_clk stream.key_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2545_ hotp.digest\[7\] _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2476_ _0808_ _0833_ _0810_ _0811_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_110_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4215_ net169 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[442\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold461_I hotp.block.sha1.mixer.w\[148\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4146_ net506 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[373\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4452__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4077_ net127 clknet_leaf_41_clk hotp.block.sha1.mixer.w\[304\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold726_I hotp.block.sha1.mixer.w\[202\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3028_ _1258_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2675__A2 _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4134__D net401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3973__D net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2330_ stream.digest\[19\] stream.digest\[20\] _0712_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2261_ _0657_ _0669_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4000_ net145 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[227\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2192_ stream.counter\[1\] stream.counter\[0\] _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_9_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ _0454_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold307_I hotp.block.sha1.mixer.w\[396\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3715_ net636 clknet_leaf_86_clk hotp.block.sha1.mixer.d\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3646_ net816 clknet_leaf_93_clk hotp.block.sha1.mixer.b\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3577_ _0150_ clknet_leaf_63_clk hotp.digest\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2528_ _0839_ _0881_ _0882_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_hold676_I hotp.block.sha1.mixer.w\[92\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold15 hotp.block.sha1.mixer.w\[297\] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2459_ _0808_ _0810_ _0815_ _0816_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xhold37 hotp.block.sha1.mixer.w\[456\] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold26 hotp.block.sha1.mixer.w\[42\] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3842__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold48 hotp.block.sha1.mixer.w\[303\] net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold59 hotp.block.sha1.mixer.w\[453\] net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4219__D net322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4129_ net365 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[356\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_6_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__D net739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ hotp.block.sha1.mixer.e\[0\] _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3500_ net565 clknet_leaf_20_clk stream.key_buf\[152\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1761_ hotp.block.mixer.msg\[128\] _1519_ _1520_ _1521_ _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_96_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1692_ _1456_ _1459_ _1443_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold507 hotp.block.sha1.mixer.w\[237\] net527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold518 hotp.block.sha1.mixer.e\[5\] net538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3431_ net615 clknet_leaf_35_clk stream.key_buf\[83\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold529 hotp.block.sha1.mixer.w\[185\] net549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3362_ net826 clknet_leaf_49_clk stream.key_buf\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2313_ _0690_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3293_ _0034_ clknet_leaf_38_clk stream.msg_buf\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2244_ stream.digest\[16\] stream.digest\[20\] stream.digest\[24\] stream.digest\[28\]
+ _0653_ _0654_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2175_ _0594_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_49_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3878__D net634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3395__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1959_ hotp.block.sha1.mixer.b\[0\] hotp.block.sha1.mixer.c\[0\] _0438_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3629_ net414 clknet_leaf_77_clk hotp.block.sha1.mixer.a\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput16 net16 out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3788__D net792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3980_ net203 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[207\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2931_ _1202_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_99_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2862_ hotp.block.mixer.msg\[1\] hotp.block.mixer.msg\[2\] _1162_ _1164_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2793_ hotp.index\[0\] _0809_ _1110_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1813_ hotp.block.magic.step\[0\] _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1744_ _1497_ _1499_ _1504_ _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_13_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold304 stream.key_buf\[102\] net324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold315 stream.key_buf\[1\] net335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4463_ _0363_ clknet_leaf_71_clk hotp.block.magic.step\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold326 hotp.block.sha1.mixer.w\[505\] net346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3414_ net818 clknet_leaf_53_clk stream.key_buf\[66\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1675_ _1436_ _1437_ _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold337 hotp.block.sha1.mixer.w\[479\] net357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold348 hotp.block.sha1.mixer.w\[70\] net368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_1_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold359 hotp.block.sha1.mixer.b\[26\] net379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_68_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ _0295_ clknet_leaf_61_clk hotp.block.mixer.msg\[106\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3345_ _0082_ clknet_leaf_16_clk seg.digit\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3276_ _0017_ clknet_leaf_39_clk stream.msg_buf\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold374_I hotp.block.sha1.mixer.w\[407\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2227_ _0640_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_107_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4193__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2158_ stream.msg_buf\[51\] stream.msg_buf\[52\] _0582_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2089_ stream.msg_buf\[21\] stream.msg_buf\[22\] _0545_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_24_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4232__D net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_hold3_I hotp.block.sha1.mixer.w\[253\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4142__D net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4066__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3981__D net748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3130_ _1316_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3061_ _1266_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_54_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2012_ _0489_ _0474_ _0490_ _1621_ _1562_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_102_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3963_ net390 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[190\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3894_ net226 clknet_leaf_27_clk hotp.block.sha1.mixer.w\[121\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2914_ _1193_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_93_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2845_ _1143_ _1145_ _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2776_ _0639_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold101 hotp.block.sha1.mixer.w\[294\] net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold112 hotp.block.sha1.mixer.w\[264\] net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1727_ _1475_ _1477_ _1486_ _1489_ net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold134 hotp.block.sha1.mixer.w\[402\] net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold123 hotp.block.sha1.mixer.w\[381\] net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_106_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold167 stream.key_buf\[20\] net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1658_ stream.msg_state\[2\] _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold589_I hotp.block.sha1.mixer.w\[203\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold156 hotp.block.sha1.mixer.w\[391\] net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold145 hotp.block.sha1.mixer.a\[28\] net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4446_ _0347_ clknet_leaf_95_clk hotp.block.mixer.msg\[158\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold189 stream.key_buf\[79\] net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4377_ _0278_ clknet_leaf_60_clk hotp.block.mixer.msg\[89\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold178 hotp.block.sha1.mixer.w\[175\] net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_113_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3328_ _0069_ clknet_leaf_40_clk stream.msg_buf\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_31_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3259_ _1610_ _1588_ _1375_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_clkbuf_leaf_46_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4089__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_104_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold690 hotp.block.sha1.mixer.w\[490\] net710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1902__I _1578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4137__D net622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3976__D net484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2630_ _0945_ _0971_ _0972_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2561_ _0908_ _0898_ _0911_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2492_ _0829_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4300_ _0201_ clknet_leaf_104_clk hotp.block.mixer.msg\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4231_ net497 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[458\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4162_ net205 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[389\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4093_ net831 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[320\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3113_ _1306_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3044_ hotp.block.mixer.msg\[79\] hotp.block.mixer.msg\[80\] _1267_ _1268_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold337_I hotp.block.sha1.mixer.w\[479\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3946_ net626 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[173\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold504_I hotp.block.sha1.mixer.w\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3877_ net478 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[104\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2828_ hotp.digest\[38\] _0857_ _1129_ hotp.digest\[37\] _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2759_ _0850_ _1086_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_57_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4429_ _0330_ clknet_leaf_69_clk hotp.block.mixer.msg\[141\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_70_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output19_I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3800_ net325 clknet_leaf_107_clk hotp.block.sha1.mixer.w\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1992_ _1556_ _0466_ _0467_ _0470_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3731_ net707 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1956__A2 _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3662_ net758 clknet_leaf_78_clk hotp.block.sha1.mixer.b\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_99_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3593_ _0166_ clknet_leaf_46_clk stream.key_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2613_ hotp.digest\[13\] _0937_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1807__I hotp.block.magic.step\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2544_ _0884_ _0895_ _0896_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2475_ _0375_ hotp.index\[0\] _0427_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_110_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4214_ net691 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[441\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold287_I hotp.block.sha1.mixer.w\[224\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4145_ net762 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[372\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold454_I hotp.block.sha1.mixer.w\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4076_ net645 clknet_leaf_41_clk hotp.block.sha1.mixer.w\[303\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3027_ hotp.block.mixer.msg\[72\] hotp.block.mixer.msg\[73\] _1256_ _1258_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold719_I hotp.block.sha1.mixer.w\[196\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold621_I hotp.block.sha1.mixer.w\[160\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3929_ net594 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[156\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4240__D net529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1880__C _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4277__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold63_I stream.key_buf\[147\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4150__D net770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2260_ stream.digest\[2\] stream.digest\[6\] stream.digest\[10\] stream.digest\[14\]
+ _0658_ _0659_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2191_ _0604_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1975_ _1512_ _0441_ _0447_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_114_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3714_ net442 clknet_leaf_86_clk hotp.block.sha1.mixer.d\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold202_I hotp.block.sha1.mixer.w\[187\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3645_ net40 clknet_leaf_69_clk hotp.block.sha1.mixer.b\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3576_ _0149_ clknet_leaf_63_clk hotp.digest\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2527_ _0867_ _0876_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2458_ _1499_ hotp.index\[3\] _1518_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold571_I hotp.block.sha1.mixer.w\[101\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold27 hotp.block.sha1.mixer.w\[275\] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold16 hotp.block.sha1.mixer.w\[88\] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold38 hotp.block.sha1.mixer.c\[19\] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2389_ _0747_ _0751_ _0757_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold49 hotp.block.sha1.mixer.w\[462\] net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_97_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4128_ net539 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[355\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4059_ net576 clknet_leaf_19_clk hotp.block.sha1.mixer.w\[286\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4235__D net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_65_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3667__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4145__D net762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2281__A1 _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3984__D net688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1760_ _1496_ _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1691_ _1405_ _1458_ _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold508 hotp.block.sha1.mixer.w\[60\] net528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3430_ net334 clknet_leaf_35_clk stream.key_buf\[82\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold519 hotp.block.sha1.mixer.w\[356\] net539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3361_ net745 clknet_leaf_49_clk stream.key_buf\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2312_ _0705_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3292_ _0033_ clknet_leaf_36_clk stream.msg_buf\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2243_ net5 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2174_ stream.msg_buf\[58\] stream.msg_buf\[59\] _0592_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_49_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3894__D net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1958_ hotp.block.sha1.mixer.b\[0\] hotp.block.sha1.mixer.d\[0\] hotp.block.sha1.mixer.c\[0\]
+ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_43_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1889_ _1545_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3628_ net511 clknet_leaf_77_clk hotp.block.sha1.mixer.a\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput17 net17 out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_3559_ _0006_ clknet_leaf_45_clk stream.key_state\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_67_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2015__A1 _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2002__S _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold26_I hotp.block.sha1.mixer.w\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3979__D net713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2930_ _1160_ _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2006__A1 _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2861_ _1158_ _1162_ _1163_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2792_ _1109_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1812_ _1496_ _1535_ _1572_ _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3832__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1743_ _1501_ _1503_ _1504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_41_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1674_ _1433_ _1440_ _1443_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4462_ _0362_ clknet_leaf_62_clk hotp.block.magic.step\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xhold305 hotp.block.sha1.mixer.w\[28\] net325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold316 hotp.block.sha1.mixer.w\[9\] net336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3413_ net230 clknet_leaf_52_clk stream.key_buf\[65\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold327 stream.key_buf\[146\] net347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold338 hotp.block.sha1.mixer.w\[66\] net358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold349 hotp.block.sha1.mixer.w\[161\] net369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4393_ _0294_ clknet_leaf_61_clk hotp.block.mixer.msg\[105\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3344_ _0081_ clknet_leaf_16_clk seg.digit\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3275_ _0016_ clknet_leaf_39_clk stream.msg_buf\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2226_ stream.key_counter\[7\] _1407_ _0639_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_107_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2157_ _0584_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2088_ _0529_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_89_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold534_I hotp.block.sha1.mixer.w\[217\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_5_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_110_clk clknet_4_0_0_clk clknet_leaf_110_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1725__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_101_clk clknet_4_3_0_clk clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_10_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3060_ _1276_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2011_ _0458_ _0455_ _0453_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output9_I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3962_ net836 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[189\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3893_ net133 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[120\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2913_ hotp.block.mixer.msg\[23\] hotp.block.mixer.msg\[24\] _1192_ _1193_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2844_ hotp.block.sha1.mixer.a_carry\[1\] _0503_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3027__I0 hotp.block.mixer.msg\[72\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2775_ _0638_ _1095_ _1097_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_81_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold113 hotp.block.sha1.mixer.w\[121\] net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1726_ seg.digit\[3\] _1487_ _1488_ _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold124 hotp.block.sha1.mixer.w\[384\] net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold102 hotp.block.sha1.mixer.c\[8\] net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold135 hotp.block.sha1.mixer.w\[472\] net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1657_ net3 _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold168 hotp.block.sha1.mixer.a\[10\] net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold157 hotp.block.sha1.mixer.w\[103\] net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold146 hotp.block.sha1.mixer.e\[26\] net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4445_ _0346_ clknet_leaf_95_clk hotp.block.mixer.msg\[157\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4376_ _0277_ clknet_leaf_60_clk hotp.block.mixer.msg\[88\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold179 hotp.block.sha1.mixer.w\[486\] net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3327_ _0068_ clknet_leaf_40_clk stream.msg_buf\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3728__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3258_ _1391_ _1393_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2209_ _0615_ _0622_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3189_ _1349_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4243__D net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold680 hotp.block.sha1.mixer.w\[483\] net700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold691 hotp.block.sha1.mixer.w\[242\] net711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_19_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold93_I hotp.block.sha1.mixer.w\[77\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2235__B _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4153__D net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3992__D net429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2560_ _0909_ _0910_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2491_ hotp.digest\[39\] _0848_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4230_ net338 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[457\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4161_ net623 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[388\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4092_ net521 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[319\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3112_ hotp.block.mixer.msg\[109\] hotp.block.mixer.msg\[110\] _1303_ _1306_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3043_ _1266_ _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_59_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold232_I hotp.block.sha1.mixer.w\[248\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3945_ net668 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[172\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3400__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3876_ net553 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[103\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2827_ _1135_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2758_ _1083_ _1084_ _1085_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1709_ _1472_ _1445_ _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2689_ _0991_ _1024_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4428_ _0329_ clknet_leaf_78_clk hotp.block.mixer.msg\[140\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4359_ _0260_ clknet_leaf_74_clk hotp.block.mixer.msg\[71\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_100_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4238__D net803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_92_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4148__D net343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3987__D net397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3730_ net472 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1991_ _0468_ _0469_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_30_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3661_ net679 clknet_leaf_78_clk hotp.block.sha1.mixer.b\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2612_ hotp.digest\[14\] _0940_ _0956_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3592_ _0165_ clknet_leaf_66_clk hotp.digest\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2543_ hotp.digest\[5\] _0876_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_45_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2474_ _0824_ _0830_ _0831_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_110_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4213_ net718 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[440\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3016__S _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4144_ net772 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[371\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4075_ net68 clknet_leaf_33_clk hotp.block.sha1.mixer.w\[302\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1892__A2 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_103_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3026_ _1257_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_90_clk clknet_4_8_0_clk clknet_leaf_90_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_hold614_I hotp.block.sha1.mixer.w\[106\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3928_ net518 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[155\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3859_ net271 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[86\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2564__I _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_81_clk clknet_4_10_0_clk clknet_leaf_81_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4221__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2190_ stream.counter\[6\] _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3939__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2407__C _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_72_clk clknet_4_11_0_clk clknet_leaf_72_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1974_ _0452_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ net778 clknet_leaf_86_clk hotp.block.sha1.mixer.d\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3644_ _0008_ clknet_leaf_95_clk hotp.block.sha1.mixer.a\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3575_ _0148_ clknet_leaf_64_clk hotp.digest\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2526_ _0878_ _0860_ _0880_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold397_I hotp.block.sha1.mixer.w\[233\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2457_ hotp.index\[0\] _0809_ _0814_ _0364_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_54_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold17 hotp.block.sha1.mixer.w\[62\] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_hold564_I hotp.block.sha1.mixer.w\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold28 hotp.block.sha1.mixer.w\[397\] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold39 hotp.block.sha1.mixer.w\[333\] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2388_ _0619_ _0606_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4127_ net261 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[354\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4058_ net421 clknet_leaf_19_clk hotp.block.sha1.mixer.w\[285\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3009_ hotp.block.mixer.msg\[64\] hotp.block.mixer.msg\[65\] _1246_ _1248_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_63_clk clknet_4_15_0_clk clknet_leaf_63_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4251__D net357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1891__C _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_54_clk clknet_4_13_0_clk clknet_leaf_54_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4161__D net623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1690_ _1422_ _1457_ _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1792__A1 _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold509 hotp.block.sha1.mixer.w\[468\] net529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3360_ net202 clknet_leaf_51_clk stream.key_buf\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2311_ stream.digest\[11\] stream.digest\[12\] _0701_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3291_ _0032_ clknet_leaf_37_clk stream.msg_buf\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2242_ net4 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2173_ _0593_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_45_clk clknet_4_12_0_clk clknet_leaf_45_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold312_I hotp.block.sha1.mixer.w\[368\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4267__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1957_ hotp.block.sha1.mixer.b\[27\] hotp.block.sha1.mixer.a\[27\] _0435_ _0436_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1888_ _1588_ _0379_ _0380_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3627_ net225 clknet_leaf_76_clk hotp.block.sha1.mixer.a\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput18 net18 out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3558_ _0005_ clknet_leaf_47_clk stream.key_state\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2509_ hotp.digest\[1\] _0857_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3489_ net400 clknet_leaf_26_clk stream.key_buf\[141\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4246__D net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_clk clknet_4_7_0_clk clknet_leaf_36_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_27_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4156__D net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_27_clk clknet_4_4_0_clk clknet_leaf_27_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3995__D net422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2860_ hotp.block.mixer.msg\[1\] _1162_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1811_ hotp.block.mixer.round\[0\] _1542_ _1572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2791_ _0824_ _1107_ _1108_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_4_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1742_ _1502_ _1503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1765__A1 hotp.block.mixer.msg\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold317 hotp.block.sha1.mixer.w\[145\] net337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1673_ _1442_ _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4461_ _0361_ clknet_leaf_71_clk hotp.block.magic.step\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xhold306 hotp.block.sha1.mixer.d\[17\] net326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3412_ net643 clknet_leaf_52_clk stream.key_buf\[64\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold328 stream.key_buf\[49\] net348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_22_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold339 hotp.block.sha1.mixer.w\[492\] net359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4392_ _0293_ clknet_leaf_61_clk hotp.block.mixer.msg\[104\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3343_ _0080_ clknet_leaf_44_clk stream.state\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3274_ _0015_ clknet_leaf_39_clk stream.msg_buf\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2225_ stream.key_counter\[4\] _0638_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_107_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2156_ stream.msg_buf\[50\] stream.msg_buf\[51\] _0582_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2087_ _0544_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_18_clk clknet_4_4_0_clk clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_hold527_I hotp.block.sha1.mixer.w\[69\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2989_ hotp.block.mixer.msg\[56\] hotp.block.mixer.msg\[57\] _1234_ _1236_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_118_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1942__S _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4432__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1995__A1 _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ _0458_ _0444_ _0382_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3961_ net510 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[188\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_102_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2912_ _1181_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3892_ net311 clknet_leaf_21_clk hotp.block.sha1.mixer.w\[119\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3027__I1 hotp.block.mixer.msg\[73\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2843_ _1138_ _1148_ _0734_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2774_ stream.key_counter\[3\] _0637_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1725_ net7 _1488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold114 hotp.block.sha1.mixer.w\[302\] net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_79_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold103 hotp.block.sha1.mixer.w\[461\] net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold125 hotp.block.sha1.mixer.w\[228\] net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold158 hotp.block.sha1.mixer.w\[308\] net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1656_ _1421_ _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold136 hotp.block.sha1.mixer.w\[49\] net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold147 hotp.block.sha1.mixer.d\[8\] net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4444_ _0345_ clknet_leaf_95_clk hotp.block.mixer.msg\[156\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_7_clk clknet_4_1_0_clk clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4375_ _0276_ clknet_leaf_60_clk hotp.block.mixer.msg\[87\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold169 hotp.block.sha1.mixer.w\[236\] net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_42_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3326_ _0067_ clknet_leaf_40_clk stream.msg_buf\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold477_I hotp.block.sha1.mixer.w\[459\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3257_ _0685_ _1392_ _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2208_ _0616_ _0618_ _0621_ _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3188_ hotp.block.mixer.msg\[142\] hotp.block.mixer.msg\[143\] _1345_ _1349_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2139_ _0574_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1977__A1 _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold670 stream.key_buf\[75\] net690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold681 stream.key_buf\[136\] net701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_102_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_31_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold692 stream.key_buf\[25\] net712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2490_ hotp.digest\[2\] _0844_ _0845_ _0372_ _0847_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_4160_ net823 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[387\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3111_ _1305_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4091_ net393 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[318\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3042_ _1244_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2426__B _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3944_ net786 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[171\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3875_ net177 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[102\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold225_I hotp.block.sha1.mixer.w\[258\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2826_ hotp.digest\[37\] _1122_ _1129_ hotp.digest\[36\] _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_116_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2757_ _1067_ _1070_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1708_ stream.msg_state\[1\] _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2688_ hotp.digest\[21\] _1022_ _1023_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1639_ _1409_ _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4427_ _0328_ clknet_leaf_77_clk hotp.block.mixer.msg\[139\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3845__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4358_ _0259_ clknet_leaf_74_clk hotp.block.mixer.msg\[70\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3309_ _0050_ clknet_leaf_34_clk stream.msg_buf\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4289_ _0190_ clknet_leaf_95_clk hotp.block.mixer.msg\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1990_ _0440_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4164__D net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4150__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3660_ net44 clknet_leaf_77_clk hotp.block.sha1.mixer.b\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2611_ _0954_ _0955_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3591_ _0164_ clknet_leaf_66_clk hotp.digest\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2542_ hotp.digest\[6\] _0860_ _0894_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3868__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2473_ _1505_ _0823_ _0827_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_55_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4212_ net629 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[439\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4143_ net649 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[370\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4074_ net134 clknet_leaf_41_clk hotp.block.sha1.mixer.w\[301\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3025_ hotp.block.mixer.msg\[71\] hotp.block.mixer.msg\[72\] _1256_ _1257_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold342_I hotp.block.sha1.mixer.w\[420\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3398__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3927_ net475 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[154\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3858_ net447 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[85\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2809_ _1005_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_59_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3789_ net395 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4023__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold49_I hotp.block.sha1.mixer.w\[462\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4159__D net735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3998__D net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ _0442_ _0439_ _1513_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_44_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3712_ net644 clknet_leaf_93_clk hotp.block.sha1.mixer.d\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3643_ net147 clknet_leaf_94_clk hotp.block.sha1.mixer.a\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3574_ _0147_ clknet_leaf_57_clk hotp.digest\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2525_ _0868_ _0879_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3027__S _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2456_ hotp.index\[2\] _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_54_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold29 stream.key_buf\[5\] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold18 hotp.block.sha1.mixer.w\[198\] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_2387_ _0619_ _0748_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4126_ net508 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[353\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4196__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4057_ net364 clknet_leaf_19_clk hotp.block.sha1.mixer.w\[284\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3008_ _1247_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_91_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_44_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_59_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_102_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3290_ _0031_ clknet_leaf_37_clk stream.msg_buf\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2310_ _0704_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3906__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2241_ net6 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2172_ stream.msg_buf\[57\] stream.msg_buf\[58\] _0592_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_49_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_69_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1829__I _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold138_I hotp.block.sha1.mixer.w\[261\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1956_ _0371_ _1548_ _0369_ _0375_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_7_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_78_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1887_ _0375_ _0371_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3626_ net513 clknet_leaf_76_clk hotp.block.sha1.mixer.a\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput19 net19 out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_3557_ _0004_ clknet_leaf_45_clk stream.key_state\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2508_ hotp.digest\[2\] _0860_ _0864_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_hold674_I hotp.block.sha1.mixer.w\[380\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3488_ net86 clknet_leaf_28_clk stream.key_buf\[140\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2439_ _0752_ _0798_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4109_ net61 clknet_leaf_21_clk hotp.block.sha1.mixer.w\[336\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_67_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1810_ _1557_ _1536_ _1554_ _1571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2790_ hotp.rst_n _0826_ _1538_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_53_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1741_ hotp.block.mixer.round\[2\] _1502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1672_ _1441_ _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4460_ _0360_ clknet_leaf_71_clk hotp.block.magic.step\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold307 hotp.block.sha1.mixer.w\[396\] net327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3411_ net544 clknet_leaf_52_clk stream.key_buf\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4391_ _0292_ clknet_leaf_61_clk hotp.block.mixer.msg\[103\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold318 hotp.block.sha1.mixer.w\[458\] net338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold329 hotp.block.sha1.mixer.d\[16\] net349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_68_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3342_ _0079_ clknet_leaf_44_clk stream.state\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3273_ _0014_ clknet_leaf_46_clk stream.msg_buf\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2224_ stream.key_counter\[3\] _0637_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_107_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2155_ _0583_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold255_I hotp.block.sha1.mixer.w\[383\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2086_ stream.msg_buf\[20\] stream.msg_buf\[21\] _0540_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_86_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2988_ _1235_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1939_ _0416_ _0421_ _0422_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3609_ _0182_ clknet_leaf_45_clk hotp.digest\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2705__A1 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_95_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1995__A2 _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_93_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4167__D net560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3960_ net409 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[187\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_102_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2911_ _1191_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3891_ net807 clknet_leaf_21_clk hotp.block.sha1.mixer.w\[118\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2842_ _0502_ _1146_ _1147_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2773_ _0637_ _1095_ _1096_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_72_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1724_ seg.digit\[2\] _1481_ _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_14_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold126 stream.key_buf\[43\] net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold104 stream.key_buf\[4\] net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold115 hotp.block.sha1.mixer.c\[6\] net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1655_ _1402_ _1423_ _1425_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold159 hotp.block.sha1.mixer.w\[211\] net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold137 hotp.block.sha1.mixer.w\[64\] net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold148 hotp.block.sha1.mixer.w\[417\] net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4443_ _0344_ clknet_leaf_95_clk hotp.block.mixer.msg\[155\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4374_ _0275_ clknet_leaf_59_clk hotp.block.mixer.msg\[86\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3325_ _0066_ clknet_leaf_41_clk stream.msg_buf\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold372_I hotp.block.sha1.mixer.w\[361\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3256_ _1589_ _1375_ _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2207_ stream.counter\[4\] stream.counter\[3\] _0619_ _0620_ _0621_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3187_ _1348_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2138_ stream.msg_buf\[42\] stream.msg_buf\[43\] _0572_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2069_ _0534_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold804_I hotp.block.sha1.mixer.w\[162\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold671 hotp.block.sha1.mixer.w\[442\] net691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold660 hotp.block.sha1.mixer.w\[199\] net680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold682 hotp.block.sha1.mixer.d\[15\] net702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold693 hotp.block.sha1.mixer.w\[207\] net713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_87_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3110_ hotp.block.mixer.msg\[108\] hotp.block.mixer.msg\[109\] _1303_ _1305_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4090_ net419 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[317\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3041_ _1265_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3943_ net446 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[170\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1959__A2 hotp.block.sha1.mixer.c\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3874_ net228 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[101\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2825_ _1134_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_hold218_I hotp.block.sha1.mixer.w\[197\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold120_I hotp.block.sha1.mixer.w\[422\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2756_ _1066_ _1076_ _1050_ hotp.digest\[28\] _1069_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_5_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1707_ _1469_ _1470_ _1471_ _1403_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2687_ _1007_ _1009_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_42_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1638_ _1406_ _1407_ _1408_ _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4426_ _0327_ clknet_leaf_77_clk hotp.block.mixer.msg\[138\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4357_ _0258_ clknet_leaf_74_clk hotp.block.mixer.msg\[69\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3308_ _0049_ clknet_leaf_34_clk stream.msg_buf\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4288_ _0189_ clknet_leaf_97_clk hotp.block.mixer.msg\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3239_ _1508_ _1378_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4270__D net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold490 hotp.block.sha1.mixer.w\[189\] net510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1657__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4180__D net603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2610_ _0939_ _0949_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3590_ _0163_ clknet_leaf_45_clk hotp.digest\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2541_ _0868_ _0893_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2472_ _0829_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4211_ net310 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[438\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4142_ net108 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[369\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4073_ net637 clknet_leaf_41_clk hotp.block.sha1.mixer.w\[300\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3024_ _1245_ _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_50_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold335_I hotp.block.sha1.mixer.w\[250\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3926_ net663 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[153\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold502_I hotp.block.sha1.mixer.w\[180\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3857_ net402 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[84\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2808_ _1121_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_59_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3788_ net792 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2739_ _0365_ _0846_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4409_ _0310_ clknet_leaf_62_clk hotp.block.mixer.msg\[121\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1868__A1 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output17_I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3835__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1972_ _0438_ _0445_ _0450_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_44_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3711_ net45 clknet_leaf_85_clk hotp.block.sha1.mixer.d\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3642_ net489 clknet_leaf_94_clk hotp.block.sha1.mixer.a\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3573_ _0146_ clknet_leaf_64_clk hotp.digest\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2524_ hotp.digest\[2\] _0871_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2455_ _1628_ _0807_ _0812_ _0397_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2386_ _0735_ _0755_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_hold285_I hotp.block.sha1.mixer.w\[89\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold19 hotp.block.sha1.mixer.a\[23\] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4125_ net350 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[352\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3270__C _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4056_ net750 clknet_leaf_19_clk hotp.block.sha1.mixer.w\[283\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4085__D net502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3007_ hotp.block.mixer.msg\[63\] hotp.block.mixer.msg\[64\] _1246_ _1247_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3909_ net543 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[136\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3708__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_115_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2240_ _0649_ _0651_ _1443_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2171_ _0515_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_49_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2009__A1 _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1955_ _0419_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1886_ _0374_ _0377_ _0378_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_hold200_I hotp.block.sha1.mixer.w\[218\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3625_ net183 clknet_leaf_75_clk hotp.block.sha1.mixer.a\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3556_ _0133_ clknet_leaf_17_clk stream.counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2507_ _0862_ _0863_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3487_ net652 clknet_leaf_29_clk stream.key_buf\[139\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2438_ _0795_ _0611_ _0787_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2369_ stream.counter\[0\] _0739_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4108_ net569 clknet_leaf_21_clk hotp.block.sha1.mixer.w\[335\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4039_ net493 clknet_leaf_14_clk hotp.block.sha1.mixer.w\[266\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_113_clk clknet_4_0_0_clk clknet_leaf_113_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_34_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2487__A1 _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_104_clk clknet_4_2_0_clk clknet_leaf_104_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4186__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1740_ _1500_ _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold308 stream.key_buf\[121\] net328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_80_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1671_ net8 _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_34_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3410_ net351 clknet_leaf_52_clk stream.key_buf\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4390_ _0291_ clknet_leaf_61_clk hotp.block.mixer.msg\[102\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold319 hotp.block.sha1.mixer.w\[465\] net339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3341_ _0078_ clknet_leaf_44_clk stream.debug\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_0_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3272_ _0378_ _1399_ _0734_ _1395_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2223_ stream.key_counter\[2\] _0636_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2154_ stream.msg_buf\[49\] stream.msg_buf\[50\] _0582_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_107_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_90_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2085_ _0543_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3403__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold415_I hotp.block.sha1.mixer.w\[436\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2987_ hotp.block.mixer.msg\[55\] hotp.block.mixer.msg\[56\] _1234_ _1235_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1938_ hotp.block.sha1.mixer.c\[30\] _0421_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1869_ _1499_ _1628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3608_ _0181_ clknet_leaf_45_clk hotp.digest\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_43_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3539_ _0116_ clknet_leaf_14_clk stream.digest\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_58_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_101_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4273__D net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2910_ hotp.block.mixer.msg\[22\] hotp.block.mixer.msg\[23\] _1187_ _1191_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4183__D net695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3890_ net186 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[117\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2841_ _0502_ _1146_ _0503_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2772_ stream.key_counter\[2\] _0636_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1723_ _1478_ _1485_ _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_54_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold105 hotp.block.sha1.mixer.w\[10\] net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold116 hotp.block.sha1.mixer.w\[425\] net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4442_ _0343_ clknet_leaf_91_clk hotp.block.mixer.msg\[154\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1654_ _1424_ _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold149 hotp.block.sha1.mixer.w\[443\] net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold138 hotp.block.sha1.mixer.w\[261\] net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold127 hotp.block.sha1.mixer.a\[31\] net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4373_ _0274_ clknet_leaf_59_clk hotp.block.mixer.msg\[85\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3324_ _0065_ clknet_leaf_42_clk stream.msg_buf\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3255_ _1589_ _1375_ _1391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2206_ stream.counter\[10\] stream.counter\[9\] stream.counter\[8\] _0399_ _0620_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3186_ hotp.block.mixer.msg\[141\] hotp.block.mixer.msg\[142\] _1345_ _1348_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2137_ _0573_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2068_ stream.msg_buf\[12\] stream.msg_buf\[13\] _0530_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3919__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold661 stream.key_buf\[98\] net681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold672 hotp.block.sha1.mixer.w\[124\] net692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold650 hotp.block.sha1.mixer.e\[10\] net670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold683 hotp.block.sha1.mixer.w\[274\] net703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold694 hotp.block.sha1.mixer.w\[222\] net714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3900__D net455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3040_ hotp.block.mixer.msg\[78\] hotp.block.mixer.msg\[79\] _1261_ _1265_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3810__D net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3942_ net102 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[169\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3873_ net591 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[100\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2824_ hotp.digest\[36\] _1122_ _1116_ hotp.digest\[35\] _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2755_ _1066_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1706_ _1405_ _1411_ _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2686_ _1021_ _1009_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1637_ stream.key_counter\[1\] stream.key_counter\[0\] _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_74_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4425_ _0326_ clknet_leaf_69_clk hotp.block.mixer.msg\[137\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold482_I hotp.block.sha1.mixer.w\[313\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4356_ _0257_ clknet_leaf_74_clk hotp.block.mixer.msg\[68\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3307_ _0048_ clknet_leaf_36_clk stream.msg_buf\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4287_ _0188_ clknet_leaf_97_clk hotp.block.sha1.mixer.a_carry\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3238_ _1377_ _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3169_ _1338_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_93_clk clknet_4_9_0_clk clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold480 hotp.block.sha1.mixer.e\[16\] net500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold491 hotp.block.sha1.mixer.a\[16\] net511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_59_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_84_clk clknet_4_10_0_clk clknet_leaf_84_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_hold91_I hotp.block.sha1.mixer.w\[450\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2540_ _0878_ _0888_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_23_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1673__I _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2471_ _0822_ _1604_ hotp.block.mixer.stage\[0\] _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__3805__D net632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4210_ net148 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[437\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4141_ net354 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[368\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4072_ net388 clknet_leaf_41_clk hotp.block.sha1.mixer.w\[299\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3023_ _1255_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_75_clk clknet_4_11_0_clk clknet_leaf_75_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3925_ net423 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[152\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3856_ net31 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[83\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2807_ hotp.digest\[32\] _1065_ _1116_ _1120_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3787_ net372 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2738_ _1067_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ _0309_ clknet_leaf_62_clk hotp.block.mixer.msg\[120\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2669_ hotp.digest\[19\] hotp.digest\[20\] hotp.digest\[21\] _1007_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4339_ _0240_ clknet_leaf_86_clk hotp.block.mixer.msg\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_clk clknet_4_12_0_clk clknet_leaf_66_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2363__B _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3637__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_57_clk clknet_4_15_0_clk clknet_leaf_57_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_62_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3710_ net468 clknet_leaf_85_clk hotp.block.sha1.mixer.d\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1971_ hotp.block.sha1.mixer.b\[0\] hotp.block.sha1.mixer.c\[0\] _0449_ _0450_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4191__D net534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3641_ net383 clknet_leaf_94_clk hotp.block.sha1.mixer.a\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3572_ _0145_ clknet_leaf_57_clk hotp.digest\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2523_ hotp.digest\[4\] _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2454_ _0808_ _0810_ _0811_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2385_ stream.counter\[1\] _0748_ _0751_ _0754_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4124_ net208 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[351\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold180_I hotp.block.sha1.mixer.w\[181\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 in[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_48_clk clknet_4_13_0_clk clknet_leaf_48_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4055_ net250 clknet_leaf_17_clk hotp.block.sha1.mixer.w\[282\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4092__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3006_ _1245_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_hold445_I hotp.block.sha1.mixer.w\[216\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold612_I hotp.block.sha1.mixer.w\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3908_ net551 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[135\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3839_ net559 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[66\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_39_clk clknet_4_7_0_clk clknet_leaf_39_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_2_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_9_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2170_ _0591_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_109_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1954_ _0433_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1885_ _1560_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3624_ net231 clknet_leaf_76_clk hotp.block.sha1.mixer.a\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3555_ _0132_ clknet_leaf_16_clk stream.counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3486_ net415 clknet_leaf_29_clk stream.key_buf\[138\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2506_ hotp.digest\[0\] _0849_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_12_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2437_ _0603_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2368_ _1438_ _0505_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3482__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4107_ net116 clknet_leaf_20_clk hotp.block.sha1.mixer.w\[334\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2299_ _0698_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4038_ net558 clknet_leaf_14_clk hotp.block.sha1.mixer.w\[265\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_2_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3028__I _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3825__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1998__A1 _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1670_ _1434_ stream.msg_state\[3\] _1430_ _1439_ _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold309 stream.key_buf\[9\] net329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3340_ _0003_ clknet_leaf_43_clk stream.msg_state\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3271_ _1400_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3813__D net524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2222_ stream.key_counter\[1\] stream.key_counter\[0\] _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_84_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2153_ _0571_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2084_ stream.msg_buf\[19\] stream.msg_buf\[20\] _0540_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4130__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2986_ _1223_ _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1937_ _0419_ _0420_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_17_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1868_ _1617_ _1514_ _1533_ _1626_ _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3607_ _0180_ clknet_leaf_45_clk hotp.digest\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold810 hotp.block.sha1.mixer.w\[168\] net830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_31_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3538_ _0115_ clknet_leaf_14_clk stream.digest\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1799_ _1559_ _1560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_hold777_I hotp.block.sha1.mixer.w\[421\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3848__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1913__A1 _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3469_ net839 clknet_leaf_29_clk stream.key_buf\[121\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2641__A2 _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold17_I hotp.block.sha1.mixer.w\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2840_ _1143_ _1145_ _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_72_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2771_ _1408_ _0636_ _1095_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_26_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1722_ _1479_ _1480_ _1484_ _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold106 stream.key_buf\[60\] net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1653_ net8 _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold117 hotp.block.sha1.mixer.w\[177\] net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4441_ _0342_ clknet_leaf_91_clk hotp.block.mixer.msg\[153\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_117_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold128 hotp.block.sha1.mixer.w\[438\] net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold139 hotp.block.sha1.mixer.e\[17\] net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4372_ _0273_ clknet_leaf_60_clk hotp.block.mixer.msg\[84\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3323_ _0064_ clknet_leaf_42_clk stream.msg_buf\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3254_ _1380_ _1390_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2205_ stream.counter\[2\] _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3185_ _1347_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2136_ stream.msg_buf\[41\] stream.msg_buf\[42\] _0572_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2067_ _0533_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold525_I hotp.block.sha1.mixer.w\[195\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2969_ hotp.block.mixer.msg\[47\] hotp.block.mixer.msg\[48\] _1224_ _1225_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_79_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3670__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold651 hotp.block.sha1.mixer.w\[292\] net671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold640 hotp.block.sha1.mixer.w\[348\] net660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold662 hotp.block.sha1.mixer.w\[347\] net682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold673 stream.key_buf\[85\] net693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold695 hotp.block.sha1.mixer.w\[299\] net715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold684 hotp.block.sha1.mixer.b\[20\] net704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2934__I0 hotp.block.mixer.msg\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4176__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2991__S _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4194__D net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3941_ net370 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[168\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_42_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3872_ net738 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[99\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2823_ _1133_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_14_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2754_ hotp.digest\[31\] _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_57_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1705_ stream.key_state\[1\] _1449_ _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2685_ _0990_ _1000_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_100_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1636_ stream.key_counter\[5\] stream.key_counter\[6\] _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_74_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4424_ _0325_ clknet_leaf_70_clk hotp.block.mixer.msg\[136\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4355_ _0256_ clknet_leaf_73_clk hotp.block.mixer.msg\[67\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4199__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3306_ _0047_ clknet_leaf_36_clk stream.msg_buf\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4286_ _0187_ clknet_leaf_96_clk hotp.block.sha1.mixer.a_carry\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3237_ _1377_ _1378_ _1379_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3168_ hotp.block.mixer.msg\[133\] hotp.block.mixer.msg\[134\] _1335_ _1338_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2119_ stream.msg_buf\[34\] stream.msg_buf\[35\] _0561_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3099_ hotp.block.mixer.msg\[103\] hotp.block.mixer.msg\[104\] _1298_ _1299_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold470 hotp.block.sha1.mixer.d\[14\] net490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold481 hotp.block.sha1.mixer.w\[230\] net501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold492 stream.key_buf\[82\] net512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_95_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3911__D net596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2835__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold84_I hotp.block.sha1.mixer.w\[463\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2470_ _1519_ _0825_ _0827_ _1504_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_2_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3909__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4140_ net332 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[367\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4071_ net715 clknet_leaf_41_clk hotp.block.sha1.mixer.w\[298\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3022_ hotp.block.mixer.msg\[70\] hotp.block.mixer.msg\[71\] _1251_ _1255_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_39_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3924_ net152 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[151\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3855_ net263 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[82\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2806_ _1082_ _1119_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3786_ net483 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2737_ hotp.digest\[28\] hotp.digest\[27\] hotp.digest\[29\] _1067_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2668_ _1005_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_hold592_I hotp.block.sha1.mixer.w\[475\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4407_ _0308_ clknet_leaf_62_clk hotp.block.mixer.msg\[119\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2599_ _0883_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4338_ _0239_ clknet_leaf_86_clk hotp.block.mixer.msg\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4269_ net577 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[496\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2136__S _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3242__A2 _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1774__I _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_5_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1970_ _0448_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3640_ net165 clknet_leaf_93_clk hotp.block.sha1.mixer.a\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3571_ _0144_ clknet_leaf_64_clk hotp.digest\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3731__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3816__D net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2522_ _0839_ _0874_ _0877_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2453_ _1521_ hotp.index\[2\] _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2384_ _0606_ _0616_ _0753_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3881__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4123_ net378 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[350\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput2 in[1] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4054_ net53 clknet_leaf_18_clk hotp.block.sha1.mixer.w\[281\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3005_ _1244_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4237__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold605_I hotp.block.sha1.mixer.w\[364\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3907_ net719 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[134\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3838_ net358 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[65\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3769_ net65 clknet_leaf_85_clk hotp.block.sha1.mixer.e\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold47_I hotp.block.sha1.mixer.w\[501\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_109_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_64_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ hotp.block.sha1.mixer.w_fb hotp.block.sha1.mixer.w\[481\] _0432_ _0433_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1884_ _0364_ _0376_ _1535_ _1564_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_4_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3623_ net780 clknet_leaf_76_clk hotp.block.sha1.mixer.a\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3554_ _0131_ clknet_leaf_17_clk stream.counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3485_ net519 clknet_leaf_29_clk stream.key_buf\[137\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2505_ _0861_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2436_ _0794_ _0796_ _0759_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_hold290_I hotp.block.sha1.mixer.w\[439\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold388_I hotp.block.sha1.mixer.w\[476\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2367_ _0634_ _0622_ _0407_ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4106_ net828 clknet_leaf_26_clk hotp.block.sha1.mixer.w\[333\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold555_I hotp.block.sha1.mixer.w\[499\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2298_ stream.digest\[5\] stream.digest\[6\] _0696_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4037_ net427 clknet_leaf_14_clk hotp.block.sha1.mixer.w\[264\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_65_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_74_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_46_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1998__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3270_ _0376_ _0428_ _1399_ _0685_ _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2221_ _0407_ _0633_ _0634_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4197__D net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2152_ _0581_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2083_ _0542_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2985_ _1233_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1936_ _0367_ _0376_ _0372_ _0369_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA_hold303_I hotp.block.sha1.mixer.w\[206\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1867_ _1587_ _1619_ _1623_ _1625_ _1626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xhold811 hotp.block.sha1.mixer.w\[321\] net831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold800 stream.key_buf\[3\] net820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3606_ _0179_ clknet_leaf_44_clk hotp.digest\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1798_ hotp.block.magic.step\[4\] _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_3_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3537_ _0114_ clknet_leaf_14_clk stream.digest\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2968__I _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3468_ net328 clknet_leaf_29_clk stream.key_buf\[120\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3399_ net617 clknet_leaf_51_clk stream.key_buf\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2419_ _0677_ _0775_ _0782_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2469__A3 _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_13_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3914__D net605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3942__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_91_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2770_ _1467_ _1455_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1721_ _1482_ _1483_ seg.digit\[2\] _1484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2989__S _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold107 hotp.block.sha1.mixer.w\[305\] net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_79_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1652_ _1413_ _1422_ stream.key_state\[0\] _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4440_ _0341_ clknet_leaf_91_clk hotp.block.mixer.msg\[152\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_117_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold118 stream.key_buf\[93\] net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold129 hotp.block.sha1.mixer.w\[193\] net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_clkbuf_leaf_1_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4371_ _0272_ clknet_leaf_60_clk hotp.block.mixer.msg\[83\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3824__D net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3322_ _0063_ clknet_leaf_42_clk stream.msg_buf\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3253_ _0468_ _1389_ _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2204_ _0603_ _0617_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3184_ hotp.block.mixer.msg\[140\] hotp.block.mixer.msg\[141\] _1345_ _1347_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2135_ _0571_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_28_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2066_ stream.msg_buf\[11\] stream.msg_buf\[12\] _0530_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2968_ _1223_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_79_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1919_ _1478_ _1476_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2899__S _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2899_ hotp.block.mixer.msg\[17\] hotp.block.mixer.msg\[18\] _1182_ _1185_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold630 stream.key_buf\[34\] net650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_92_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold641 hotp.block.sha1.mixer.e\[15\] net661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold663 hotp.block.sha1.mixer.c\[4\] net683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold652 hotp.block.sha1.mixer.w\[22\] net672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold696 stream.key_buf\[143\] net716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold674 hotp.block.sha1.mixer.w\[380\] net694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold685 hotp.block.sha1.mixer.c\[18\] net705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3909__D net543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2550__A2 _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4270__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3940_ net830 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[167\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3838__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ net485 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[98\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2822_ hotp.digest\[35\] _1122_ _1116_ _1132_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_54_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2753_ _1065_ _1080_ _1081_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1704_ _1402_ _1467_ _1468_ _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2684_ _0841_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1635_ stream.key_counter\[3\] stream.key_counter\[2\] stream.key_counter\[4\] stream.key_counter\[7\]
+ _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_74_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4423_ _0324_ clknet_leaf_70_clk hotp.block.mixer.msg\[135\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4354_ _0255_ clknet_leaf_72_clk hotp.block.mixer.msg\[66\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3305_ _0046_ clknet_leaf_36_clk stream.msg_buf\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold370_I hotp.block.sha1.mixer.w\[191\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4285_ _0186_ clknet_leaf_96_clk hotp.block.sha1.mixer.a_carry\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3236_ _1106_ _0431_ _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3167_ _1337_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2118_ _0562_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3098_ _1287_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2049_ stream.msg_buf\[4\] stream.msg_buf\[5\] _0519_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold471 stream.key_buf\[127\] net491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold460 hotp.block.sha1.mixer.w\[382\] net480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_25_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold482 hotp.block.sha1.mixer.w\[313\] net502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold493 hotp.block.sha1.mixer.a\[14\] net513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_87_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_1_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1877__A4 _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4070_ net732 clknet_leaf_41_clk hotp.block.sha1.mixer.w\[297\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3021_ _1254_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3923_ net798 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[150\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3854_ net32 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[81\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2805_ hotp.digest\[34\] _1118_ _1107_ _1069_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA_hold216_I hotp.block.sha1.mixer.w\[431\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3785_ net297 clknet_leaf_104_clk hotp.block.sha1.mixer.w\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2736_ hotp.digest\[29\] _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2211__A1 _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2667_ _0837_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold585_I hotp.block.sha1.mixer.w\[142\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4406_ _0307_ clknet_leaf_63_clk hotp.block.mixer.msg\[118\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2598_ _0914_ _0943_ _0944_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_hold752_I hotp.block.sha1.mixer.w\[372\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4337_ _0238_ clknet_leaf_92_clk hotp.block.mixer.msg\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4268_ net477 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[495\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3219_ hotp.block.mixer.msg\[155\] hotp.block.mixer.msg\[156\] _1366_ _1367_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_87_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4199_ net542 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[426\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3047__I _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_41_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold290 hotp.block.sha1.mixer.w\[439\] net310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3922__D net620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_56_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4189__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_114_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1965__I _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3570_ _0143_ clknet_leaf_55_clk hotp.digest\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_58_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2521_ hotp.digest\[2\] _0876_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2452_ _1624_ _0809_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2383_ _1448_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3832__D net528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4122_ net204 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[349\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4053_ net437 clknet_leaf_18_clk hotp.block.sha1.mixer.w\[280\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput3 in[2] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3004_ _1159_ _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_69_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3406__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_82_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3906_ net387 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[133\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold500_I hotp.block.sha1.mixer.w\[227\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1875__I _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3837_ net206 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[64\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3768_ net115 clknet_leaf_78_clk hotp.block.sha1.mixer.e\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2719_ _1050_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3699_ net436 clknet_leaf_85_clk hotp.block.sha1.mixer.c\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4331__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output15_I net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3917__D net337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_107_clk clknet_4_2_0_clk clknet_leaf_107_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1952_ _1514_ _0431_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1883_ _0375_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3622_ net188 clknet_leaf_75_clk hotp.block.sha1.mixer.a\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3553_ _0130_ clknet_leaf_16_clk stream.counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_45_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3484_ net556 clknet_leaf_29_clk stream.key_buf\[136\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2504_ _0840_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_102_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2435_ _0795_ _0780_ _0791_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4204__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold283_I hotp.block.sha1.mixer.w\[429\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4105_ net59 clknet_leaf_27_clk hotp.block.sha1.mixer.w\[332\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2366_ _0407_ _0736_ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2297_ _0697_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4036_ net132 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[263\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold715_I hotp.block.sha1.mixer.w\[387\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_111_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3871__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2220_ _0615_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2151_ stream.msg_buf\[48\] stream.msg_buf\[49\] _0577_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2082_ stream.msg_buf\[18\] stream.msg_buf\[19\] _0540_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_66_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2635__A1 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2984_ hotp.block.mixer.msg\[54\] hotp.block.mixer.msg\[55\] _1229_ _1233_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1935_ _0418_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_hold129_I hotp.block.sha1.mixer.w\[193\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1866_ _1568_ _1624_ _1625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3605_ _0178_ clknet_leaf_66_clk hotp.digest\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold801 hotp.block.sha1.mixer.b\[9\] net821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold812 hotp.block.sha1.mixer.b\[7\] net832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1797_ _1555_ _1557_ _1558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_77_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3536_ _0113_ clknet_leaf_14_clk stream.digest\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold498_I hotp.block.sha1.mixer.w\[156\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3467_ net171 clknet_leaf_32_clk stream.key_buf\[119\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold665_I hotp.block.sha1.mixer.w\[71\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3398_ net420 clknet_leaf_51_clk stream.key_buf\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2418_ _0632_ _0613_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2349_ _0726_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4019_ net720 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[246\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3930__D net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2843__B _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2335__S _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1720_ seg.digit\[0\] _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1651_ _1421_ _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold108 hotp.block.sha1.mixer.e\[30\] net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_117_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold119 stream.key_buf\[95\] net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_81_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4370_ _0271_ clknet_leaf_73_clk hotp.block.mixer.msg\[82\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3321_ _0062_ clknet_leaf_41_clk stream.msg_buf\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4001__D net555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3252_ _0469_ _1383_ _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2203_ stream.counter\[12\] stream.counter\[7\] _0605_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input6_I in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3183_ _1346_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2134_ _0514_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2065_ _0532_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold246_I hotp.block.sha1.mixer.w\[385\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2967_ _1160_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_79_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1918_ _0404_ net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2898_ _1184_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1849_ hotp.block.main_in _1607_ _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold782_I hotp.block.sha1.mixer.w\[109\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold620 hotp.block.sha1.mixer.e\[25\] net640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold631 stream.key_buf\[114\] net651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold642 stream.key_buf\[57\] net662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold653 stream.key_buf\[32\] net673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold697 stream.key_buf\[30\] net717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold664 stream.key_buf\[154\] net684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold686 hotp.block.sha1.mixer.w\[108\] net706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold675 hotp.block.sha1.mixer.w\[411\] net695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3519_ _0096_ clknet_leaf_98_clk stream.digest\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_96_clk clknet_4_9_0_clk clknet_leaf_96_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_20_clk clknet_4_4_0_clk clknet_leaf_20_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3925__D net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_87_clk clknet_4_8_0_clk clknet_leaf_87_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2838__A1 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3870_ net760 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[97\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2821_ hotp.digest\[34\] _1126_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2752_ _1066_ _1058_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_11_clk clknet_4_1_0_clk clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1703_ stream.key_state\[0\] stream.key_state\[2\] _1429_ _1468_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2683_ hotp.digest\[23\] _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4422_ _0323_ clknet_leaf_70_clk hotp.block.mixer.msg\[134\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3835__D net486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1634_ stream.key_state\[3\] _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_74_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4353_ _0254_ clknet_leaf_72_clk hotp.block.mixer.msg\[65\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3304_ _0045_ clknet_leaf_36_clk stream.msg_buf\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4284_ _0012_ clknet_leaf_97_clk hotp.block.sha1.mixer.w\[511\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3235_ _1106_ _0430_ _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_78_clk clknet_4_10_0_clk clknet_leaf_78_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4095__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3166_ hotp.block.mixer.msg\[132\] hotp.block.mixer.msg\[133\] _1335_ _1337_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2117_ stream.msg_buf\[33\] stream.msg_buf\[34\] _0561_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3097_ _1297_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2048_ _0522_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3999_ net520 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[226\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3932__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold450 stream.key_buf\[71\] net470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold461 hotp.block.sha1.mixer.w\[148\] net481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold472 hotp.block.sha1.mixer.w\[184\] net492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold494 stream.key_buf\[87\] net514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold483 hotp.block.sha1.mixer.w\[91\] net503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xclkbuf_leaf_69_clk clknet_4_11_0_clk clknet_leaf_69_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1788__I _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3245__A1 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0_clk clknet_4_0_0_clk clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3020_ hotp.block.mixer.msg\[69\] hotp.block.mixer.msg\[70\] _1251_ _1254_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3236__A1 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ net620 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[149\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3853_ net598 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[80\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2804_ _1117_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3784_ net201 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2735_ _1005_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2666_ _0973_ _1003_ _1004_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4405_ _0306_ clknet_leaf_63_clk hotp.block.mixer.msg\[117\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2597_ _0930_ _0937_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4336_ _0237_ clknet_leaf_90_clk hotp.block.mixer.msg\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold578_I hotp.block.sha1.mixer.w\[81\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3153__I _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4267_ net631 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[494\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3218_ _1350_ _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4198_ net434 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[425\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3149_ hotp.block.mixer.msg\[125\] hotp.block.mixer.msg\[126\] _1324_ _1327_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3002__I1 hotp.block.mixer.msg\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3828__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold280 hotp.block.sha1.mixer.w\[1\] net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold291 hotp.block.sha1.mixer.w\[120\] net311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3358__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2520_ _0875_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2451_ hotp.index\[1\] _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2382_ _0626_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4121_ net233 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[348\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4052_ net779 clknet_leaf_18_clk hotp.block.sha1.mixer.w\[279\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput4 in[3] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3003_ _1243_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_69_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold159_I hotp.block.sha1.mixer.w\[211\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3905_ net416 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[132\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3836_ net157 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3767_ net274 clknet_leaf_84_clk hotp.block.sha1.mixer.e\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2718_ hotp.digest\[27\] _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3698_ net708 clknet_leaf_85_clk hotp.block.sha1.mixer.c\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2649_ _0973_ _0988_ _0989_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4319_ _0220_ clknet_leaf_90_clk hotp.block.mixer.msg\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3933__D net369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1951_ _0430_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1882_ _1568_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3621_ net450 clknet_leaf_75_clk hotp.block.sha1.mixer.a\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3552_ _0129_ clknet_leaf_16_clk stream.counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4004__D net613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2503_ _0859_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3483_ net701 clknet_leaf_29_clk stream.key_buf\[135\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3843__D net685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2434_ _0610_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2365_ _0624_ _1416_ _0632_ _0615_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4104_ net793 clknet_leaf_27_clk hotp.block.sha1.mixer.w\[331\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2296_ stream.digest\[4\] stream.digest\[5\] _0696_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ net366 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[262\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_40_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3673__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3819_ net809 clknet_leaf_107_clk hotp.block.sha1.mixer.w\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_55_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4179__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_113_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1796__I _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3928__D net518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold52_I hotp.block.sha1.mixer.w\[460\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2150_ _0580_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2081_ _0541_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2983_ _1232_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3838__D net358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1934_ _1549_ _0417_ _1514_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1865_ hotp.block.magic.step\[4\] _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold802 stream.key_buf\[6\] net822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3604_ _0177_ clknet_leaf_66_clk hotp.index\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1796_ _1556_ _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_77_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1655__B _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3535_ _0112_ clknet_leaf_18_clk stream.digest\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold813 hotp.block.sha1.mixer.e\[11\] net833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3466_ net602 clknet_leaf_32_clk stream.key_buf\[118\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2417_ _0677_ _0775_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3397_ net377 clknet_leaf_51_clk stream.key_buf\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2348_ stream.digest\[27\] stream.digest\[28\] _0722_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold658_I hotp.block.sha1.mixer.w\[246\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2279_ _0684_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4018_ net678 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[245\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1650_ _1420_ _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2351__S _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold109 hotp.block.sha1.mixer.w\[315\] net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_81_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3320_ _0061_ clknet_leaf_41_clk stream.msg_buf\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3251_ _0469_ _1383_ _1388_ _1380_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2202_ stream.counter\[1\] stream.counter\[0\] _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3182_ hotp.block.mixer.msg\[139\] hotp.block.mixer.msg\[140\] _1345_ _1346_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2133_ _0570_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2064_ stream.msg_buf\[10\] stream.msg_buf\[11\] _0530_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold141_I hotp.block.sha1.mixer.w\[231\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2966_ _1222_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_79_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1917_ _1581_ _0403_ _1476_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2897_ hotp.block.mixer.msg\[16\] hotp.block.mixer.msg\[17\] _1182_ _1184_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1848_ _1606_ _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold610 stream.key_buf\[76\] net630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold621 hotp.block.sha1.mixer.w\[160\] net641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold654 stream.key_buf\[131\] net674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold632 stream.key_buf\[140\] net652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_hold775_I hotp.block.sha1.mixer.w\[260\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold643 hotp.block.sha1.mixer.w\[154\] net663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1779_ _1537_ _1539_ _1540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold665 hotp.block.sha1.mixer.w\[71\] net685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold676 hotp.block.sha1.mixer.w\[92\] net696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold687 hotp.block.sha1.mixer.d\[23\] net707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3518_ _0095_ clknet_leaf_99_clk stream.digest\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3449_ net324 clknet_leaf_30_clk stream.key_buf\[101\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold698 hotp.block.sha1.mixer.w\[441\] net718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2995__I _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4217__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3941__D net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2138__I1 stream.msg_buf\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2346__S _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2820_ _1126_ _1130_ _1131_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_14_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2751_ _1076_ _0862_ _1077_ _1079_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3734__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1702_ _1424_ _1467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2682_ _1006_ _1017_ _1018_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1633_ stream.key_state\[2\] _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4421_ _0322_ clknet_leaf_70_clk hotp.block.mixer.msg\[133\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4012__D net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3884__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4352_ _0253_ clknet_leaf_72_clk hotp.block.mixer.msg\[64\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3303_ _0044_ clknet_leaf_36_clk stream.msg_buf\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3851__D net548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4283_ net254 clknet_leaf_96_clk hotp.block.sha1.mixer.w\[510\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3234_ _0684_ _1376_ _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3165_ _1336_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2116_ _0550_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3096_ hotp.block.mixer.msg\[102\] hotp.block.mixer.msg\[103\] _1293_ _1297_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2047_ stream.msg_buf\[3\] stream.msg_buf\[4\] _0519_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold523_I hotp.block.sha1.mixer.w\[137\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3998_ net234 clknet_leaf_114_clk hotp.block.sha1.mixer.w\[225\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2949_ _1202_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_45_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold462 hotp.block.sha1.mixer.w\[262\] net482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold440 hotp.block.sha1.mixer.w\[31\] net460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold451 hotp.block.sha1.mixer.b\[13\] net471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold473 hotp.block.sha1.mixer.w\[267\] net493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold495 hotp.block.sha1.mixer.c\[15\] net515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold484 hotp.block.sha1.mixer.w\[6\] net504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3936__D net805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3921_ net766 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[148\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4007__D net530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3852_ net110 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[79\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2803_ hotp.digest\[31\] hotp.digest\[32\] hotp.digest\[33\] _1117_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3783_ net131 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3846__D net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2734_ _1035_ _1063_ _1064_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2665_ _0990_ _0998_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2596_ _0939_ _0940_ _0942_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4404_ _0305_ clknet_leaf_63_clk hotp.block.mixer.msg\[116\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4335_ _0236_ clknet_leaf_88_clk hotp.block.mixer.msg\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4266_ net740 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[493\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3217_ _1365_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4197_ net136 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[424\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3148_ _1326_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3079_ _1244_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold270 hotp.block.sha1.mixer.w\[464\] net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold281 stream.key_buf\[94\] net301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold292 hotp.block.sha1.mixer.w\[341\] net312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_102_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold82_I hotp.block.sha1.mixer.w\[170\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2450_ _1568_ hotp.index\[0\] hotp.index\[1\] _1624_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_20_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2381_ _1448_ _0750_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4120_ net660 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[347\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4051_ net294 clknet_leaf_17_clk hotp.block.sha1.mixer.w\[278\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3922__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 in[4] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3002_ hotp.block.mixer.msg\[62\] hotp.block.mixer.msg\[63\] _1239_ _1243_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_69_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3904_ net309 clknet_leaf_25_clk hotp.block.sha1.mixer.w\[131\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold319_I hotp.block.sha1.mixer.w\[465\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold221_I hotp.block.sha1.mixer.w\[186\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3835_ net486 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_43_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3766_ net166 clknet_leaf_78_clk hotp.block.sha1.mixer.e\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2717_ _1035_ _1048_ _1049_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3697_ net173 clknet_leaf_84_clk hotp.block.sha1.mixer.c\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2648_ hotp.digest\[17\] _0966_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2579_ hotp.digest\[10\] _0898_ _0927_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4200__D net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4318_ _0219_ clknet_leaf_91_clk hotp.block.mixer.msg\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4249_ net827 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[476\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2671__C _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2243__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1950_ _0428_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1881_ _0371_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3620_ net774 clknet_leaf_75_clk hotp.block.sha1.mixer.a\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3551_ _0128_ clknet_leaf_17_clk stream.counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2502_ _0840_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3482_ net94 clknet_leaf_28_clk stream.key_buf\[134\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2433_ _0749_ _0792_ _0610_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2364_ _1442_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4020__D net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4103_ net194 clknet_leaf_26_clk hotp.block.sha1.mixer.w\[330\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_16_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2295_ _0690_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4034_ net482 clknet_leaf_15_clk hotp.block.sha1.mixer.w\[261\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold269_I hotp.block.sha1.mixer.w\[146\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold603_I hotp.block.sha1.mixer.w\[389\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3818_ net109 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3749_ net29 clknet_leaf_75_clk hotp.block.sha1.mixer.e\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_104_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_43_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3944__D net786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2080_ stream.msg_buf\[17\] stream.msg_buf\[18\] _0540_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4273__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_61_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2982_ hotp.block.mixer.msg\[53\] hotp.block.mixer.msg\[54\] _1229_ _1232_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_83_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1933_ _1517_ _1518_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4015__D net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3603_ _0176_ clknet_leaf_66_clk hotp.index\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1864_ _1610_ _1621_ _1622_ _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold803 hotp.block.sha1.mixer.w\[388\] net823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3854__D net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1795_ _1547_ _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3534_ _0111_ clknet_leaf_17_clk stream.digest\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2020__A1 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold814 hotp.block.sha1.mixer.w\[256\] net834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3465_ net494 clknet_leaf_32_clk stream.key_buf\[117\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2416_ _0736_ _0738_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3396_ net348 clknet_leaf_51_clk stream.key_buf\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2347_ _0725_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2278_ hotp.rst_n _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_hold553_I hotp.block.sha1.mixer.w\[467\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4017_ net608 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[244\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3640__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2011__A1 _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_106_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3939__D net535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1761__B1 _1520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3250_ _1528_ _1386_ _0819_ _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2201_ _1414_ _0508_ stream.debug\[1\] _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3181_ _1329_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2132_ stream.msg_buf\[40\] stream.msg_buf\[41\] _0566_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _0531_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_54_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3849__D net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2965_ hotp.block.mixer.msg\[46\] hotp.block.mixer.msg\[47\] _1218_ _1222_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_69_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1916_ hotp.digest\[0\] _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold301_I hotp.block.sha1.mixer.w\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2896_ _1183_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1847_ _1604_ _1605_ _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_112_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold600 hotp.block.sha1.mixer.w\[150\] net620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold611 hotp.block.sha1.mixer.w\[495\] net631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold644 stream.key_buf\[73\] net664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold622 stream.key_buf\[47\] net642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold633 stream.key_buf\[48\] net653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1778_ hotp.block.mixer.round\[0\] _1530_ _1538_ _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3517_ _0094_ clknet_leaf_99_clk stream.digest\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold677 hotp.block.sha1.mixer.w\[127\] net697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold666 stream.key_buf\[148\] net686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_69_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold688 hotp.block.sha1.mixer.c\[22\] net708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold655 hotp.block.sha1.mixer.w\[24\] net675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3448_ net817 clknet_leaf_30_clk stream.key_buf\[100\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold699 hotp.block.sha1.mixer.w\[135\] net719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_hold768_I hotp.block.sha1.mixer.w\[238\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3379_ net673 clknet_leaf_56_clk stream.key_buf\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3172__I _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2251__I _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2750_ _0980_ _1078_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1701_ _1463_ _1466_ _1443_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2681_ hotp.digest\[21\] _0998_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1632_ stream.key_state\[1\] _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4420_ _0321_ clknet_leaf_70_clk hotp.block.mixer.msg\[132\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4351_ _0252_ clknet_leaf_70_clk hotp.block.mixer.msg\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3302_ _0043_ clknet_leaf_36_clk stream.msg_buf\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4282_ net75 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[509\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3233_ hotp.stage\[2\] _1606_ _1375_ _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3164_ hotp.block.mixer.msg\[131\] hotp.block.mixer.msg\[132\] _1335_ _1336_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2115_ _0560_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3095_ _1296_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2046_ _0521_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold251_I hotp.block.sha1.mixer.w\[87\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold349_I hotp.block.sha1.mixer.w\[161\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3997_ net141 clknet_leaf_113_clk hotp.block.sha1.mixer.w\[224\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2948_ _1212_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2879_ _1173_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4203__D net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold441 hotp.block.sha1.mixer.w\[254\] net461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold452 hotp.block.sha1.mixer.d\[22\] net472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold430 hotp.block.sha1.mixer.a\[9\] net450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold463 hotp.block.sha1.mixer.w\[14\] net483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold474 stream.key_buf\[118\] net494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold496 hotp.block.sha1.mixer.w\[322\] net516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_8_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold485 hotp.block.sha1.mixer.c\[26\] net505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2246__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2910__S _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3952__D net522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2357__S _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3920_ net481 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[147\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3851_ net548 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[78\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2802_ _1115_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3851__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3782_ net125 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2733_ _1051_ _1058_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4023__D net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2664_ _1000_ _0985_ _1002_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4207__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2595_ _0909_ _0941_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4403_ _0304_ clknet_leaf_57_clk hotp.block.mixer.msg\[115\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3862__D net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4334_ _0235_ clknet_leaf_90_clk hotp.block.mixer.msg\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4265_ net495 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[492\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold466_I hotp.block.sha1.mixer.w\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3216_ hotp.block.mixer.msg\[154\] hotp.block.mixer.msg\[155\] _1361_ _1365_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4196_ net267 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[423\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3147_ hotp.block.mixer.msg\[124\] hotp.block.mixer.msg\[125\] _1324_ _1326_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3078_ _1286_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2029_ _0506_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_108_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2015__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold260 hotp.block.sha1.mixer.c\[24\] net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold271 hotp.block.sha1.mixer.w\[488\] net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold293 hotp.block.sha1.mixer.w\[296\] net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold282 hotp.block.sha1.mixer.w\[182\] net302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3874__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3947__D net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold75_I hotp.block.sha1.mixer.w\[358\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2380_ _0745_ _0749_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4050_ net42 clknet_leaf_18_clk hotp.block.sha1.mixer.w\[277\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput6 in[5] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3001_ _1242_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4018__D net678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3903_ net164 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[130\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3857__D net402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3834_ net37 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_43_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold214_I hotp.block.sha1.mixer.w\[226\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_89_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3765_ net640 clknet_leaf_78_clk hotp.block.sha1.mixer.e\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2716_ hotp.digest\[25\] _1027_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3696_ net229 clknet_leaf_83_clk hotp.block.sha1.mixer.c\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2647_ hotp.digest\[18\] _0985_ _0987_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold583_I hotp.block.sha1.mixer.w\[408\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2578_ _0909_ _0926_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4317_ _0218_ clknet_leaf_104_clk hotp.block.mixer.msg\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4248_ net408 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[475\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold750_I hotp.block.sha1.mixer.w\[378\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_98_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4179_ net394 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[406\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_109_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_64_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1880_ _0366_ _0370_ _1623_ _1587_ _0372_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_36_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3550_ _0127_ clknet_leaf_19_clk stream.counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2501_ _0839_ _0854_ _0858_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3481_ net287 clknet_leaf_33_clk stream.key_buf\[133\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2432_ _0611_ _0790_ _0793_ _0646_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2363_ _0732_ _0733_ _0734_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4102_ net54 clknet_leaf_27_clk hotp.block.sha1.mixer.w\[329\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2294_ _0695_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4033_ net158 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[260\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3817_ net781 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3748_ net540 clknet_leaf_75_clk hotp.block.sha1.mixer.e\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4211__D net310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3679_ net219 clknet_leaf_79_clk hotp.block.sha1.mixer.c\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output13_I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_50_clk clknet_4_13_0_clk clknet_leaf_50_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3912__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3960__D net409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2981_ _1231_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_41_clk clknet_4_6_0_clk clknet_leaf_41_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1932_ hotp.block.sha1.mixer.b\[0\] _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1863_ _1604_ _1552_ _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3602_ _0175_ clknet_leaf_65_clk hotp.index\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1794_ _1554_ _1555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3533_ _0110_ clknet_leaf_17_clk stream.digest\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold815 hotp.block.sha1.mixer.w\[375\] net835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold804 hotp.block.sha1.mixer.w\[162\] net824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4031__D net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3464_ net571 clknet_leaf_32_clk stream.key_buf\[116\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2415_ _0779_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3870__D net760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3395_ net653 clknet_leaf_51_clk stream.key_buf\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4098__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2346_ stream.digest\[26\] stream.digest\[27\] _0722_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2277_ _0675_ _0682_ _0683_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4016_ net819 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[243\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold713_I hotp.block.sha1.mixer.w\[366\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3935__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_32_clk clknet_4_5_0_clk clknet_leaf_32_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4206__D net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold8_I hotp.block.sha1.mixer.w\[73\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_99_clk clknet_4_3_0_clk clknet_leaf_99_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_23_clk clknet_4_4_0_clk clknet_leaf_23_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_61_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3955__D net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4240__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2200_ stream.debug\[1\] _1445_ _0509_ _0613_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3180_ _1344_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2131_ _0569_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2062_ stream.msg_buf\[9\] stream.msg_buf\[10\] _0530_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2964_ _1221_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4026__D net461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1915_ _1482_ _1477_ _0402_ net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xclkbuf_leaf_14_clk clknet_4_3_0_clk clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_79_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2895_ hotp.block.mixer.msg\[15\] hotp.block.mixer.msg\[16\] _1182_ _1183_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3865__D net771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ _1495_ _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1777_ _1507_ _1523_ _1502_ _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_8_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold612 hotp.block.sha1.mixer.w\[33\] net632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold601 hotp.block.sha1.mixer.w\[68\] net621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold623 stream.key_buf\[65\] net643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_102_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold634 hotp.block.sha1.mixer.e\[7\] net654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold645 hotp.block.sha1.mixer.b\[23\] net665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3516_ _0093_ clknet_leaf_99_clk stream.digest\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold667 stream.key_buf\[38\] net687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1682__B net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold678 hotp.block.sha1.mixer.w\[37\] net698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold656 hotp.block.sha1.mixer.e\[20\] net676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3447_ net639 clknet_leaf_30_clk stream.key_buf\[99\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3488__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold689 stream.key_buf\[151\] net709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3378_ net441 clknet_leaf_56_clk stream.key_buf\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2329_ _0715_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3257__A1 _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_36_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_80_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4263__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1991__A1 _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2908__S _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1700_ stream.msg_state\[3\] _1465_ _1466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2680_ hotp.digest\[22\] _0985_ _1016_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1631_ _1401_ _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4350_ _0251_ clknet_leaf_84_clk hotp.block.mixer.msg\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3301_ _0042_ clknet_leaf_36_clk stream.msg_buf\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4281_ net463 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[508\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3232_ _0468_ _1525_ _0430_ _1374_ _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
Xclkbuf_leaf_3_clk clknet_4_0_0_clk clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3163_ _1329_ _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2114_ stream.msg_buf\[32\] stream.msg_buf\[33\] _0556_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3094_ hotp.block.mixer.msg\[101\] hotp.block.mixer.msg\[102\] _1293_ _1296_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2045_ stream.msg_buf\[2\] stream.msg_buf\[3\] _0519_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4136__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold244_I hotp.block.sha1.mixer.w\[158\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3996_ net307 clknet_leaf_114_clk hotp.block.sha1.mixer.w\[223\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2947_ hotp.block.mixer.msg\[38\] hotp.block.mixer.msg\[39\] _1208_ _1212_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold509_I hotp.block.sha1.mixer.w\[468\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2878_ hotp.block.mixer.msg\[8\] hotp.block.mixer.msg\[9\] _1171_ _1173_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold420 stream.key_buf\[128\] net440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1829_ _1588_ _1589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold442 stream.key_buf\[69\] net462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold453 stream.key_buf\[78\] net473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold431 hotp.block.sha1.mixer.w\[94\] net451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_96_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold486 hotp.block.sha1.mixer.w\[374\] net506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold464 hotp.block.sha1.mixer.w\[204\] net484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold475 hotp.block.sha1.mixer.w\[493\] net495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold497 stream.key_buf\[39\] net517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_109_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_11_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_53_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_118_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_68_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_111_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3850_ net299 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[77\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2801_ _0830_ _0855_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3781_ net336 clknet_leaf_100_clk hotp.block.sha1.mixer.w\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2732_ _1060_ _0842_ _1062_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2663_ _0991_ _1001_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2594_ hotp.digest\[10\] _0933_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4402_ _0303_ clknet_leaf_58_clk hotp.block.mixer.msg\[114\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4333_ _0234_ clknet_leaf_89_clk hotp.block.mixer.msg\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4264_ net359 clknet_leaf_100_clk hotp.block.sha1.mixer.w\[491\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3215_ _1364_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4195_ net525 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[422\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3146_ _1325_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold459_I hotp.block.sha1.mixer.w\[437\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3077_ hotp.block.mixer.msg\[94\] hotp.block.mixer.msg\[95\] _1282_ _1286_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2028_ _1427_ _1438_ _0505_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_hold626_I hotp.block.sha1.mixer.w\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3676__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4214__D net691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3979_ net713 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[206\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold261 hotp.block.sha1.mixer.e\[13\] net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold250 hotp.block.sha1.mixer.w\[54\] net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold283 hotp.block.sha1.mixer.w\[429\] net303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold294 hotp.block.sha1.mixer.b\[15\] net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold272 hotp.block.sha1.mixer.w\[482\] net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4451__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3963__D net390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput7 in[6] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3000_ hotp.block.mixer.msg\[61\] hotp.block.mixer.msg\[62\] _1239_ _1242_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_69_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3902_ net773 clknet_leaf_25_clk hotp.block.sha1.mixer.w\[129\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3833_ net321 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3764_ net286 clknet_leaf_79_clk hotp.block.sha1.mixer.e\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2715_ hotp.digest\[26\] _1020_ _1047_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3873__D net591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3695_ net58 clknet_leaf_86_clk hotp.block.sha1.mixer.c\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2646_ _0954_ _0986_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2577_ _0908_ _0921_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_77_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold576_I hotp.block.sha1.mixer.w\[139\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4316_ _0217_ clknet_leaf_104_clk hotp.block.mixer.msg\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4247_ net612 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[474\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4178_ net570 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[405\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4209__D net479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3129_ hotp.block.mixer.msg\[116\] hotp.block.mixer.msg\[117\] _1314_ _1316_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_2_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3841__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3958__D net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3480_ net611 clknet_leaf_33_clk stream.key_buf\[132\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2500_ _0403_ _0857_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2431_ stream.counter\[9\] _0749_ _0782_ _0792_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2362_ _0431_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4101_ net81 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[328\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2293_ stream.digest\[3\] stream.digest\[4\] _0691_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4032_ net795 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[259\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4029__D net363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold157_I hotp.block.sha1.mixer.w\[103\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3868__D net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3816_ net276 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3747_ net654 clknet_leaf_75_clk hotp.block.sha1.mixer.e\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_95_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold693_I hotp.block.sha1.mixer.w\[207\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3678_ net87 clknet_leaf_85_clk hotp.block.sha1.mixer.c\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2629_ _0959_ _0966_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_7_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3394__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_66_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2980_ hotp.block.mixer.msg\[52\] hotp.block.mixer.msg\[53\] _1229_ _1231_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1931_ _0412_ _0415_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3737__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1862_ _1620_ _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3601_ _0174_ clknet_leaf_65_clk hotp.index\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1793_ hotp.block.magic.step\[1\] _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3532_ _0109_ clknet_leaf_17_clk stream.digest\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold805 hotp.block.sha1.mixer.a\[4\] net825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold816 hotp.block.sha1.mixer.w\[190\] net836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3463_ net184 clknet_leaf_31_clk stream.key_buf\[115\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2414_ _0604_ _0774_ _0778_ _1425_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_58_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3394_ net642 clknet_leaf_51_clk stream.key_buf\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2345_ _0724_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2276_ hotp.block.main_in _0675_ _1467_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4015_ net24 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[242\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold441_I hotp.block.sha1.mixer.w\[254\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold539_I hotp.block.sha1.mixer.w\[67\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4222__D net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4192__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4132__D net599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3971__D net680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2130_ stream.msg_buf\[39\] stream.msg_buf\[40\] _0566_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2061_ _0529_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2963_ hotp.block.mixer.msg\[45\] hotp.block.mixer.msg\[46\] _1218_ _1221_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1914_ stream.debug\[1\] _1602_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2894_ _1181_ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_72_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1845_ hotp.block.mixer.stage\[1\] _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1776_ _1536_ _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold602 hotp.block.sha1.mixer.w\[365\] net622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_4_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold635 hotp.block.sha1.mixer.w\[126\] net655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3881__D net802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold613 hotp.block.sha1.mixer.w\[445\] net633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold624 hotp.block.sha1.mixer.d\[4\] net644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3515_ _0092_ clknet_leaf_99_clk stream.digest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold657 stream.key_buf\[53\] net677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold646 hotp.block.sha1.mixer.w\[455\] net666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold668 hotp.block.sha1.mixer.w\[212\] net688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold391_I hotp.block.sha1.mixer.w\[214\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold679 hotp.block.sha1.mixer.w\[8\] net699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3446_ net439 clknet_leaf_30_clk stream.key_buf\[98\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3377_ net717 clknet_leaf_56_clk stream.key_buf\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2328_ stream.digest\[18\] stream.digest\[19\] _0712_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2259_ _0652_ _0667_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4217__D net633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_112_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3966__D net424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1630_ net2 _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1982__A2 _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3300_ _0041_ clknet_leaf_40_clk stream.msg_buf\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ net191 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[507\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3231_ _0819_ _0826_ _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3162_ _1334_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2113_ _0559_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3093_ _1295_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2044_ _0520_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_85_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold237_I hotp.block.sha1.mixer.w\[74\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3876__D net553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3995_ net422 clknet_leaf_114_clk hotp.block.sha1.mixer.w\[222\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2946_ _1211_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold404_I hotp.block.sha1.mixer.w\[194\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2877_ _1172_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ _1587_ _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold410 hotp.block.sha1.mixer.w\[205\] net430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold421 stream.key_buf\[31\] net441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold432 hotp.block.sha1.mixer.w\[448\] net452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1759_ hotp.block.mixer.msg\[64\] hotp.block.mixer.msg\[96\] _1498_ _1520_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold443 hotp.block.sha1.mixer.w\[509\] net463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold454 hotp.block.sha1.mixer.w\[57\] net474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold773_I hotp.block.sha1.mixer.w\[332\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold487 hotp.block.sha1.mixer.w\[138\] net507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold465 hotp.block.sha1.mixer.w\[99\] net485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold476 hotp.block.sha1.mixer.a\[19\] net496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3429_ net512 clknet_leaf_35_clk stream.key_buf\[81\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold498 hotp.block.sha1.mixer.w\[156\] net518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__1712__I hotp.block.debug\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3948__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_19_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2800_ _1593_ _1110_ _1114_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_30_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3780_ net699 clknet_leaf_100_clk hotp.block.sha1.mixer.w\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2731_ _1030_ _1061_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4401_ _0302_ clknet_leaf_58_clk hotp.block.mixer.msg\[113\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2662_ hotp.digest\[18\] _0994_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2593_ _0859_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4332_ _0233_ clknet_leaf_89_clk hotp.block.mixer.msg\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4263_ net120 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[490\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3214_ hotp.block.mixer.msg\[153\] hotp.block.mixer.msg\[154\] _1361_ _1364_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4194_ net140 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[421\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_87_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3145_ hotp.block.mixer.msg\[123\] hotp.block.mixer.msg\[124\] _1324_ _1325_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3076_ _1285_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold354_I hotp.block.sha1.mixer.w\[219\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2027_ stream.msg_state\[3\] _1472_ stream.msg_state\[2\] _0505_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3978_ net323 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[205\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2929_ _1201_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_98_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold262 stream.key_buf\[96\] net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4230__D net338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold251 hotp.block.sha1.mixer.w\[87\] net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold240 hotp.block.sha1.mixer.w\[52\] net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_102_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold284 stream.key_buf\[44\] net304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold295 hotp.block.sha1.mixer.w\[403\] net315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold273 hotp.block.sha1.mixer.w\[90\] net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_102_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1937__A2 _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4140__D net332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4276__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 rst_n net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_69_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3901_ net763 clknet_leaf_25_clk hotp.block.sha1.mixer.w\[128\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3832_ net528 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3763_ net426 clknet_leaf_79_clk hotp.block.sha1.mixer.e\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2714_ _1030_ _1046_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3694_ net705 clknet_leaf_87_clk hotp.block.sha1.mixer.c\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2645_ _0968_ _0979_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_100_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2576_ _0914_ _0924_ _0925_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4315_ _0216_ clknet_leaf_104_clk hotp.block.mixer.msg\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4246_ net60 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[473\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4177_ net433 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[404\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3128_ _1315_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3643__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3059_ hotp.block.mixer.msg\[86\] hotp.block.mixer.msg\[87\] _1272_ _1276_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_52_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_67_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_110_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4135__D net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold80_I hotp.block.sha1.mixer.w\[367\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3974__D net746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2430_ _0738_ _0791_ _0737_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2361_ hotp.block.sha1.mixer.e\[0\] _1591_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4100_ net78 clknet_leaf_27_clk hotp.block.sha1.mixer.w\[327\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2292_ _0694_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4031_ net41 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[258\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold317_I hotp.block.sha1.mixer.w\[145\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3815_ net627 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3746_ net837 clknet_leaf_77_clk hotp.block.sha1.mixer.e\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_95_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2574__A2 _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3677_ net160 clknet_leaf_84_clk hotp.block.sha1.mixer.c\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold686_I hotp.block.sha1.mixer.w\[108\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2628_ _0968_ _0940_ _0970_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2559_ hotp.digest\[6\] _0902_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4229_ net172 clknet_leaf_14_clk hotp.block.sha1.mixer.w\[456\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_21_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3969__D net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1630__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1930_ _1402_ _0413_ net1 _0414_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_29_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1861_ _1545_ _1620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3600_ _0173_ clknet_leaf_46_clk stream.key_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3531_ _0108_ clknet_leaf_17_clk stream.digest\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1792_ _1552_ _1543_ _1553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold806 stream.key_buf\[15\] net826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold817 hotp.block.sha1.mixer.e\[6\] net837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3462_ net794 clknet_leaf_31_clk stream.key_buf\[114\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3393_ net223 clknet_leaf_49_clk stream.key_buf\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2413_ _1426_ _0775_ _0777_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_90_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2344_ stream.digest\[25\] stream.digest\[26\] _0722_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2275_ stream.msg_buf\[0\] _0650_ _0681_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3879__D net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4014_ net711 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[241\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3241__B _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold601_I hotp.block.sha1.mixer.w\[68\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3831__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3729_ net581 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_100_clk clknet_4_3_0_clk clknet_leaf_100_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_72_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2060_ _0515_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2962_ _1220_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3854__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1913_ _0400_ _1477_ _0401_ net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_45_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2893_ _1160_ _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1844_ _1582_ _1597_ _1487_ _1603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1775_ hotp.block.magic.step\[3\] _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_13_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold603 hotp.block.sha1.mixer.w\[389\] net623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold625 hotp.block.sha1.mixer.w\[304\] net645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold614 hotp.block.sha1.mixer.w\[106\] net634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_69_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold636 hotp.block.sha1.mixer.w\[4\] net656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3514_ _0091_ clknet_leaf_98_clk stream.digest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold669 stream.key_buf\[86\] net689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3445_ net681 clknet_leaf_30_clk stream.key_buf\[97\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold647 hotp.block.sha1.mixer.d\[12\] net667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold658 hotp.block.sha1.mixer.w\[246\] net678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3376_ net22 clknet_leaf_55_clk stream.key_buf\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2327_ _0714_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2258_ stream.digest\[18\] stream.digest\[22\] stream.digest\[26\] stream.digest\[30\]
+ _0653_ _0654_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2189_ stream.counter\[11\] _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold816_I hotp.block.sha1.mixer.w\[190\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4233__D net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3727__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4143__D net649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3982__D net601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3230_ _1593_ _0434_ _1373_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3161_ hotp.block.mixer.msg\[130\] hotp.block.mixer.msg\[131\] _1330_ _1334_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2112_ stream.msg_buf\[31\] stream.msg_buf\[32\] _0556_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3092_ hotp.block.mixer.msg\[100\] hotp.block.mixer.msg\[101\] _1293_ _1295_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2043_ stream.msg_buf\[1\] stream.msg_buf\[2\] _0519_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold132_I hotp.block.sha1.mixer.w\[152\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3994_ net714 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[221\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2945_ hotp.block.mixer.msg\[37\] hotp.block.mixer.msg\[38\] _1208_ _1211_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2876_ hotp.block.mixer.msg\[7\] hotp.block.mixer.msg\[8\] _1171_ _1172_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1827_ _1495_ _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold400 stream.key_buf\[51\] net420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold411 hotp.block.sha1.mixer.c\[16\] net431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold433 stream.key_buf\[126\] net453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1758_ _1496_ _1498_ _1519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold444 hotp.block.sha1.mixer.c\[14\] net464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold422 hotp.block.sha1.mixer.d\[6\] net442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1689_ _1401_ _1410_ _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold477 hotp.block.sha1.mixer.w\[459\] net497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold466 hotp.block.sha1.mixer.w\[63\] net486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold455 hotp.block.sha1.mixer.w\[155\] net475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3428_ net247 clknet_leaf_36_clk stream.key_buf\[80\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold499 stream.key_buf\[138\] net519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold488 hotp.block.sha1.mixer.w\[354\] net508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_hold766_I hotp.block.sha1.mixer.w\[172\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3359_ net317 clknet_leaf_50_clk stream.key_buf\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4138__D net733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3977__D net430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2730_ hotp.digest\[26\] _1054_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2661_ hotp.digest\[20\] _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4400_ _0301_ clknet_leaf_63_clk hotp.block.mixer.msg\[112\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2592_ hotp.digest\[12\] _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ _0232_ clknet_leaf_88_clk hotp.block.mixer.msg\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4262_ net710 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[489\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3213_ _1363_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4193_ net797 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[420\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3144_ _1308_ _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_87_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3075_ hotp.block.mixer.msg\[93\] hotp.block.mixer.msg\[94\] _1282_ _1285_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2026_ _1595_ _0434_ _0504_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2140__I0 stream.msg_buf\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_hold514_I hotp.block.sha1.mixer.w\[419\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3977_ net430 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[204\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2928_ hotp.block.mixer.msg\[30\] hotp.block.mixer.msg\[31\] _1197_ _1201_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2859_ _1161_ _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold230 hotp.block.sha1.mixer.w\[283\] net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold241 hotp.block.sha1.mixer.w\[355\] net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold252 hotp.block.sha1.mixer.w\[38\] net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold263 hotp.block.sha1.mixer.w\[316\] net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold296 hotp.block.sha1.mixer.w\[444\] net316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_68_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold274 hotp.block.sha1.mixer.w\[279\] net294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold285 hotp.block.sha1.mixer.w\[89\] net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_68_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_77_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_80_clk clknet_4_10_0_clk clknet_leaf_80_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_69_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3900_ net455 clknet_leaf_25_clk hotp.block.sha1.mixer.w\[127\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_71_clk clknet_4_11_0_clk clknet_leaf_71_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3831_ net619 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3762_ net604 clknet_leaf_79_clk hotp.block.sha1.mixer.e\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_43_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2713_ _1029_ _1041_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3693_ net98 clknet_leaf_83_clk hotp.block.sha1.mixer.c\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2644_ _0859_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2575_ _0908_ _0906_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4314_ _0215_ clknet_leaf_105_clk hotp.block.mixer.msg\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4220__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4245_ net278 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[472\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold464_I hotp.block.sha1.mixer.w\[204\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4176_ net541 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[403\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3127_ hotp.block.mixer.msg\[115\] hotp.block.mixer.msg\[116\] _1314_ _1315_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1864__A2 _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3058_ _1275_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold729_I hotp.block.sha1.mixer.w\[400\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_62_clk clknet_4_14_0_clk clknet_leaf_62_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2009_ _1621_ _0483_ _0487_ hotp.block.magic.step\[3\] _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__D net564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2549__I _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_53_clk clknet_4_13_0_clk clknet_leaf_53_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold73_I hotp.block.sha1.mixer.w\[107\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_37_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_94_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4151__D net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4243__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3990__D net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ hotp.block.sha1.mixer.h_carry _1580_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2291_ stream.digest\[2\] stream.digest\[3\] _0691_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_9_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4030_ net245 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[257\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_44_clk clknet_4_12_0_clk clknet_leaf_44_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_75_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3814_ net46 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3745_ net538 clknet_leaf_77_clk hotp.block.sha1.mixer.e\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_95_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3676_ hotp.block.debug\[0\] clknet_leaf_94_clk hotp.block.sha1.mixer.b\[31\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2627_ _0954_ _0969_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold581_I hotp.block.sha1.mixer.w\[210\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2558_ _0861_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2489_ _0846_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_11_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4228_ net57 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[455\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4159_ net735 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[386\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4236__D net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_35_clk clknet_4_7_0_clk clknet_leaf_35_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4266__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4146__D net506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_26_clk clknet_4_5_0_clk clknet_leaf_26_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3985__D net537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1860_ _1618_ _1552_ _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1791_ _1551_ _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3530_ _0107_ clknet_leaf_17_clk stream.digest\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold818 hotp.block.sha1.mixer.a\[27\] net838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold807 hotp.block.sha1.mixer.w\[477\] net827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3461_ net651 clknet_leaf_31_clk stream.key_buf\[113\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3392_ net195 clknet_leaf_51_clk stream.key_buf\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2412_ _0604_ _0745_ _0776_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_51_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2343_ _0723_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3783__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2274_ _0679_ _0680_ _0650_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4013_ net249 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[240\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_66_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4139__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold162_I hotp.block.sha1.mixer.w\[434\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_17_clk clknet_4_6_0_clk clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_hold427_I hotp.block.sha1.mixer.w\[86\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1989_ _0460_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3728_ net443 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3659_ net314 clknet_leaf_79_clk hotp.block.sha1.mixer.b\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_19_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output11_I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1994__A1 _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_hold36_I hotp.block.sha1.mixer.w\[471\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4431__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2961_ hotp.block.mixer.msg\[44\] hotp.block.mixer.msg\[45\] _1218_ _1220_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1912_ _1601_ _1476_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2892_ _1180_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1985__A1 _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1843_ _1488_ _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1774_ _1534_ _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold604 hotp.block.sha1.mixer.w\[504\] net624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold615 hotp.block.sha1.mixer.w\[76\] net635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_8_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold626 hotp.block.sha1.mixer.w\[34\] net646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3513_ _0090_ clknet_leaf_98_clk stream.digest\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold637 stream.key_buf\[62\] net657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3444_ net163 clknet_leaf_31_clk stream.key_buf\[96\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold648 hotp.block.sha1.mixer.w\[173\] net668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold659 hotp.block.sha1.mixer.b\[17\] net679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_6_clk clknet_4_1_0_clk clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3375_ net456 clknet_leaf_55_clk stream.key_buf\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2326_ stream.digest\[17\] stream.digest\[18\] _0712_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold377_I hotp.block.sha1.mixer.w\[215\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2257_ _0664_ _0666_ _0662_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_hold544_I hotp.block.sha1.mixer.w\[469\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2188_ stream.counter\[12\] _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_hold809_I hotp.block.sha1.mixer.w\[163\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold6_I hotp.block.sha1.mixer.w\[201\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4454__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3160_ _1333_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2111_ _0558_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold1 stream.key_buf\[26\] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3091_ _1294_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2042_ _0516_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_85_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3993_ net785 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[220\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold125_I hotp.block.sha1.mixer.w\[228\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2944_ _1210_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2875_ _1161_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1826_ _1586_ net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2930__I _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold401 hotp.block.sha1.mixer.w\[286\] net421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1757_ _1503_ _1518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold423 hotp.block.sha1.mixer.d\[20\] net443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold445 hotp.block.sha1.mixer.w\[216\] net465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold412 hotp.block.sha1.mixer.c\[12\] net432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold434 hotp.block.sha1.mixer.w\[484\] net454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold456 hotp.block.sha1.mixer.w\[306\] net476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1688_ _1455_ _1456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold478 hotp.block.sha1.mixer.w\[58\] net498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold467 hotp.block.sha1.mixer.c\[13\] net487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3427_ net381 clknet_leaf_36_clk stream.key_buf\[79\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold489 hotp.block.sha1.mixer.b\[12\] net509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3358_ net117 clknet_leaf_51_clk stream.key_buf\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2309_ stream.digest\[10\] stream.digest\[11\] _0701_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3289_ _0030_ clknet_leaf_37_clk stream.msg_buf\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4244__D net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3844__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_19_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4154__D net480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3993__D net785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ _0973_ _0997_ _0999_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2591_ _0914_ _0936_ _0938_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4330_ _0231_ clknet_leaf_88_clk hotp.block.mixer.msg\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4261_ net659 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[488\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_105_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3212_ hotp.block.mixer.msg\[152\] hotp.block.mixer.msg\[153\] _1361_ _1363_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input2_I in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4192_ net362 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[419\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3143_ _1323_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3074_ _1284_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2025_ _0501_ _0502_ _0503_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3022__S _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_114_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3976_ net484 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[203\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold507_I hotp.block.sha1.mixer.w\[237\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3717__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2927_ _1200_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2858_ _1160_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2789_ _1106_ _1537_ _1563_ _0378_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1809_ _1568_ _1542_ _1569_ _1570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold220 hotp.block.sha1.mixer.w\[379\] net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold231 stream.key_buf\[18\] net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold242 stream.key_buf\[19\] net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold253 hotp.block.sha1.mixer.b\[6\] net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold275 hotp.block.sha1.mixer.w\[314\] net295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4459_ _0359_ clknet_leaf_71_clk hotp.block.magic.step\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold286 hotp.block.sha1.mixer.w\[165\] net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold264 hotp.block.sha1.mixer.w\[72\] net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold297 stream.key_buf\[12\] net317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4239__D net573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3397__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4022__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__D net593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3988__D net465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3830_ net498 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3761_ net567 clknet_leaf_79_clk hotp.block.sha1.mixer.e\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_43_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2712_ _1035_ _1044_ _1045_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3692_ net431 clknet_leaf_83_clk hotp.block.sha1.mixer.c\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2643_ _0973_ _0983_ _0984_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2574_ hotp.digest\[9\] _0915_ _0921_ _0923_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4313_ _0214_ clknet_leaf_105_clk hotp.block.mixer.msg\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold192_I hotp.block.sha1.mixer.w\[432\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4244_ net155 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[471\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4175_ net315 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[402\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3126_ _1308_ _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3057_ hotp.block.mixer.msg\[85\] hotp.block.mixer.msg\[86\] _1272_ _1275_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2008_ _0484_ _0485_ _0486_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_92_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3959_ net222 clknet_leaf_1_clk hotp.block.sha1.mixer.w\[186\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4195__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2290_ _0693_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3813_ net524 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3744_ net360 clknet_leaf_77_clk hotp.block.sha1.mixer.e\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3675_ net606 clknet_leaf_94_clk hotp.block.sha1.mixer.b\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_95_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2626_ hotp.digest\[14\] _0962_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2557_ hotp.digest\[8\] _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_hold574_I hotp.block.sha1.mixer.w\[157\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2488_ _1504_ _0428_ _0827_ _0825_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3905__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4227_ net666 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[454\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4158_ net43 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[385\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4089_ net578 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[316\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3109_ _1304_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2789__A1 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4210__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4162__D net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_8_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1790_ _1550_ _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold819 stream.key_buf\[122\] net839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold808 hotp.block.sha1.mixer.w\[334\] net828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_24_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3460_ net449 clknet_leaf_31_clk stream.key_buf\[112\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3391_ net304 clknet_leaf_54_clk stream.key_buf\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2411_ _0737_ _0746_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2342_ stream.digest\[24\] stream.digest\[25\] _0722_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2273_ hotp.block.main_in _1435_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4012_ net180 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[239\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3727_ net380 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1988_ _1530_ _1548_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_hold691_I hotp.block.sha1.mixer.w\[242\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3658_ net34 clknet_leaf_76_clk hotp.block.sha1.mixer.b\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2609_ _0861_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3589_ _0162_ clknet_leaf_45_clk hotp.digest\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_3_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3004__I _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4157__D net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3996__D net307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2960_ _1219_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1911_ _0399_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2891_ hotp.block.mixer.msg\[14\] hotp.block.mixer.msg\[15\] _1176_ _1180_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1842_ _1483_ _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1773_ _1513_ _1533_ _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3512_ _0089_ clknet_leaf_98_clk stream.digest\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold616 hotp.block.sha1.mixer.d\[7\] net636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold605 hotp.block.sha1.mixer.w\[364\] net625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold627 hotp.block.sha1.mixer.b\[28\] net647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3443_ net282 clknet_leaf_30_clk stream.key_buf\[95\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold638 stream.key_buf\[56\] net658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold649 hotp.block.sha1.mixer.c\[28\] net669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3374_ stream.key_buf\[27\] clknet_leaf_56_clk stream.key_buf\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2325_ _0713_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3025__S _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2256_ _0657_ _0665_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4067__D net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2187_ _0598_ _0517_ _0601_ _0513_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_88_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_50_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_65_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4129__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2110_ stream.msg_buf\[30\] stream.msg_buf\[31\] _0556_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold2 stream.key_buf\[29\] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3090_ hotp.block.mixer.msg\[99\] hotp.block.mixer.msg\[100\] _1293_ _1294_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2041_ _0518_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3992_ net429 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[219\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_18_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2943_ hotp.block.mixer.msg\[36\] hotp.block.mixer.msg\[37\] _1208_ _1210_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_33_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2874_ _1170_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1825_ _1580_ _1584_ _1585_ _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1756_ _1501_ _1517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold402 hotp.block.sha1.mixer.w\[223\] net422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold435 hotp.block.sha1.mixer.w\[128\] net455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_64_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold413 hotp.block.sha1.mixer.w\[405\] net433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold424 hotp.block.sha1.mixer.c\[10\] net444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1687_ stream.key_state\[0\] stream.key_state\[2\] _1418_ _1401_ _1455_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
Xhold468 hotp.block.sha1.mixer.w\[32\] net488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold446 hotp.block.sha1.mixer.w\[39\] net466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold457 hotp.block.sha1.mixer.w\[496\] net477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3426_ net209 clknet_leaf_37_clk stream.key_buf\[78\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold479 hotp.block.sha1.mixer.w\[144\] net499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold487_I hotp.block.sha1.mixer.w\[138\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3357_ net232 clknet_leaf_49_clk stream.key_buf\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2308_ _0703_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3646__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3288_ _0029_ clknet_leaf_37_clk stream.msg_buf\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2239_ _0650_ _0615_ _0628_ _0408_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_95_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2590_ hotp.digest\[10\] _0937_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3669__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4260_ net291 clknet_leaf_99_clk hotp.block.sha1.mixer.w\[487\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3211_ _1362_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4191_ net534 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[418\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3142_ hotp.block.mixer.msg\[122\] hotp.block.mixer.msg\[123\] _1319_ _1323_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_87_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3073_ hotp.block.mixer.msg\[92\] hotp.block.mixer.msg\[93\] _1282_ _1284_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2024_ _0419_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold235_I hotp.block.sha1.mixer.w\[433\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3975_ net609 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[202\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2926_ hotp.block.mixer.msg\[29\] hotp.block.mixer.msg\[30\] _1197_ _1200_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold402_I hotp.block.sha1.mixer.w\[223\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2857_ _1159_ _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1808_ hotp.block.magic.step\[3\] _1535_ _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold210 stream.key_buf\[66\] net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2788_ _0365_ _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold243 hotp.block.sha1.mixer.w\[83\] net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold232 hotp.block.sha1.mixer.w\[248\] net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold221 hotp.block.sha1.mixer.w\[186\] net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1739_ hotp.block.mixer.round\[3\] _1500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4458_ _0358_ clknet_leaf_67_clk hotp.stage\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold276 hotp.block.sha1.mixer.w\[507\] net296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold287 hotp.block.sha1.mixer.w\[224\] net307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold254 hotp.block.sha1.mixer.e\[27\] net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold265 hotp.block.sha1.mixer.c\[31\] net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3409_ net657 clknet_leaf_52_clk stream.key_buf\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold298 hotp.block.sha1.mixer.w\[30\] net318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4389_ _0290_ clknet_leaf_61_clk hotp.block.mixer.msg\[101\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1867__A1 _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold11_I hotp.block.sha1.mixer.w\[84\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4165__D net727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3760_ net676 clknet_leaf_79_clk hotp.block.sha1.mixer.e\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_43_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2711_ _1029_ _1027_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3691_ net515 clknet_leaf_83_clk hotp.block.sha1.mixer.c\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2642_ _0968_ _0966_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2573_ _0851_ _0922_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _0213_ clknet_leaf_106_clk hotp.block.mixer.msg\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4243_ net56 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[470\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold185_I hotp.block.sha1.mixer.w\[390\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4174_ net154 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[401\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1849__A1 hotp.block.main_in vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3125_ _1313_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3056_ _1274_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold352_I hotp.block.sha1.mixer.w\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2007_ _1562_ _0480_ hotp.block.magic.step\[1\] _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3958_ net241 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[185\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3889_ net352 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[116\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2909_ _1190_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_4_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3999__D net520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3707__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3812_ net595 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3743_ net597 clknet_leaf_77_clk hotp.block.sha1.mixer.e\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3674_ net438 clknet_leaf_94_clk hotp.block.sha1.mixer.b\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2625_ hotp.digest\[16\] _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2556_ _0884_ _0905_ _0907_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2487_ _1497_ _1537_ _1560_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_4226_ net563 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[453\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4157_ net266 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[384\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3108_ hotp.block.mixer.msg\[107\] hotp.block.mixer.msg\[108\] _1303_ _1304_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold734_I hotp.block.sha1.mixer.w\[97\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4088_ net283 clknet_leaf_33_clk hotp.block.sha1.mixer.w\[315\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3039_ _1264_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_26_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_112_clk clknet_4_0_0_clk clknet_leaf_112_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1997__B1 _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_103_clk clknet_4_2_0_clk clknet_leaf_103_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_80_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold809 hotp.block.sha1.mixer.w\[163\] net829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2410_ _0605_ _0399_ _0765_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3390_ net146 clknet_leaf_49_clk stream.key_buf\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2341_ _0711_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_90_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2272_ stream.key_buf\[0\] _1436_ _0678_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ net768 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[238\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3029__I0 hotp.block.mixer.msg\[73\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1987_ _0454_ _0444_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2401__A1 _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3726_ net731 clknet_leaf_88_clk hotp.block.sha1.mixer.d\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4185__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3657_ net471 clknet_leaf_76_clk hotp.block.sha1.mixer.b\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2608_ _0945_ _0952_ _0953_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3588_ _0161_ clknet_leaf_65_clk hotp.digest\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2539_ _0884_ _0891_ _0892_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_3_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4209_ net479 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[436\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1994__A3 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1910_ stream.counter\[5\] _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2890_ _1179_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1841_ _1585_ _1595_ _1600_ net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1772_ _1498_ _1500_ _1502_ _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_13_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold617 hotp.block.sha1.mixer.w\[301\] net637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3511_ _0088_ clknet_leaf_97_clk stream.digest\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold606 hotp.block.sha1.mixer.w\[174\] net626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3442_ net139 clknet_leaf_31_clk stream.key_buf\[94\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold628 stream.key_buf\[24\] net648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold639 hotp.block.sha1.mixer.w\[489\] net659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3373_ net21 clknet_leaf_55_clk stream.key_buf\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2324_ stream.digest\[16\] stream.digest\[17\] _0712_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2255_ stream.digest\[1\] stream.digest\[5\] stream.digest\[9\] stream.digest\[13\]
+ _0658_ _0659_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2186_ stream.msg_buf\[0\] _0408_ _0600_ net1 _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold432_I hotp.block.sha1.mixer.w\[448\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3709_ net404 clknet_leaf_85_clk hotp.block.sha1.mixer.d\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_4_12_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4200__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold3 hotp.block.sha1.mixer.w\[253\] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4168__D net327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2040_ stream.msg_buf\[0\] stream.msg_buf\[1\] _0517_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ net374 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[218\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2942_ _1209_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_33_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1958__A3 hotp.block.sha1.mixer.c\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2873_ hotp.block.mixer.msg\[6\] hotp.block.mixer.msg\[7\] _1166_ _1170_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1824_ _1488_ _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_26_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1755_ _1506_ _1515_ _1516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold436 stream.key_buf\[28\] net456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_52_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold414 hotp.block.sha1.mixer.w\[426\] net434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_13_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold403 hotp.block.sha1.mixer.w\[153\] net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold425 hotp.block.sha1.mixer.w\[51\] net445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_20_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold458 hotp.block.sha1.mixer.w\[105\] net478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1686_ _1450_ _1454_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold469 hotp.block.sha1.mixer.a\[30\] net489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold447 hotp.block.sha1.mixer.a\[21\] net467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3425_ net473 clknet_leaf_37_clk stream.key_buf\[77\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3356_ net329 clknet_leaf_49_clk stream.key_buf\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold382_I hotp.block.sha1.mixer.w\[85\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3287_ _0028_ clknet_leaf_38_clk stream.msg_buf\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2307_ stream.digest\[9\] stream.digest\[10\] _0701_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2238_ _0510_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2169_ stream.msg_buf\[56\] stream.msg_buf\[57\] _0587_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_92_clk clknet_4_8_0_clk clknet_leaf_92_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_hold814_I hotp.block.sha1.mixer.w\[256\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_83_clk clknet_4_10_0_clk clknet_leaf_83_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2533__B _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4246__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3210_ hotp.block.mixer.msg\[151\] hotp.block.mixer.msg\[152\] _1361_ _1362_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4190_ net213 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[417\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3141_ _1322_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3072_ _1283_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_19_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2023_ hotp.block.debug\[1\] _0500_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_74_clk clknet_4_11_0_clk clknet_leaf_74_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ net746 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[201\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2925_ _1199_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2856_ _1611_ _0418_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_26_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1807_ hotp.block.magic.step\[3\] _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2787_ _1100_ _1105_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold211 hotp.block.sha1.mixer.a\[12\] net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold200 hotp.block.sha1.mixer.w\[218\] net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold233 stream.key_buf\[42\] net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold244 hotp.block.sha1.mixer.w\[158\] net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1738_ _1498_ _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold222 hotp.block.sha1.mixer.w\[192\] net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1669_ _1438_ _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4457_ _0357_ clknet_leaf_67_clk hotp.block.mixer.stage\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold255 hotp.block.sha1.mixer.w\[383\] net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold266 hotp.block.sha1.mixer.e\[24\] net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold277 hotp.block.sha1.mixer.w\[13\] net297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3408_ net801 clknet_leaf_53_clk stream.key_buf\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold764_I hotp.block.sha1.mixer.w\[159\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold288 hotp.block.sha1.mixer.w\[276\] net308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold299 hotp.block.sha1.mixer.b\[10\] net319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4388_ _0289_ clknet_leaf_60_clk hotp.block.mixer.msg\[100\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3339_ _0002_ clknet_leaf_43_clk stream.msg_state\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_37_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_64_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_65_clk clknet_4_14_0_clk clknet_leaf_65_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_79_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4269__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__D net575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_17_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_56_clk clknet_4_15_0_clk clknet_leaf_56_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3232__A1 _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2710_ hotp.digest\[25\] _0862_ _1041_ _1043_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3636__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_0_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4181__D net574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3690_ net464 clknet_leaf_83_clk hotp.block.sha1.mixer.c\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2641_ hotp.digest\[17\] _0915_ _0979_ _0982_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_23_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2572_ _0897_ _0920_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2489__I _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4311_ _0212_ clknet_leaf_106_clk hotp.block.mixer.msg\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_73_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4242_ net808 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[469\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4173_ net256 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[400\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3124_ hotp.block.mixer.msg\[114\] hotp.block.mixer.msg\[115\] _1309_ _1313_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold178_I hotp.block.sha1.mixer.w\[175\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3055_ hotp.block.mixer.msg\[84\] hotp.block.mixer.msg\[85\] _1272_ _1274_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_47_clk clknet_4_12_0_clk clknet_leaf_47_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2006_ _0453_ _0455_ _1551_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3957_ net549 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[184\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2908_ hotp.block.mixer.msg\[21\] hotp.block.mixer.msg\[22\] _1187_ _1190_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3888_ net587 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[115\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2839_ _0436_ _0499_ _1144_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_38_clk clknet_4_7_0_clk clknet_leaf_38_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_68_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4091__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_29_clk clknet_4_5_0_clk clknet_leaf_29_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_48_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3811_ net466 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_99_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3742_ net396 clknet_leaf_77_clk hotp.block.sha1.mixer.e\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3673_ net755 clknet_leaf_94_clk hotp.block.sha1.mixer.b\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_81_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2624_ _0945_ _0965_ _0967_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2555_ hotp.digest\[6\] _0906_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2486_ hotp.digest\[1\] _0843_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4225_ net79 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[452\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4156_ net144 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[383\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3107_ _1287_ _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4087_ net129 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[314\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold727_I hotp.block.sha1.mixer.w\[143\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3038_ hotp.block.mixer.msg\[77\] hotp.block.mixer.msg\[78\] _1261_ _1264_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2857__I _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1997__A1 _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold71_I hotp.block.sha1.mixer.w\[255\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2340_ _0721_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1671__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2271_ _0604_ _0676_ _0677_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4010_ net788 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[237\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1988__A1 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3029__I1 hotp.block.mixer.msg\[74\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1986_ _0382_ _0459_ _0462_ _0464_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_71_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3725_ net326 clknet_leaf_87_clk hotp.block.sha1.mixer.d\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_9_clk clknet_4_1_0_clk clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3656_ net509 clknet_leaf_76_clk hotp.block.sha1.mixer.b\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2607_ _0939_ _0937_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3587_ _0160_ clknet_leaf_65_clk hotp.digest\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold677_I hotp.block.sha1.mixer.w\[127\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2538_ _0878_ _0876_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2469_ _0819_ _0826_ _0468_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_4208_ net435 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[435\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_3_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ net100 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[366\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1957__S _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_76_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3847__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1840_ _1585_ _1599_ _1600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1771_ hotp.block.mixer.msg\[0\] _1516_ _1527_ _1531_ _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_3510_ _0087_ clknet_leaf_98_clk stream.digest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold618 stream.key_buf\[77\] net638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold607 hotp.block.sha1.mixer.w\[43\] net627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3441_ net301 clknet_leaf_30_clk stream.key_buf\[93\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold629 hotp.block.sha1.mixer.w\[371\] net649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3372_ net712 clknet_leaf_55_clk stream.key_buf\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2323_ _0711_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2254_ _0652_ _0663_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2185_ _1463_ _1464_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold160_I hotp.block.sha1.mixer.w\[240\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold258_I hotp.block.sha1.mixer.w\[473\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ _0442_ _0446_ _0447_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3708_ _0010_ clknet_leaf_93_clk hotp.block.sha1.mixer.c\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3639_ net838 clknet_leaf_93_clk hotp.block.sha1.mixer.a\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4274__D net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4025__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold4 hotp.block.sha1.mixer.w\[243\] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_89_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4184__D net526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3990_ net220 clknet_leaf_114_clk hotp.block.sha1.mixer.w\[217\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2941_ hotp.block.mixer.msg\[35\] hotp.block.mixer.msg\[36\] _1208_ _1209_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_33_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2872_ _1169_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1823_ _1581_ _1582_ _1478_ _1583_ _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_44_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1754_ _1503_ _1509_ _1514_ _1501_ _1515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xhold426 hotp.block.sha1.mixer.w\[171\] net446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold404 hotp.block.sha1.mixer.w\[194\] net424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold415 hotp.block.sha1.mixer.w\[436\] net435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_110_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3424_ net638 clknet_leaf_37_clk stream.key_buf\[76\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1685_ stream.msg_state\[3\] _1453_ _1428_ _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold448 hotp.block.sha1.mixer.d\[2\] net468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold459 hotp.block.sha1.mixer.w\[437\] net479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold437 hotp.block.sha1.mixer.a\[24\] net457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3355_ net320 clknet_leaf_50_clk stream.key_buf\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3286_ _0027_ clknet_leaf_38_clk stream.msg_buf\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2306_ _0702_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2237_ _0624_ _0630_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2168_ _0590_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2099_ stream.msg_buf\[25\] stream.msg_buf\[26\] _0551_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold4_I hotp.block.sha1.mixer.w\[243\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4198__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3026__I _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3901__D net763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2834__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4179__D net394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3140_ hotp.block.mixer.msg\[121\] hotp.block.mixer.msg\[122\] _1319_ _1322_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3071_ hotp.block.mixer.msg\[91\] hotp.block.mixer.msg\[92\] _1282_ _1283_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3811__D net466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2022_ hotp.block.debug\[1\] _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_18_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3973_ net26 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[200\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2924_ hotp.block.mixer.msg\[28\] hotp.block.mixer.msg\[29\] _1197_ _1199_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold123_I hotp.block.sha1.mixer.w\[381\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2855_ hotp.block.mixer.msg\[0\] _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_115_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1806_ _1549_ _1565_ _1566_ hotp.block.magic.step\[4\] _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold201 stream.key_buf\[150\] net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2786_ stream.key_counter\[7\] _1103_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold212 stream.key_buf\[10\] net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold223 hotp.block.sha1.mixer.w\[3\] net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold234 hotp.block.sha1.mixer.w\[511\] net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1737_ hotp.block.mixer.round\[1\] _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold267 stream.key_buf\[134\] net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1668_ _1436_ _1437_ _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4456_ _0356_ clknet_leaf_67_clk hotp.block.mixer.stage\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold256 hotp.block.sha1.mixer.w\[44\] net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold245 hotp.block.sha1.mixer.w\[183\] net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold278 hotp.block.sha1.mixer.c\[7\] net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3407_ net126 clknet_leaf_52_clk stream.key_buf\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold289 hotp.block.sha1.mixer.w\[132\] net309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3908__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4387_ _0288_ clknet_leaf_60_clk hotp.block.mixer.msg\[99\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3338_ _0001_ clknet_leaf_43_clk stream.msg_state\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3269_ _0367_ _0368_ _0916_ _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_101_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold790 hotp.block.sha1.mixer.c\[9\] net810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_86_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4213__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2640_ _0980_ _0981_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2571_ hotp.digest\[7\] _0920_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3806__D net646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4310_ _0211_ clknet_leaf_105_clk hotp.block.mixer.msg\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4241_ net564 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[468\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4172_ net749 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[399\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3123_ _1312_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3054_ _1273_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2005_ _0480_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_hold240_I hotp.block.sha1.mixer.w\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold338_I hotp.block.sha1.mixer.w\[66\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3956_ net492 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[183\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2907_ _1189_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold505_I hotp.block.sha1.mixer.w\[423\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3887_ net399 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[114\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2838_ _0457_ _0498_ _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2769_ stream.key_counter\[0\] _1456_ _0735_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3730__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4439_ _0340_ clknet_leaf_91_clk hotp.block.mixer.msg\[151\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3880__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3810_ net272 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4192__D net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3741_ net342 clknet_leaf_74_clk hotp.block.sha1.mixer.e\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3672_ net647 clknet_leaf_94_clk hotp.block.sha1.mixer.b\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2623_ hotp.digest\[14\] _0966_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2554_ _0875_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_63_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2485_ hotp.digest\[0\] hotp.digest\[39\] _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_10_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4224_ net239 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[451\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_78_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4155_ net275 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[382\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3106_ _1302_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold455_I hotp.block.sha1.mixer.w\[155\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4086_ net295 clknet_leaf_33_clk hotp.block.sha1.mixer.w\[313\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3037_ _1263_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_16_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3939_ net535 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[166\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1758__A2 _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1930__A2 _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2270_ stream.counter\[7\] _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1988__A2 _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1985_ _1574_ _0448_ _0463_ _1620_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_55_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3724_ net349 clknet_leaf_87_clk hotp.block.sha1.mixer.d\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3655_ net389 clknet_leaf_76_clk hotp.block.sha1.mixer.b\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2606_ hotp.digest\[13\] _0915_ _0949_ _0951_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_101_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3586_ _0159_ clknet_leaf_65_clk hotp.digest\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2537_ hotp.digest\[5\] _0842_ _0888_ _0890_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2468_ _1528_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_3_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ net244 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[434\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2399_ _0607_ _0765_ _0747_ _0751_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4138_ net733 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[365\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4069_ net35 clknet_leaf_20_clk hotp.block.sha1.mixer.w\[296\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_50_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1770_ _1530_ _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold608 hotp.block.sha1.mixer.w\[398\] net628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold619 stream.key_buf\[100\] net639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3440_ net138 clknet_leaf_31_clk stream.key_buf\[92\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3371_ net648 clknet_leaf_55_clk stream.key_buf\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3814__D net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2322_ _0689_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3941__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2253_ stream.digest\[17\] stream.digest\[21\] stream.digest\[25\] stream.digest\[29\]
+ _0653_ _0654_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2184_ _0598_ _0517_ _0599_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1968_ _1500_ hotp.block.mixer.round\[2\] _1511_ _1510_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_114_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1899_ _1582_ _1601_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3707_ net285 clknet_leaf_94_clk hotp.block.sha1.mixer.c\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3638_ net376 clknet_leaf_93_clk hotp.block.sha1.mixer.a\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3569_ _0142_ clknet_leaf_48_clk hotp.digest\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1888__A1 _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold5 hotp.block.sha1.mixer.w\[410\] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_89_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2940_ _1202_ _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2871_ hotp.block.mixer.msg\[5\] hotp.block.mixer.msg\[6\] _1166_ _1169_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3494__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1822_ _1479_ _1483_ _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_13_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1753_ _1513_ _1514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold405 hotp.block.sha1.mixer.w\[323\] net425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1684_ _1452_ _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold427 hotp.block.sha1.mixer.w\[86\] net447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold416 hotp.block.sha1.mixer.c\[23\] net436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3423_ net630 clknet_leaf_37_clk stream.key_buf\[75\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold438 hotp.block.sha1.mixer.d\[24\] net458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold449 hotp.block.sha1.mixer.w\[21\] net469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3354_ net118 clknet_leaf_49_clk stream.key_buf\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3285_ _0026_ clknet_leaf_38_clk stream.msg_buf\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2305_ stream.digest\[8\] stream.digest\[9\] _0701_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2236_ _0631_ _0630_ _0648_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_hold270_I hotp.block.sha1.mixer.w\[464\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2167_ stream.msg_buf\[55\] stream.msg_buf\[56\] _0587_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2098_ _0550_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold535_I hotp.block.sha1.mixer.w\[229\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3837__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4142__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3070_ _1266_ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_38_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4195__D net525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2021_ _0436_ _0499_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ net775 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[199\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2923_ _1198_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2854_ _1152_ _0434_ _1157_ _1155_ _0431_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_45_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2785_ _1102_ _1104_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1805_ _1555_ _1557_ _1534_ _1566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_5_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold116_I hotp.block.sha1.mixer.w\[425\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1736_ _1496_ _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold202 hotp.block.sha1.mixer.w\[187\] net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold213 hotp.block.sha1.mixer.w\[349\] net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold235 hotp.block.sha1.mixer.w\[433\] net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold224 hotp.block.sha1.mixer.w\[435\] net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold257 hotp.block.sha1.mixer.w\[338\] net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1667_ stream.counter\[7\] stream.counter\[6\] _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold268 hotp.block.sha1.mixer.w\[50\] net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold246 hotp.block.sha1.mixer.w\[385\] net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4455_ _0355_ clknet_leaf_68_clk hotp.block.mixer.round\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3406_ net190 clknet_leaf_51_clk stream.key_buf\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4386_ _0287_ clknet_leaf_62_clk hotp.block.mixer.msg\[98\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold279 hotp.block.sha1.mixer.w\[78\] net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3337_ _0000_ clknet_leaf_46_clk stream.msg_state\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3268_ _1395_ _0428_ _1398_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2219_ _1415_ _0632_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3199_ _1355_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3449__D net324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2142__S _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold780 hotp.block.sha1.mixer.w\[342\] net800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold791 hotp.block.sha1.mixer.w\[480\] net811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3912__D net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold94_I hotp.block.sha1.mixer.w\[359\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_97_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2570_ _0916_ _0917_ _0919_ hotp.digest\[10\] _0847_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_77_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2987__S _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4240_ net529 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[467\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4171_ net592 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[398\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3122_ hotp.block.mixer.msg\[113\] hotp.block.mixer.msg\[114\] _1309_ _1312_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3053_ hotp.block.mixer.msg\[83\] hotp.block.mixer.msg\[84\] _1272_ _1273_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ _1543_ _0481_ _0482_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_106_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3955_ net265 clknet_leaf_1_clk hotp.block.sha1.mixer.w\[182\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2906_ hotp.block.mixer.msg\[20\] hotp.block.mixer.msg\[21\] _1187_ _1189_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4188__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3886_ net812 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[113\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2837_ hotp.block.sha1.mixer.a_carry\[1\] _1142_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2768_ _1065_ _1093_ _1094_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2699_ _1019_ _1027_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1719_ _1481_ _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2897__S _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4438_ _0339_ clknet_leaf_91_clk hotp.block.mixer.msg\[150\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4369_ _0270_ clknet_leaf_72_clk hotp.block.mixer.msg\[81\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3405__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3907__D net719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1775__I hotp.block.magic.step\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4330__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_106_clk clknet_4_2_0_clk clknet_leaf_106_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3740_ hotp.block.sha1.mixer.c\[0\] clknet_leaf_86_clk hotp.block.sha1.mixer.d\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ net725 clknet_leaf_93_clk hotp.block.sha1.mixer.b\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2622_ _0875_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2553_ _0897_ _0898_ _0904_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2484_ _0841_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4223_ net130 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[450\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_52_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold183_I hotp.block.sha1.mixer.w\[208\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4154_ net480 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[381\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4085_ net502 clknet_leaf_33_clk hotp.block.sha1.mixer.w\[312\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3105_ hotp.block.mixer.msg\[106\] hotp.block.mixer.msg\[107\] _1298_ _1302_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3036_ hotp.block.mixer.msg\[76\] hotp.block.mixer.msg\[77\] _1261_ _1263_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold350_I hotp.block.sha1.mixer.w\[169\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold615_I hotp.block.sha1.mixer.w\[76\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3938_ net185 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[165\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3869_ net754 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[96\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_14_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4203__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1930__A3 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_94_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold57_I hotp.block.sha1.mixer.w\[414\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1984_ _0460_ _0441_ _0447_ _1550_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3870__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3723_ net702 clknet_leaf_87_clk hotp.block.sha1.mixer.d\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3654_ net319 clknet_leaf_80_clk hotp.block.sha1.mixer.b\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2605_ _0851_ _0950_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3585_ _0158_ clknet_leaf_65_clk hotp.digest\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2536_ _0851_ _0889_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2467_ _1521_ _1508_ _1625_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4206_ net182 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[433\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2398_ stream.counter\[4\] _0607_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4137_ net622 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[364\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4068_ net313 clknet_leaf_41_clk hotp.block.sha1.mixer.w\[295\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_65_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3019_ _1253_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3045__I _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3920__D net481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_62_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold609 hotp.block.sha1.mixer.w\[440\] net629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_69_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3370_ net782 clknet_leaf_55_clk stream.key_buf\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2321_ _0710_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4198__D net434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2252_ _0656_ _0661_ _0662_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_15_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2183_ stream.msg_buf\[62\] _0517_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3706_ _0009_ clknet_leaf_93_clk hotp.block.sha1.mixer.c\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1967_ hotp.block.mixer.round\[5\] _1511_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1898_ _1609_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3637_ net566 clknet_leaf_93_clk hotp.block.sha1.mixer.a\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3568_ _0141_ clknet_leaf_48_clk hotp.digest\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2519_ _0855_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3499_ net333 clknet_leaf_20_clk stream.key_buf\[151\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_71_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3740__D hotp.block.sha1.mixer.c\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_95_clk clknet_4_9_0_clk clknet_leaf_95_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3915__D net747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold6 hotp.block.sha1.mixer.w\[201\] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_86_clk clknet_4_8_0_clk clknet_leaf_86_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_89_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3639__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2870_ _1168_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1821_ _1481_ _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_10_clk clknet_4_1_0_clk clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1752_ _1510_ _1511_ _1512_ _1513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_111_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1683_ _1420_ _1451_ _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold417 hotp.block.sha1.mixer.w\[281\] net437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_52_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold406 hotp.block.sha1.mixer.e\[23\] net426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3422_ net690 clknet_leaf_37_clk stream.key_buf\[74\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold439 hotp.block.sha1.mixer.d\[13\] net459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold428 hotp.block.sha1.mixer.w\[234\] net448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3353_ net822 clknet_leaf_47_clk stream.key_buf\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3284_ _0025_ clknet_leaf_38_clk stream.msg_buf\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2304_ _0690_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2235_ _0630_ _0647_ _0413_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_77_clk clknet_4_11_0_clk clknet_leaf_77_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2166_ _0589_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2097_ _0515_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold528_I hotp.block.sha1.mixer.w\[79\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3253__A1 _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2999_ _1241_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_73_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_68_clk clknet_4_9_0_clk clknet_leaf_68_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4094__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3931__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_59_clk clknet_4_14_0_clk clknet_leaf_59_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_38_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2020_ _0457_ _0498_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3971_ net680 clknet_leaf_108_clk hotp.block.sha1.mixer.w\[198\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3235__A1 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2922_ hotp.block.mixer.msg\[27\] hotp.block.mixer.msg\[28\] _1197_ _1198_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2853_ hotp.block.sha1.mixer.a_carry\[2\] hotp.block.sha1.mixer.a_carry\[1\] _1142_
+ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2784_ _0413_ _1456_ _1103_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1804_ _1563_ _1564_ _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1735_ hotp.block.mixer.round\[0\] _1496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_113_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold203 stream.key_buf\[46\] net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold225 hotp.block.sha1.mixer.w\[258\] net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold214 hotp.block.sha1.mixer.w\[226\] net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1666_ stream.counter\[8\] _1435_ _1436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold247 hotp.block.sha1.mixer.w\[424\] net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold236 hotp.block.sha1.mixer.w\[401\] net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold269 hotp.block.sha1.mixer.w\[146\] net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold258 hotp.block.sha1.mixer.w\[473\] net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _0354_ clknet_leaf_94_clk hotp.block.mixer.round\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3405_ net616 clknet_leaf_51_clk stream.key_buf\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4385_ _0286_ clknet_leaf_71_clk hotp.block.mixer.msg\[97\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3336_ _0077_ clknet_leaf_43_clk stream.msg_buf\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3267_ _0367_ _0368_ _0372_ _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2218_ stream.state\[2\] _0631_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3198_ hotp.block.mixer.msg\[146\] hotp.block.mixer.msg\[147\] _1351_ _1355_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2149_ stream.msg_buf\[47\] stream.msg_buf\[48\] _0577_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold781 stream.key_buf\[61\] net801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold770 stream.key_buf\[16\] net790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold792 hotp.block.sha1.mixer.w\[114\] net812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_86_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_24_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2333__S _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4170_ net628 clknet_leaf_109_clk hotp.block.sha1.mixer.w\[397\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3827__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3121_ _1311_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_42_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3052_ _1266_ _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2003_ _1551_ _0455_ _0449_ _0461_ hotp.block.magic.step\[2\] _0482_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_TAPCELL_ROW_106_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3954_ net302 clknet_leaf_0_clk hotp.block.sha1.mixer.w\[181\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3885_ net730 clknet_leaf_23_clk hotp.block.sha1.mixer.w\[112\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_51_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2905_ _1188_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2836_ _1139_ _1140_ _1141_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2767_ _1082_ _0838_ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2698_ _1029_ _1020_ _1032_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1718_ seg.digit\[1\] _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1649_ _1418_ _1419_ _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2977__I _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4437_ _0338_ clknet_leaf_91_clk hotp.block.mixer.msg\[149\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4368_ _0269_ clknet_leaf_73_clk hotp.block.mixer.msg\[80\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3319_ _0060_ clknet_leaf_41_clk stream.msg_buf\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4299_ _0200_ clknet_leaf_104_clk hotp.block.mixer.msg\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2186__B2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1791__I _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3923__D net798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3670_ net379 clknet_leaf_93_clk hotp.block.sha1.mixer.b\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2621_ _0959_ _0940_ _0964_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2552_ _0868_ _0903_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2483_ _0840_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4222_ net111 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[449\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3833__D net321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4153_ net143 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[380\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4084_ net580 clknet_leaf_33_clk hotp.block.sha1.mixer.w\[311\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3104_ _1301_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3035_ _1262_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold608_I hotp.block.sha1.mixer.w\[398\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold510_I hotp.block.sha1.mixer.w\[235\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3937_ net306 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[164\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3868_ net105 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[95\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2819_ hotp.digest\[34\] _0838_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3799_ net742 clknet_leaf_107_clk hotp.block.sha1.mixer.w\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_6_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_45_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3918__D net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3672__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4178__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1983_ _0461_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3722_ net490 clknet_leaf_87_clk hotp.block.sha1.mixer.d\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3653_ net821 clknet_leaf_80_clk hotp.block.sha1.mixer.b\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2604_ _0930_ _0948_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3584_ _0157_ clknet_leaf_65_clk hotp.digest\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2535_ _0867_ _0887_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2466_ _0418_ _0823_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4205_ net255 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[432\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2397_ _0748_ _0763_ stream.counter\[4\] _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4136_ net625 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[363\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold460_I hotp.block.sha1.mixer.w\[382\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4067_ net50 clknet_leaf_20_clk hotp.block.sha1.mixer.w\[294\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_65_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3018_ hotp.block.mixer.msg\[68\] hotp.block.mixer.msg\[69\] _1251_ _1253_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2320_ stream.digest\[15\] stream.digest\[16\] _0706_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2251_ _1442_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2182_ stream.msg_buf\[63\] _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_34_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1966_ _0416_ _0444_ hotp.block.sha1.mixer.d\[0\] _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3705_ net63 clknet_leaf_92_clk hotp.block.sha1.mixer.c\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1897_ _1601_ _1602_ _1603_ _0389_ net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_31_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3636_ net457 clknet_leaf_93_clk hotp.block.sha1.mixer.a\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3567_ _0140_ clknet_leaf_48_clk hotp.digest\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2518_ _0867_ _0860_ _0873_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_hold675_I hotp.block.sha1.mixer.w\[411\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3498_ net709 clknet_leaf_19_clk stream.key_buf\[150\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2449_ hotp.index\[3\] _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_71_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4119_ net682 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[346\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3860__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3931__D net784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold7 hotp.block.sha1.mixer.b\[24\] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_89_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ _1479_ _1581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_13_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1751_ hotp.block.mixer.round\[6\] _1512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1682_ _1428_ stream.msg_state\[0\] _1417_ net3 _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xhold407 hotp.block.sha1.mixer.w\[265\] net427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_52_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold418 hotp.block.sha1.mixer.b\[30\] net438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold429 stream.key_buf\[113\] net449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3421_ net55 clknet_leaf_52_clk stream.key_buf\[73\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3352_ net49 clknet_leaf_48_clk stream.key_buf\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4002__D net501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2303_ _0700_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_111_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3283_ _0024_ clknet_leaf_38_clk stream.msg_buf\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3841__D net547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2234_ _1401_ _1434_ _0633_ _0643_ _1429_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2165_ stream.msg_buf\[54\] stream.msg_buf\[55\] _0587_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2096_ _0549_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2998_ hotp.block.mixer.msg\[60\] hotp.block.mixer.msg\[61\] _1239_ _1241_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1949_ _1537_ _1560_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_17_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3733__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3619_ net741 clknet_leaf_75_clk hotp.block.sha1.mixer.a\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_61_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3883__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4239__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_76_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_88_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_14_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3926__D net663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_97_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_29_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3970_ net38 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[197\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2921_ _1181_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2852_ _1149_ _1156_ _0734_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2783_ stream.key_counter\[5\] stream.key_counter\[6\] _1098_ _1103_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_72_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1803_ _1554_ _1557_ _1564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3836__D net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1734_ hotp.block.mixer.stage\[0\] _1495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold204 stream.key_buf\[36\] net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold226 hotp.block.sha1.mixer.w\[346\] net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold215 hotp.block.sha1.mixer.b\[4\] net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4453_ _0353_ clknet_leaf_94_clk hotp.block.mixer.round\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_113_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3404_ net662 clknet_leaf_51_clk stream.key_buf\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold248 hotp.block.sha1.mixer.w\[344\] net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1665_ stream.counter\[12\] stream.counter\[11\] stream.counter\[10\] stream.counter\[9\]
+ _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
Xhold237 hotp.block.sha1.mixer.w\[74\] net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold259 hotp.block.sha1.mixer.d\[27\] net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4384_ _0285_ clknet_leaf_71_clk hotp.block.mixer.msg\[96\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3335_ _0076_ clknet_leaf_43_clk stream.msg_buf\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3266_ _1397_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2217_ _0508_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_hold540_I hotp.block.sha1.mixer.w\[395\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3197_ _1354_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2148_ _0579_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2079_ _0529_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3746__D net837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold782 hotp.block.sha1.mixer.w\[109\] net802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold771 hotp.block.sha1.mixer.e\[14\] net791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold760 hotp.block.sha1.mixer.a\[11\] net780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold793 hotp.block.sha1.mixer.b\[8\] net813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_93_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1779__A2 _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3120_ hotp.block.mixer.msg\[112\] hotp.block.mixer.msg\[113\] _1309_ _1311_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3051_ _1271_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2002_ _0452_ _0480_ _1547_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3953_ net200 clknet_leaf_1_clk hotp.block.sha1.mixer.w\[180\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3884_ net181 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[111\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2904_ hotp.block.mixer.msg\[19\] hotp.block.mixer.msg\[20\] _1187_ _1188_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold121_I hotp.block.sha1.mixer.w\[225\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2835_ _1590_ _0497_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_60_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2766_ _0403_ _1091_ _1092_ _0862_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2697_ _1030_ _1031_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1717_ seg.digit\[1\] seg.digit\[0\] _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1648_ net2 net3 _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_hold490_I hotp.block.sha1.mixer.w\[189\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4436_ _0337_ clknet_leaf_92_clk hotp.block.mixer.msg\[148\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3154__I _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4367_ _0268_ clknet_leaf_73_clk hotp.block.mixer.msg\[79\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3318_ _0059_ clknet_leaf_41_clk stream.msg_buf\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold755_I hotp.block.sha1.mixer.w\[200\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4298_ _0199_ clknet_leaf_91_clk hotp.block.mixer.msg\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3921__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3249_ _1380_ _1387_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold590 stream.key_buf\[105\] net610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2852__B _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2344__S _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2620_ _0954_ _0963_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2551_ hotp.digest\[5\] _0900_ _0902_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2482_ _0829_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4221_ net583 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[448\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_52_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4010__D net788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4152_ net694 clknet_leaf_110_clk hotp.block.sha1.mixer.w\[379\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4083_ net531 clknet_leaf_33_clk hotp.block.sha1.mixer.w\[310\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3103_ hotp.block.mixer.msg\[105\] hotp.block.mixer.msg\[106\] _1298_ _1301_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_108_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3034_ hotp.block.mixer.msg\[75\] hotp.block.mixer.msg\[76\] _1261_ _1262_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold169_I hotp.block.sha1.mixer.w\[236\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3936_ net805 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[163\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_63_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3867_ net258 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[94\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2818_ hotp.digest\[33\] _1128_ _1129_ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3798_ net214 clknet_leaf_106_clk hotp.block.sha1.mixer.w\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2749_ _1050_ _1071_ _1060_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4419_ _0320_ clknet_leaf_72_clk hotp.block.mixer.msg\[131\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3934__D net824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2339__S _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _0460_ _1547_ _1529_ _0441_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_71_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3721_ net459 clknet_leaf_87_clk hotp.block.sha1.mixer.d\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4005__D net417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3652_ net813 clknet_leaf_80_clk hotp.block.sha1.mixer.b\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2603_ hotp.digest\[11\] _0948_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3583_ _0156_ clknet_leaf_65_clk hotp.digest\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_2_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3844__D net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2534_ hotp.digest\[3\] _0887_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2465_ _0822_ hotp.block.mixer.stage\[1\] hotp.block.mixer.stage\[0\] _0823_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_54_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2396_ _1426_ _0746_ _0608_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_hold286_I hotp.block.sha1.mixer.w\[165\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4204_ net212 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[431\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4135_ net197 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[362\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_3_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4066_ net121 clknet_leaf_28_clk hotp.block.sha1.mixer.w\[293\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4272__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3017_ _1252_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold718_I hotp.block.sha1.mixer.w\[100\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3919_ net787 clknet_leaf_7_clk hotp.block.sha1.mixer.w\[146\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2010__A1 _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3929__D net594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2250_ _0657_ _0660_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_108_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2181_ _0597_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3839__D net559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_117_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_60_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1965_ _0443_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3704_ net669 clknet_leaf_92_clk hotp.block.sha1.mixer.c\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1896_ _1602_ _0388_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3635_ net39 clknet_leaf_85_clk hotp.block.sha1.mixer.a\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3566_ _0139_ clknet_leaf_48_clk hotp.digest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2517_ _0868_ _0872_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3497_ net221 clknet_leaf_42_clk stream.key_buf\[149\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2448_ _0804_ _0806_ _0759_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_hold668_I hotp.block.sha1.mixer.w\[212\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2379_ _1453_ _0643_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_71_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4118_ net246 clknet_leaf_18_clk hotp.block.sha1.mixer.w\[345\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4049_ net806 clknet_leaf_18_clk hotp.block.sha1.mixer.w\[276\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2241__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3031__I0 hotp.block.mixer.msg\[74\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold8 hotp.block.sha1.mixer.w\[73\] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_89_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1750_ hotp.block.mixer.round\[4\] _1511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold408 stream.key_buf\[107\] net428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1681_ _1445_ _1447_ _1449_ _1428_ _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3420_ net664 clknet_leaf_52_clk stream.key_buf\[72\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold419 stream.key_buf\[99\] net439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3351_ net124 clknet_leaf_49_clk stream.key_buf\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2302_ stream.digest\[7\] stream.digest\[8\] _0696_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_111_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3282_ _0023_ clknet_leaf_39_clk stream.msg_buf\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2233_ _1415_ _0630_ _0645_ _0646_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2164_ _0588_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2095_ stream.msg_buf\[24\] stream.msg_buf\[25\] _0545_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2997_ _1240_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1948_ _0427_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1879_ _0371_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold785_I hotp.block.sha1.mixer.w\[164\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3618_ net783 clknet_leaf_75_clk hotp.block.sha1.mixer.a\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3549_ _0126_ clknet_leaf_19_clk stream.counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3942__D net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2920_ _1196_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2851_ _1151_ _1154_ _1155_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2782_ stream.key_counter\[5\] _1098_ stream.key_counter\[6\] _1102_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1802_ _1562_ _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1733_ _1490_ _1491_ _1489_ _1494_ net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_25_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4013__D net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold216 hotp.block.sha1.mixer.w\[431\] net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4452_ _0352_ clknet_leaf_94_clk hotp.block.mixer.round\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold205 hotp.block.sha1.mixer.a\[15\] net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold227 stream.key_buf\[81\] net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold249 stream.key_buf\[130\] net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3403_ net658 clknet_leaf_51_clk stream.key_buf\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1664_ _1427_ _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold238 hotp.block.sha1.mixer.w\[95\] net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_111_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4383_ _0284_ clknet_leaf_71_clk hotp.block.mixer.msg\[95\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3852__D net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3334_ _0075_ clknet_leaf_43_clk stream.msg_buf\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3265_ _0685_ _1548_ _1575_ _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2216_ _0629_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3196_ hotp.block.mixer.msg\[145\] hotp.block.mixer.msg\[146\] _1351_ _1354_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_37_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2147_ stream.msg_buf\[46\] stream.msg_buf\[47\] _0577_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2078_ _0539_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold533_I hotp.block.sha1.mixer.w\[104\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold700_I hotp.block.sha1.mixer.w\[247\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4206__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold761 hotp.block.sha1.mixer.w\[45\] net781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold750 hotp.block.sha1.mixer.w\[378\] net770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold772 hotp.block.sha1.mixer.w\[16\] net792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold794 stream.key_buf\[22\] net814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold783 hotp.block.sha1.mixer.w\[466\] net803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_86_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3937__D net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3050_ hotp.block.mixer.msg\[82\] hotp.block.mixer.msg\[83\] _1267_ _1271_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2001_ _0460_ _1550_ _1529_ _0469_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__4008__D net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_109_clk clknet_4_2_0_clk clknet_leaf_109_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_106_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_60_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3873__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ net522 clknet_leaf_1_clk hotp.block.sha1.mixer.w\[179\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3883_ net582 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[110\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2903_ _1181_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3847__D net796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2834_ _1590_ _0497_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_115_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_75_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2765_ _1076_ _1085_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2696_ hotp.digest\[22\] _1023_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1716_ seg.digit\[2\] _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1647_ _1417_ _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4435_ _0336_ clknet_leaf_92_clk hotp.block.mixer.msg\[147\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4366_ _0267_ clknet_leaf_73_clk hotp.block.mixer.msg\[78\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold483_I hotp.block.sha1.mixer.w\[91\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3317_ _0058_ clknet_leaf_41_clk stream.msg_buf\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4297_ _0198_ clknet_leaf_91_clk hotp.block.mixer.msg\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_13_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold748_I hotp.block.sha1.mixer.w\[239\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3248_ _0826_ _1386_ _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3179_ hotp.block.mixer.msg\[138\] hotp.block.mixer.msg\[139\] _1340_ _1344_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_28_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold580 hotp.block.sha1.mixer.w\[446\] net600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold591 stream.key_buf\[133\] net611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_92_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold92_I hotp.block.sha1.mixer.w\[498\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2550_ _0901_ _0845_ _0886_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_50_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2481_ _0838_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4220_ net452 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[447\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_52_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4151_ net240 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[378\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4082_ net561 clknet_leaf_33_clk hotp.block.sha1.mixer.w\[309\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3102_ _1300_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3033_ _1245_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1860__A2 _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3935_ net829 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[162\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3866_ net451 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[93\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2817_ _1115_ _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3797_ net103 clknet_leaf_105_clk hotp.block.sha1.mixer.w\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold698_I hotp.block.sha1.mixer.w\[441\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2748_ _1060_ _1051_ _1071_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_14_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2679_ _0991_ _1015_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4418_ _0319_ clknet_leaf_70_clk hotp.block.mixer.msg\[130\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4201__D net303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4349_ _0250_ clknet_leaf_84_clk hotp.block.mixer.msg\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_45_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_94_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3950__D net341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2355__S _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3720_ net667 clknet_leaf_87_clk hotp.block.sha1.mixer.d\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1981_ _1512_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_40_clk clknet_4_7_0_clk clknet_leaf_40_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3911__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3651_ net832 clknet_leaf_80_clk hotp.block.sha1.mixer.b\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2602_ hotp.digest\[14\] _0947_ _0917_ _0847_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3582_ _0155_ clknet_leaf_62_clk hotp.digest\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2533_ hotp.digest\[6\] _0886_ _0845_ _0847_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_12_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4021__D net533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2464_ hotp.stage\[2\] _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2395_ _0735_ _0762_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3860__D net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4203_ net236 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[430\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4134_ net401 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[361\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold279_I hotp.block.sha1.mixer.w\[78\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4065_ net71 clknet_leaf_20_clk hotp.block.sha1.mixer.w\[292\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3016_ hotp.block.mixer.msg\[67\] hotp.block.mixer.msg\[68\] _1251_ _1252_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold446_I hotp.block.sha1.mixer.w\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold613_I hotp.block.sha1.mixer.w\[445\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_clk clknet_4_5_0_clk clknet_leaf_31_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3918_ net289 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[145\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3849_ net113 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[76\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_76_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98_clk clknet_4_3_0_clk clknet_leaf_98_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4097__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3934__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_22_clk clknet_4_4_0_clk clknet_leaf_22_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3945__D net668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2180_ stream.msg_buf\[61\] stream.msg_buf\[62\] _0516_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_89_clk clknet_4_8_0_clk clknet_leaf_89_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3265__A1 _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1964_ _0439_ _0441_ _0442_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_13_clk clknet_4_3_0_clk clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3703_ net99 clknet_leaf_86_clk hotp.block.sha1.mixer.c\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3855__D net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1895_ _1615_ _0387_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3634_ net101 clknet_leaf_78_clk hotp.block.sha1.mixer.a\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3565_ _0138_ clknet_leaf_47_clk hotp.digest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2516_ hotp.digest\[1\] _0870_ _0871_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3496_ net89 clknet_leaf_27_clk stream.key_buf\[148\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2447_ _0776_ _0805_ stream.counter\[12\] _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2378_ _0745_ _0746_ _0747_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_71_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4117_ net193 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[344\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4048_ net308 clknet_leaf_17_clk hotp.block.sha1.mixer.w\[275\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold9 hotp.block.sha1.mixer.e\[9\] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_89_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1680_ _1441_ _1448_ _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_64_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold409 hotp.block.sha1.mixer.w\[220\] net429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3022__I1 hotp.block.mixer.msg\[71\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4262__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3350_ net820 clknet_leaf_47_clk stream.key_buf\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2301_ _0699_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_111_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3281_ _0022_ clknet_leaf_39_clk stream.msg_buf\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2232_ _1446_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2163_ stream.msg_buf\[53\] stream.msg_buf\[54\] _0587_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2094_ _0548_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold409_I hotp.block.sha1.mixer.w\[220\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2996_ hotp.block.mixer.msg\[59\] hotp.block.mixer.msg\[60\] _1239_ _1240_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1947_ _1563_ _1575_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1878_ _1543_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3617_ net815 clknet_leaf_75_clk hotp.block.sha1.mixer.a\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3548_ _0125_ clknet_leaf_42_clk stream.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold778_I hotp.block.sha1.mixer.w\[151\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3479_ net340 clknet_leaf_33_clk stream.key_buf\[131\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4135__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold18_I hotp.block.sha1.mixer.w\[198\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2850_ _1151_ _1154_ _0419_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1801_ hotp.block.magic.step\[2\] _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2781_ _1100_ _1101_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1732_ _1478_ _1493_ _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xhold206 hotp.block.sha1.mixer.w\[122\] net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1663_ stream.msg_state\[1\] _1432_ _1433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold217 hotp.block.sha1.mixer.w\[19\] net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4451_ _0351_ clknet_leaf_94_clk hotp.block.mixer.round\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_113_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold228 stream.key_buf\[37\] net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3402_ net207 clknet_leaf_38_clk stream.key_buf\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold239 hotp.block.sha1.mixer.d\[9\] net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4382_ _0283_ clknet_leaf_72_clk hotp.block.mixer.msg\[94\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3333_ _0074_ clknet_leaf_43_clk stream.msg_buf\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3264_ _1395_ _0368_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2215_ _1421_ _0628_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3195_ _1353_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2146_ _0578_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2077_ stream.msg_buf\[16\] stream.msg_buf\[17\] _0535_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2979_ _1230_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4204__D net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold773 hotp.block.sha1.mixer.w\[332\] net793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold762 stream.key_buf\[23\] net782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold740 hotp.block.sha1.mixer.w\[98\] net760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold751 hotp.block.sha1.mixer.w\[93\] net771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold784 stream.key_buf\[156\] net804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold795 hotp.block.sha1.mixer.a\[5\] net815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_86_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2247__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3675__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__D net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2361__A1 hotp.block.sha1.mixer.e\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2000_ _0465_ _0471_ _0476_ _0478_ _1562_ _1536_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XPHY_EDGE_ROW_11_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3951_ net410 clknet_leaf_1_clk hotp.block.sha1.mixer.w\[178\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2902_ _1186_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3882_ net759 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[109\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2833_ hotp.block.sha1.mixer.a_carry\[0\] _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2764_ _0831_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4024__D net764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1927__A1 _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1715_ seg.digit\[3\] _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2695_ _0850_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3863__D net503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1646_ _1414_ _1416_ _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4434_ _0335_ clknet_leaf_92_clk hotp.block.mixer.msg\[146\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4365_ _0266_ clknet_leaf_72_clk hotp.block.mixer.msg\[77\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3316_ _0057_ clknet_leaf_41_clk stream.msg_buf\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4296_ _0197_ clknet_leaf_91_clk hotp.block.mixer.msg\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3247_ _1377_ _1384_ _1386_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_hold643_I hotp.block.sha1.mixer.w\[154\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3178_ _1343_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2129_ _0568_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold810_I hotp.block.sha1.mixer.w\[168\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2530__I _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold570 stream.key_buf\[155\] net590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold581 hotp.block.sha1.mixer.w\[210\] net601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_92_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold592 hotp.block.sha1.mixer.w\[475\] net612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_9_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2906__S _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3948__D net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold85_I hotp.block.sha1.mixer.w\[96\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2480_ _0837_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4150_ net770 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[377\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3101_ hotp.block.mixer.msg\[104\] hotp.block.mixer.msg\[105\] _1298_ _1300_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4081_ net97 clknet_leaf_40_clk hotp.block.sha1.mixer.w\[308\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3032_ _1260_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4019__D net720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3858__D net447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3934_ net824 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[161\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_63_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold224_I hotp.block.sha1.mixer.w\[435\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3865_ net771 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[92\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2816_ _1127_ _1119_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3796_ net675 clknet_leaf_105_clk hotp.block.sha1.mixer.w\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2747_ hotp.digest\[30\] _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2678_ _1000_ _1010_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_hold593_I hotp.block.sha1.mixer.w\[232\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4417_ _0318_ clknet_leaf_71_clk hotp.block.mixer.msg\[129\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4348_ _0249_ clknet_leaf_84_clk hotp.block.mixer.msg\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3181__I _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4279_ net296 clknet_leaf_99_clk hotp.block.sha1.mixer.w\[506\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_94_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4219__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_74_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1980_ _0458_ _0443_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_89_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3650_ net273 clknet_leaf_79_clk hotp.block.sha1.mixer.b\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_12_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2601_ _0946_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3581_ _0154_ clknet_leaf_62_clk hotp.digest\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2532_ _0885_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_27_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2463_ _0813_ _0818_ _0820_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4202_ net361 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[429\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2394_ stream.counter\[3\] _0748_ _0751_ _0761_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4133_ net392 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[360\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_3_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4064_ net671 clknet_leaf_20_clk hotp.block.sha1.mixer.w\[291\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3015_ _1245_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold341_I hotp.block.sha1.mixer.w\[430\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold606_I hotp.block.sha1.mixer.w\[174\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3917_ net337 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[144\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ net635 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[75\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3779_ net557 clknet_leaf_100_clk hotp.block.sha1.mixer.w\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4212__D net629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3961__D net510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3265__A2 _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4191__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ hotp.block.mixer.round\[6\] _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_44_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1894_ _1616_ _0386_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_7_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3702_ net505 clknet_leaf_86_clk hotp.block.sha1.mixer.c\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3633_ net467 clknet_leaf_78_clk hotp.block.sha1.mixer.a\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4032__D net795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3564_ _0137_ clknet_leaf_47_clk hotp.digest\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3495_ net686 clknet_leaf_27_clk stream.key_buf\[147\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2515_ _0844_ _0869_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3871__D net485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2446_ _0797_ _0798_ _0738_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_58_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold389_I hotp.block.sha1.mixer.w\[188\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2377_ _0737_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_71_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4116_ net268 clknet_leaf_18_clk hotp.block.sha1.mixer.w\[343\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_3_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4047_ net47 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[274\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold723_I hotp.block.sha1.mixer.w\[394\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4207__D net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_58_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3956__D net492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3280_ _0021_ clknet_leaf_50_clk stream.msg_buf\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2300_ stream.digest\[6\] stream.digest\[7\] _0696_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_111_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_76_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2231_ _0635_ _0644_ _0629_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_111_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2162_ _0571_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2093_ stream.msg_buf\[23\] stream.msg_buf\[24\] _0545_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4027__D net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold137_I hotp.block.sha1.mixer.w\[64\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3866__D net451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2995_ _1223_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_44_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4087__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1946_ _0426_ hotp.block.sha1.mixer.w_fb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1877_ _0367_ _0368_ _0369_ _1531_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_9_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3616_ net825 clknet_leaf_75_clk hotp.block.sha1.mixer.a\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3547_ _0124_ clknet_leaf_42_clk stream.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3478_ net674 clknet_leaf_32_clk stream.key_buf\[130\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3924__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2429_ _0611_ _0787_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1800_ _1549_ _1553_ _1558_ _1542_ _1560_ _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_38_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2780_ stream.key_counter\[5\] _1098_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1731_ seg.digit\[2\] _1480_ _1492_ _1493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_54_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1662_ _1426_ _1431_ _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold207 hotp.block.sha1.mixer.w\[487\] net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4450_ _0350_ clknet_leaf_68_clk hotp.block.mixer.round\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_113_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3401_ net51 clknet_leaf_51_clk stream.key_buf\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4381_ _0282_ clknet_leaf_72_clk hotp.block.mixer.msg\[93\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold229 hotp.block.sha1.mixer.w\[241\] net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold218 hotp.block.sha1.mixer.w\[197\] net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XPHY_EDGE_ROW_84_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3332_ _0073_ clknet_leaf_43_clk stream.msg_buf\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3263_ hotp.stage\[2\] _1394_ _1396_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2214_ _0614_ _0627_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3194_ hotp.block.mixer.msg\[144\] hotp.block.mixer.msg\[145\] _1351_ _1353_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2145_ stream.msg_buf\[45\] stream.msg_buf\[46\] _0577_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_37_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2076_ _0538_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_93_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold519_I hotp.block.sha1.mixer.w\[356\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2978_ hotp.block.mixer.msg\[51\] hotp.block.mixer.msg\[52\] _1229_ _1230_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1929_ _1468_ _0409_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1945__A2 _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold730 hotp.block.sha1.mixer.w\[284\] net750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4220__D net452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold763 hotp.block.sha1.mixer.a\[6\] net783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold752 hotp.block.sha1.mixer.w\[372\] net772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold741 hotp.block.sha1.mixer.c\[11\] net761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold774 stream.key_buf\[115\] net794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold785 hotp.block.sha1.mixer.w\[164\] net805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold796 hotp.block.sha1.mixer.b\[2\] net816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4130__D net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold90 hotp.block.sha1.mixer.w\[80\] net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_26_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3950_ net341 clknet_leaf_1_clk hotp.block.sha1.mixer.w\[177\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2901_ hotp.block.mixer.msg\[18\] hotp.block.mixer.msg\[19\] _1182_ _1186_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3881_ net802 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[108\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2832_ hotp.block.sha1.mixer.a_carry\[0\] _0434_ _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2763_ _1090_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1714_ _1476_ _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2694_ hotp.digest\[24\] _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1645_ stream.state\[1\] _1415_ _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4433_ _0334_ clknet_leaf_93_clk hotp.block.mixer.msg\[145\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4364_ _0265_ clknet_leaf_73_clk hotp.block.mixer.msg\[76\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3315_ _0056_ clknet_leaf_34_clk stream.msg_buf\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4295_ _0196_ clknet_leaf_95_clk hotp.block.mixer.msg\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3246_ _1533_ _1385_ _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4275__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3177_ hotp.block.mixer.msg\[137\] hotp.block.mixer.msg\[138\] _1340_ _1343_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2128_ stream.msg_buf\[38\] stream.msg_buf\[39\] _0566_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2059_ _0528_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold803_I hotp.block.sha1.mixer.w\[388\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4215__D net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold560 hotp.block.sha1.mixer.w\[312\] net580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold571 hotp.block.sha1.mixer.w\[101\] net591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold582 stream.key_buf\[119\] net602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_92_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold593 hotp.block.sha1.mixer.w\[232\] net613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3642__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3964__D net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4148__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3100_ _1299_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4080_ net178 clknet_leaf_34_clk hotp.block.sha1.mixer.w\[307\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3031_ hotp.block.mixer.msg\[74\] hotp.block.mixer.msg\[75\] _1256_ _1260_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_108_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3933_ net369 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[160\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_63_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3864_ net696 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[91\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2815_ _1082_ hotp.digest\[32\] _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2631__I _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3795_ net403 clknet_leaf_105_clk hotp.block.sha1.mixer.w\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3874__D net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2746_ _1065_ _1074_ _1075_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2677_ _1006_ _1013_ _1014_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4416_ _0317_ clknet_leaf_71_clk hotp.block.mixer.msg\[128\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold753_I hotp.block.sha1.mixer.w\[130\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4347_ _0248_ clknet_leaf_84_clk hotp.block.mixer.msg\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4278_ net142 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[505\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3229_ _1371_ _1372_ _0503_ _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_30_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2013__A1 _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold390 hotp.block.sha1.mixer.w\[179\] net410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3959__D net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2600_ hotp.digest\[11\] hotp.digest\[12\] hotp.digest\[13\] _0946_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3580_ _0153_ clknet_leaf_62_clk hotp.digest\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2531_ hotp.digest\[3\] hotp.digest\[4\] hotp.digest\[5\] _0885_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2462_ _0819_ _1528_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4201_ net303 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[428\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2393_ _0607_ _0753_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4132_ net599 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[359\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_3_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4063_ net776 clknet_leaf_20_clk hotp.block.sha1.mixer.w\[290\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3014_ _1250_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3869__D net754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_hold334_I hotp.block.sha1.mixer.w\[369\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3916_ net499 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[143\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3847_ net796 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[74\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3778_ net504 clknet_leaf_100_clk hotp.block.sha1.mixer.w\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2729_ hotp.digest\[28\] _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output16_I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3830__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_4_7_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3360__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ _0440_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1893_ _1627_ _0373_ _0381_ _0385_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3701_ net723 clknet_leaf_86_clk hotp.block.sha1.mixer.c\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3025__I0 hotp.block.mixer.msg\[71\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3632_ net375 clknet_leaf_78_clk hotp.block.sha1.mixer.a\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_116_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3563_ _0136_ clknet_leaf_47_clk hotp.digest\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_51_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3494_ net83 clknet_leaf_28_clk stream.key_buf\[146\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2514_ _0843_ _0869_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2445_ _0602_ _0797_ _0780_ _0798_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2376_ _1453_ _0642_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_71_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4115_ net373 clknet_leaf_18_clk hotp.block.sha1.mixer.w\[342\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ net703 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[273\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_35_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3853__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_104_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_73_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4209__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_88_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_89_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_11_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2455__B2 _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_26_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3007__I0 hotp.block.mixer.msg\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4133__D net392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2230_ _1429_ _0643_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_111_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3726__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2161_ _0586_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2092_ _0547_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2994_ _1238_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_32_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1945_ hotp.block.debug\[1\] _0425_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1876_ _1624_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_44_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3615_ net799 clknet_leaf_76_clk hotp.block.sha1.mixer.a\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3546_ _0123_ clknet_leaf_42_clk stream.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3477_ net269 clknet_leaf_29_clk stream.key_buf\[129\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2428_ _0786_ _0752_ _0781_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2359_ _0396_ _0686_ _0688_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4218__D net600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4029_ net363 clknet_leaf_13_clk hotp.block.sha1.mixer.w\[256\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4031__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3967__D net545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1730_ seg.digit\[1\] _1483_ _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1661_ _1427_ _1430_ _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold208 hotp.block.sha1.mixer.w\[102\] net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3400_ net677 clknet_leaf_51_clk stream.key_buf\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold219 hotp.block.sha1.mixer.w\[452\] net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4380_ _0281_ clknet_leaf_72_clk hotp.block.mixer.msg\[92\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3331_ _0072_ clknet_leaf_40_clk stream.msg_buf\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3262_ hotp.stage\[2\] _1394_ _0684_ _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input7_I in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2213_ _0511_ _0623_ _0625_ _0626_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3193_ _1352_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2144_ _0571_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4038__D net558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2075_ stream.msg_buf\[15\] stream.msg_buf\[16\] _0535_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1890__A2 _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3877__D net478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold247_I hotp.block.sha1.mixer.w\[424\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold414_I hotp.block.sha1.mixer.w\[426\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2977_ _1223_ _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_86_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1928_ _1424_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1859_ _1604_ _1618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold720 hotp.block.sha1.mixer.w\[494\] net740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_hold783_I hotp.block.sha1.mixer.w\[466\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold731 stream.key_buf\[70\] net751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold764 hotp.block.sha1.mixer.w\[159\] net784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold753 hotp.block.sha1.mixer.w\[130\] net773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold742 hotp.block.sha1.mixer.w\[373\] net762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold797 stream.key_buf\[101\] net817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold786 hotp.block.sha1.mixer.w\[277\] net806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3529_ _0106_ clknet_leaf_16_clk stream.digest\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold775 hotp.block.sha1.mixer.w\[260\] net795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_12_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_15_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1713__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1936__A3 _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold23_I hotp.block.sha1.mixer.w\[386\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold91 hotp.block.sha1.mixer.w\[450\] net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold80 hotp.block.sha1.mixer.w\[367\] net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_106_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2900_ _1185_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3880_ net706 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[107\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_70_clk clknet_4_11_0_clk clknet_leaf_70_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2831_ _1137_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2762_ _1089_ _1076_ _0838_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1713_ net7 _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2693_ _1006_ _1026_ _1028_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4432_ _0333_ clknet_leaf_93_clk hotp.block.mixer.msg\[144\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1644_ stream.debug\[1\] _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_22_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4363_ _0264_ clknet_leaf_73_clk hotp.block.mixer.msg\[75\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3314_ _0055_ clknet_leaf_40_clk stream.msg_buf\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4294_ _0195_ clknet_leaf_104_clk hotp.block.mixer.msg\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3245_ _1106_ _0430_ _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3176_ _1342_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2127_ _0567_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_68_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1863__A2 _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2058_ stream.msg_buf\[8\] stream.msg_buf\[9\] _0524_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold531_I hotp.block.sha1.mixer.w\[136\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold629_I hotp.block.sha1.mixer.w\[371\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2364__I _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_81_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_61_clk clknet_4_14_0_clk clknet_leaf_61_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4231__D net497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold550 hotp.block.sha1.mixer.w\[406\] net570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold572 hotp.block.sha1.mixer.w\[399\] net592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold561 hotp.block.sha1.mixer.d\[21\] net581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_102_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold594 hotp.block.sha1.mixer.w\[268\] net614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold583 hotp.block.sha1.mixer.w\[408\] net603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_92_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3937__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_52_clk clknet_4_13_0_clk clknet_leaf_52_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4141__D net354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3980__D net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3030_ _1259_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43_clk clknet_4_6_0_clk clknet_leaf_43_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3932_ net641 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[159\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_63_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3863_ net503 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[90\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2814_ _1117_ _1119_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3794_ net672 clknet_leaf_105_clk hotp.block.sha1.mixer.w\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2745_ _1060_ _1058_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2676_ _1000_ _0998_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4415_ _0316_ clknet_leaf_71_clk hotp.block.mixer.msg\[127\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4242__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold579_I hotp.block.sha1.mixer.w\[360\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold481_I hotp.block.sha1.mixer.w\[230\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4346_ _0247_ clknet_leaf_83_clk hotp.block.mixer.msg\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4277_ net346 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[504\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3228_ hotp.block.mixer.msg\[159\] _1611_ _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_hold746_I hotp.block.sha1.mixer.w\[149\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3159_ hotp.block.mixer.msg\[129\] hotp.block.mixer.msg\[130\] _1330_ _1333_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_25_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_34_clk clknet_4_7_0_clk clknet_leaf_34_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1772__A1 _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold380 stream.key_buf\[142\] net400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold391 hotp.block.sha1.mixer.w\[214\] net411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4136__D net625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_25_clk clknet_4_4_0_clk clknet_leaf_25_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_hold90_I hotp.block.sha1.mixer.w\[80\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3975__D net609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4265__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_3_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2530_ _0883_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2461_ _1510_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4200_ net119 clknet_leaf_11_clk hotp.block.sha1.mixer.w\[427\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2392_ _0619_ _0606_ stream.counter\[3\] _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4131_ net114 clknet_leaf_9_clk hotp.block.sha1.mixer.w\[358\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_3_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4062_ net412 clknet_leaf_20_clk hotp.block.sha1.mixer.w\[289\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3268__A1 _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3013_ hotp.block.mixer.msg\[66\] hotp.block.mixer.msg\[67\] _1246_ _1250_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1818__A2 _1578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_clk clknet_4_6_0_clk clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3915_ net747 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[142\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3846_ net257 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[73\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3777_ net586 clknet_leaf_100_clk hotp.block.sha1.mixer.w\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2728_ _1035_ _1057_ _1059_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2659_ hotp.digest\[18\] _0998_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3782__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4329_ _0230_ clknet_leaf_89_clk hotp.block.mixer.msg\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4138__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ net280 clknet_leaf_85_clk hotp.block.sha1.mixer.c\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1961_ hotp.block.mixer.round\[3\] hotp.block.mixer.round\[5\] hotp.block.mixer.round\[4\]
+ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_60_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1892_ _1610_ _0383_ _0384_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3631_ net496 clknet_leaf_78_clk hotp.block.sha1.mixer.a\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3025__I1 hotp.block.mixer.msg\[72\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3562_ _0135_ clknet_leaf_47_clk hotp.digest\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_116_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2513_ _0848_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3493_ net347 clknet_leaf_28_clk stream.key_buf\[145\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2444_ _0646_ _0803_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_58_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_5_clk clknet_4_1_0_clk clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2375_ _0739_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_71_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4114_ net800 clknet_leaf_18_clk hotp.block.sha1.mixer.w\[341\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4045_ net618 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[272\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold709_I hotp.block.sha1.mixer.b\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3829_ net474 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_13_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold53_I hotp.block.sha1.mixer.w\[140\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ stream.msg_buf\[52\] stream.msg_buf\[53\] _0582_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4453__CLK clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2091_ stream.msg_buf\[22\] stream.msg_buf\[23\] _0545_ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2993_ hotp.block.mixer.msg\[58\] hotp.block.mixer.msg\[59\] _1234_ _1238_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_32_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1944_ hotp.block.sha1.mixer.w\[64\] hotp.block.sha1.mixer.w\[256\] hotp.block.sha1.mixer.w\[416\]
+ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1875_ _1552_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3614_ net162 clknet_leaf_77_clk hotp.block.sha1.mixer.a\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3545_ _0122_ clknet_leaf_42_clk stream.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3476_ net150 clknet_leaf_32_clk stream.key_buf\[128\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2427_ _0788_ _0789_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2358_ _0731_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2289_ stream.digest\[1\] stream.digest\[2\] _0691_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4028_ net834 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[255\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_84_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_11_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4234__D net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__D net772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3983__D net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1660_ _1428_ stream.msg_state\[0\] _1429_ _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_0_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold209 hotp.block.sha1.mixer.c\[20\] net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_33_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3330_ _0071_ clknet_leaf_39_clk stream.msg_buf\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3261_ _1618_ _1392_ _1394_ _1395_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2212_ _0624_ _0508_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3192_ hotp.block.mixer.msg\[143\] hotp.block.mixer.msg\[144\] _1351_ _1352_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3843__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2143_ _0576_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2074_ _0537_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_72_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_87_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2976_ _1228_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ _1442_ _0408_ _0411_ stream.key_buf\[0\] _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_72_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1858_ _1497_ _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_10_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold710 hotp.block.sha1.mixer.w\[113\] net730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold721 hotp.block.sha1.mixer.a\[7\] net741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold743 hotp.block.sha1.mixer.w\[129\] net763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold754 hotp.block.sha1.mixer.a\[8\] net774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold732 hotp.block.sha1.mixer.w\[478\] net752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_hold776_I hotp.block.sha1.mixer.w\[75\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1789_ hotp.block.magic.step\[0\] _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold787 hotp.block.sha1.mixer.w\[119\] net807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3528_ _0105_ clknet_leaf_16_clk stream.digest\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold765 hotp.block.sha1.mixer.w\[221\] net785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold776 hotp.block.sha1.mixer.w\[75\] net796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold798 stream.key_buf\[67\] net818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3459_ net585 clknet_leaf_31_clk stream.key_buf\[111\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_25_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_23_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_97_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold16_I hotp.block.sha1.mixer.w\[88\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4139__D net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold70 stream.key_buf\[110\] net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold92 hotp.block.sha1.mixer.w\[498\] net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold81 hotp.block.sha1.mixer.a\[22\] net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3978__D net323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2830_ hotp.digest\[39\] _0857_ _1129_ hotp.digest\[38\] _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3396__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2761_ _1082_ _1088_ _0831_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2692_ hotp.digest\[22\] _1027_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1712_ hotp.block.debug\[0\] _1475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1643_ stream.state\[2\] _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_1 net481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4431_ _0332_ clknet_leaf_93_clk hotp.block.mixer.msg\[143\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4362_ _0263_ clknet_leaf_73_clk hotp.block.mixer.msg\[74\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3313_ _0054_ clknet_leaf_34_clk stream.msg_buf\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4293_ _0194_ clknet_leaf_100_clk hotp.block.mixer.msg\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3244_ _1517_ _1383_ _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4021__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3175_ hotp.block.mixer.msg\[136\] hotp.block.mixer.msg\[137\] _1340_ _1342_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2126_ stream.msg_buf\[37\] stream.msg_buf\[38\] _0566_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_68_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2057_ _0527_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2959_ hotp.block.mixer.msg\[43\] hotp.block.mixer.msg\[44\] _1218_ _1219_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold551 stream.key_buf\[117\] net571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold562 hotp.block.sha1.mixer.w\[111\] net582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_60_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold540 hotp.block.sha1.mixer.w\[395\] net560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold595 stream.key_buf\[84\] net615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_92_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold573 hotp.block.sha1.mixer.w\[377\] net593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold584 hotp.block.sha1.mixer.e\[22\] net604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_92_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2500__A1 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1854__A3 _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2567__A1 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1917__I1 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4194__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3931_ net784 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[158\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3862_ net293 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[89\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2813_ _1125_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3793_ net469 clknet_leaf_105_clk hotp.block.sha1.mixer.w\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2744_ _1066_ _0842_ _1073_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2675_ hotp.digest\[21\] _0915_ _1010_ _1012_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_78_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4414_ _0315_ clknet_leaf_71_clk hotp.block.mixer.msg\[126\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4345_ _0246_ clknet_leaf_83_clk hotp.block.mixer.msg\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4276_ net624 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[503\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3227_ _1158_ _1607_ _1608_ _1611_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_118_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3158_ _1332_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2109_ _0557_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3089_ _1287_ _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4242__D net808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold381 hotp.block.sha1.mixer.w\[362\] net401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold370 hotp.block.sha1.mixer.w\[191\] net390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_99_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold392 hotp.block.sha1.mixer.w\[290\] net412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4152__D net694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3991__D net374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2460_ _1517_ _0817_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2391_ _0756_ _0758_ _0759_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4130_ net95 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[357\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4061_ net546 clknet_leaf_19_clk hotp.block.sha1.mixer.w\[288\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3012_ _1249_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_65_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3914_ net605 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[141\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3020__S _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold222_I hotp.block.sha1.mixer.w\[192\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3845_ net28 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[72\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3776_ net656 clknet_leaf_100_clk hotp.block.sha1.mixer.w\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2727_ hotp.digest\[26\] _1058_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2658_ _0856_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2589_ _0875_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4328_ _0229_ clknet_leaf_89_clk hotp.block.mixer.msg\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4259_ net227 clknet_leaf_100_clk hotp.block.sha1.mixer.w\[486\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3259__A2 _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4237__D net339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4147__D net835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3986__D net411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1960_ hotp.block.mixer.round\[3\] hotp.block.mixer.round\[2\] hotp.block.mixer.round\[5\]
+ hotp.block.mixer.round\[4\] _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_60_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1891_ _1555_ _1619_ _0374_ _1587_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_16_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3630_ net33 clknet_leaf_77_clk hotp.block.sha1.mixer.a\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3561_ _0134_ clknet_leaf_47_clk hotp.digest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_116_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2512_ _0861_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3492_ stream.key_buf\[145\] clknet_leaf_26_clk stream.key_buf\[144\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2443_ _0797_ _0749_ _0802_ _0408_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2374_ _0735_ _0744_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_71_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4113_ net312 clknet_leaf_19_clk hotp.block.sha1.mixer.w\[340\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold172_I hotp.block.sha1.mixer.w\[176\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4044_ net756 clknet_leaf_22_clk hotp.block.sha1.mixer.w\[271\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3828_ net589 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3759_ net579 clknet_leaf_79_clk hotp.block.sha1.mixer.e\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_18_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_89_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_27_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2090_ _0546_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_45_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2992_ _1237_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1943_ _0424_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1874_ _1555_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_54_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3613_ net218 clknet_leaf_76_clk hotp.block.debug\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4128__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3544_ _0121_ clknet_leaf_43_clk stream.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3475_ net440 clknet_leaf_32_clk stream.key_buf\[127\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold387_I hotp.block.sha1.mixer.w\[141\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2426_ _0786_ _0781_ _0413_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4278__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2357_ stream.digest\[31\] _0403_ _0727_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2288_ _0692_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold554_I hotp.block.sha1.mixer.w\[409\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4027_ net91 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[254\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_84_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_72_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4160__D net823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3260_ _0684_ _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2211_ _0400_ _0624_ _1416_ _1444_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_3191_ _1350_ _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2142_ stream.msg_buf\[44\] stream.msg_buf\[45\] _0572_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2073_ stream.msg_buf\[14\] stream.msg_buf\[15\] _0535_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold135_I hotp.block.sha1.mixer.w\[472\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2975_ hotp.block.mixer.msg\[50\] hotp.block.mixer.msg\[51\] _1224_ _1228_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1926_ _1404_ _1410_ _0410_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1857_ _1605_ hotp.block.main_in _1616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold711 hotp.block.sha1.mixer.d\[18\] net731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold700 hotp.block.sha1.mixer.w\[247\] net720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold733 hotp.block.sha1.mixer.w\[324\] net753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3527_ _0104_ clknet_leaf_16_clk stream.digest\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1788_ _1539_ _1549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold722 hotp.block.sha1.mixer.w\[27\] net742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold755 hotp.block.sha1.mixer.w\[200\] net775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold744 hotp.block.sha1.mixer.w\[252\] net764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_hold671_I hotp.block.sha1.mixer.w\[442\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold766 hotp.block.sha1.mixer.w\[172\] net786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold777 hotp.block.sha1.mixer.w\[421\] net797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold788 hotp.block.sha1.mixer.w\[470\] net808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3458_ net76 clknet_leaf_34_clk stream.key_buf\[110\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold799 hotp.block.sha1.mixer.w\[244\] net819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3389_ net253 clknet_leaf_54_clk stream.key_buf\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2409_ _0400_ _0765_ _0753_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_93_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4245__D net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold60 hotp.block.sha1.mixer.w\[327\] net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_89_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold82 hotp.block.sha1.mixer.w\[170\] net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold71 hotp.block.sha1.mixer.w\[255\] net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_89_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold93 hotp.block.sha1.mixer.w\[77\] net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4155__D net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3994__D net714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2760_ _1592_ _0841_ _1087_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1711_ _1434_ _1474_ _1425_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2691_ _0856_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1642_ _1403_ _1412_ _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_2 hotp.block.sha1.mixer.w\[151\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4430_ _0331_ clknet_leaf_69_clk hotp.block.mixer.msg\[142\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4361_ _0262_ clknet_leaf_74_clk hotp.block.mixer.msg\[73\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3312_ _0053_ clknet_leaf_34_clk stream.msg_buf\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4292_ _0193_ clknet_leaf_100_clk hotp.block.mixer.msg\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3243_ _1377_ _1382_ _1383_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3174_ _1341_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2125_ _0550_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1830__I hotp.block.sha1.mixer.e\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2056_ stream.msg_buf\[7\] stream.msg_buf\[8\] _0524_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_68_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold252_I hotp.block.sha1.mixer.w\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2273__A1 hotp.block.main_in vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold517_I hotp.block.sha1.mixer.w\[213\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2958_ _1202_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1909_ _0396_ _1477_ _0398_ net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_20_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2889_ hotp.block.mixer.msg\[13\] hotp.block.mixer.msg\[14\] _1176_ _1179_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold530 stream.key_buf\[89\] net550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold552 stream.key_buf\[125\] net572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold541 hotp.block.sha1.mixer.w\[310\] net561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold563 hotp.block.sha1.mixer.w\[449\] net583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold596 stream.key_buf\[58\] net616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold574 hotp.block.sha1.mixer.w\[157\] net594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold585 hotp.block.sha1.mixer.w\[142\] net605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_92_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3833__CLK clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_71_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_86_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3989__D net554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_47_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3930_ net264 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[157\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3861_ net305 clknet_leaf_6_clk hotp.block.sha1.mixer.w\[88\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2812_ hotp.digest\[33\] _1122_ _1116_ _1124_ _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_63_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3792_ net536 clknet_leaf_105_clk hotp.block.sha1.mixer.w\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2743_ _1051_ _1071_ _1072_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2414__C _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_39_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2674_ _0980_ _1011_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4413_ _0314_ clknet_leaf_71_clk hotp.block.mixer.msg\[125\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3018__S _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4344_ _0245_ clknet_leaf_83_clk hotp.block.mixer.msg\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4275_ net588 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[502\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3706__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3226_ _1370_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3157_ hotp.block.mixer.msg\[128\] hotp.block.mixer.msg\[129\] _1330_ _1332_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2108_ stream.msg_buf\[29\] stream.msg_buf\[30\] _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3088_ _1292_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_25_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2039_ _0516_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_25_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3856__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_111_clk clknet_4_0_0_clk clknet_leaf_111_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold371 stream.key_buf\[2\] net391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold360 hotp.block.sha1.mixer.d\[19\] net380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold393 stream.key_buf\[106\] net413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold382 hotp.block.sha1.mixer.w\[85\] net402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_99_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_102_clk clknet_4_2_0_clk clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_118_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2390_ _1446_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3729__CLK clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4060_ net367 clknet_leaf_19_clk hotp.block.sha1.mixer.w\[287\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3011_ hotp.block.mixer.msg\[65\] hotp.block.mixer.msg\[66\] _1246_ _1249_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3913_ net407 clknet_leaf_8_clk hotp.block.sha1.mixer.w\[140\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3844_ net284 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[71\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3775_ net243 clknet_leaf_99_clk hotp.block.sha1.mixer.w\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2726_ _0856_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2657_ _0990_ _0985_ _0996_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_76_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2588_ _0930_ _0898_ _0935_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4327_ _0228_ clknet_leaf_89_clk hotp.block.mixer.msg\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold751_I hotp.block.sha1.mixer.w\[93\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4258_ net199 clknet_leaf_99_clk hotp.block.sha1.mixer.w\[485\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3209_ _1350_ _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_97_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4189_ net168 clknet_leaf_101_clk hotp.block.sha1.mixer.w\[416\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4184__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold190 hotp.block.sha1.mixer.b\[5\] net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3401__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4163__D net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1890_ _0382_ _1551_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3560_ _0007_ clknet_leaf_46_clk stream.key_state\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_116_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2511_ hotp.digest\[3\] _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3491_ net744 clknet_leaf_26_clk stream.key_buf\[143\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3507__D _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2442_ _0797_ _0799_ _0801_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2373_ _0737_ _0743_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4112_ net345 clknet_leaf_19_clk hotp.block.sha1.mixer.w\[339\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4043_ net170 clknet_leaf_14_clk hotp.block.sha1.mixer.w\[270\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_hold165_I hotp.block.sha1.mixer.w\[166\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3031__S _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3827_ net330 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3758_ net356 clknet_leaf_81_clk hotp.block.sha1.mixer.e\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2709_ _0980_ _1042_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3689_ net487 clknet_leaf_83_clk hotp.block.sha1.mixer.c\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4248__D net408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output14_I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3997__D net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2991_ hotp.block.mixer.msg\[57\] hotp.block.mixer.msg\[58\] _1234_ _1237_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1942_ hotp.block.sha1.mixer.t _0388_ _1531_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_32_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1873_ _1505_ _1606_ _1629_ _0365_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3612_ _0185_ clknet_leaf_47_clk hotp.digest\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3543_ _0120_ clknet_leaf_97_clk hotp.block.sha1.mixer.h_carry vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3474_ net491 clknet_leaf_32_clk stream.key_buf\[126\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2425_ _0786_ _0776_ _0780_ _0787_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_50_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold282_I hotp.block.sha1.mixer.w\[182\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2356_ _0730_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2287_ stream.digest\[0\] stream.digest\[1\] _0691_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4026_ net461 clknet_leaf_5_clk hotp.block.sha1.mixer.w\[253\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_91_clk clknet_4_8_0_clk clknet_leaf_91_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4222__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_18_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_82_clk clknet_4_10_0_clk clknet_leaf_82_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1653__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2210_ stream.state\[2\] _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_55_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3190_ _1159_ _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2141_ _0575_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2072_ _0536_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_73_clk clknet_4_11_0_clk clknet_leaf_73_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2974_ _1227_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1925_ _1455_ _0409_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold128_I hotp.block.sha1.mixer.w\[438\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1828__I _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1856_ _1609_ _1614_ _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold712 hotp.block.sha1.mixer.w\[298\] net732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1787_ _1545_ _1547_ _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_12_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold701 hotp.block.sha1.mixer.d\[30\] net721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4245__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3526_ _0103_ clknet_leaf_15_clk stream.digest\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold723 hotp.block.sha1.mixer.w\[394\] net743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold734 hotp.block.sha1.mixer.w\[97\] net754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold745 hotp.block.sha1.mixer.e\[31\] net765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold756 hotp.block.sha1.mixer.w\[291\] net776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold778 hotp.block.sha1.mixer.w\[151\] net798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold767 hotp.block.sha1.mixer.w\[147\] net787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3457_ net90 clknet_leaf_31_clk stream.key_buf\[109\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold789 hotp.block.sha1.mixer.w\[47\] net809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3388_ net736 clknet_leaf_54_clk stream.key_buf\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2408_ _0773_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2339_ stream.digest\[23\] stream.digest\[24\] _0717_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4009_ net527 clknet_leaf_3_clk hotp.block.sha1.mixer.w\[236\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_64_clk clknet_4_15_0_clk clknet_leaf_64_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1738__I _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold50 hotp.block.sha1.mixer.w\[339\] net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1857__A2 hotp.block.main_in vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold61 hotp.block.sha1.mixer.w\[329\] net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold72 hotp.block.sha1.mixer.w\[500\] net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold83 hotp.block.sha1.mixer.w\[25\] net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold94 hotp.block.sha1.mixer.w\[359\] net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55_clk clknet_4_13_0_clk clknet_leaf_55_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4268__CLK clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1710_ _1453_ _1473_ stream.msg_state\[0\] _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2690_ _1019_ _1020_ _1025_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1641_ _1404_ _1405_ _1411_ _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_3 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ _0261_ clknet_leaf_75_clk hotp.block.mixer.msg\[72\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3311_ _0052_ clknet_leaf_34_clk stream.msg_buf\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4291_ _0192_ clknet_leaf_95_clk hotp.block.mixer.msg\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3242_ _1628_ _0397_ _1378_ _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_input5_I in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3173_ hotp.block.mixer.msg\[135\] hotp.block.mixer.msg\[136\] _1340_ _1341_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2124_ _0565_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_68_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2055_ _0526_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_46_clk clknet_4_12_0_clk clknet_leaf_46_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold245_I hotp.block.sha1.mixer.w\[183\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1759__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2957_ _1217_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1908_ _0397_ _1602_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_20_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2888_ _1178_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1839_ _1596_ _1598_ _1599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold520 hotp.block.sha1.mixer.e\[8\] net540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold542 stream.key_buf\[35\] net562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold531 hotp.block.sha1.mixer.w\[136\] net551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_60_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold553 hotp.block.sha1.mixer.w\[467\] net573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold597 stream.key_buf\[52\] net617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3509_ _0086_ clknet_leaf_66_clk hotp.rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold564 hotp.block.sha1.mixer.w\[35\] net584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold575 hotp.block.sha1.mixer.w\[40\] net595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold586 hotp.block.sha1.mixer.b\[31\] net606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_37_clk clknet_4_7_0_clk clknet_leaf_37_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold21_I hotp.block.sha1.mixer.w\[259\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_90_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_28_clk clknet_4_5_0_clk clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4166__D net743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4090__CLK clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3860_ net36 clknet_leaf_2_clk hotp.block.sha1.mixer.w\[87\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2811_ hotp.digest\[32\] _1123_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3791_ net237 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2742_ _1050_ _1071_ _0830_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2673_ _0990_ _1009_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4412_ _0313_ clknet_leaf_62_clk hotp.block.mixer.msg\[124\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1781__A4 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4343_ _0244_ clknet_leaf_83_clk hotp.block.mixer.msg\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold195_I hotp.block.sha1.mixer.w\[392\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4274_ net85 clknet_leaf_102_clk hotp.block.sha1.mixer.w\[501\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3225_ hotp.block.mixer.msg\[158\] hotp.block.mixer.msg\[159\] _1366_ _1370_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3261__C _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3156_ _1331_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4433__CLK clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2107_ _0550_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_77_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_19_clk clknet_4_6_0_clk clknet_leaf_19_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3087_ hotp.block.mixer.msg\[98\] hotp.block.mixer.msg\[99\] _1288_ _1292_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2038_ _0515_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_25_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3989_ net554 clknet_leaf_114_clk hotp.block.sha1.mixer.w\[216\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold361 stream.key_buf\[80\] net381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_7_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold350 hotp.block.sha1.mixer.w\[169\] net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold372 hotp.block.sha1.mixer.w\[361\] net392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold383 hotp.block.sha1.mixer.w\[23\] net403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold394 hotp.block.sha1.mixer.a\[17\] net414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_5_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_68_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1996__A1 _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold69_I stream.key_buf\[149\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1748__A1 _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3010_ _1248_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3912_ net73 clknet_leaf_24_clk hotp.block.sha1.mixer.w\[139\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3843_ net685 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[70\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold110_I hotp.block.sha1.mixer.w\[451\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3774_ net211 clknet_leaf_100_clk hotp.block.sha1.mixer.w\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2725_ _1051_ _1020_ _1056_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold208_I hotp.block.sha1.mixer.w\[102\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3029__S _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2656_ _0991_ _0995_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_8_clk clknet_4_1_0_clk clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2587_ _0909_ _0934_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3272__B _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4326_ _0227_ clknet_leaf_89_clk hotp.block.mixer.msg\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4257_ net385 clknet_leaf_99_clk hotp.block.sha1.mixer.w\[484\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold744_I hotp.block.sha1.mixer.w\[252\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3208_ _1360_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4188_ hotp.block.sha1.mixer.w\[416\] clknet_leaf_101_clk hotp.block.sha1.mixer.w\[415\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3139_ _1321_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_70_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_85_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold180 hotp.block.sha1.mixer.w\[181\] net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold191 hotp.block.sha1.mixer.w\[2\] net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_23_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_38_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3490_ net716 clknet_leaf_26_clk stream.key_buf\[142\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2510_ _0839_ _0865_ _0866_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2441_ _0603_ _0800_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3846__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2372_ stream.counter\[0\] _0738_ _0742_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4111_ net70 clknet_leaf_21_clk hotp.block.sha1.mixer.w\[338\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4042_ net52 clknet_leaf_10_clk hotp.block.sha1.mixer.w\[269\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3826_ net270 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3267__B _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3757_ net159 clknet_leaf_80_clk hotp.block.sha1.mixer.e\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2708_ _1019_ _1040_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold694_I hotp.block.sha1.mixer.w\[222\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3688_ net432 clknet_leaf_82_clk hotp.block.sha1.mixer.c\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2639_ _0959_ _0978_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4309_ _0210_ clknet_leaf_105_clk hotp.block.mixer.msg\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4151__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3399__CLK clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2990_ _1236_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1941_ _0416_ _0421_ _0423_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1872_ _0364_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3611_ _0184_ clknet_leaf_45_clk hotp.digest\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3542_ _0119_ clknet_leaf_66_clk stream.ready vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3473_ net453 clknet_leaf_32_clk stream.key_buf\[125\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2424_ _0786_ _0781_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2355_ stream.digest\[30\] stream.digest\[31\] _0727_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4024__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2286_ _0690_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_88_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4025_ net23 clknet_leaf_4_clk hotp.block.sha1.mixer.w\[252\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold707_I hotp.block.sha1.mixer.w\[393\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3809_ net698 clknet_leaf_112_clk hotp.block.sha1.mixer.w\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4169__D net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4197__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ stream.msg_buf\[43\] stream.msg_buf\[44\] _0572_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2071_ stream.msg_buf\[13\] stream.msg_buf\[14\] _0535_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2973_ hotp.block.mixer.msg\[49\] hotp.block.mixer.msg\[50\] _1224_ _1227_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1924_ stream.key_state\[3\] _1403_ _1409_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_8_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1855_ _1612_ _1613_ _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold702 stream.key_buf\[124\] net722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1786_ _1546_ _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold724 stream.key_buf\[144\] net744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3525_ _0102_ clknet_leaf_15_clk stream.digest\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold746 hotp.block.sha1.mixer.w\[149\] net766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold713 hotp.block.sha1.mixer.w\[366\] net733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold735 hotp.block.sha1.mixer.b\[29\] net755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold757 hotp.block.sha1.mixer.w\[123\] net777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold768 hotp.block.sha1.mixer.w\[238\] net788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold779 hotp.block.sha1.mixer.a\[3\] net799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3456_ net74 clknet_leaf_34_clk stream.key_buf\[108\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_110_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3387_ net726 clknet_leaf_54_clk stream.key_buf\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2407_ _0676_ _0747_ _0772_ _1425_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2338_ _0720_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2269_ stream.counter\[5\] _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4008_ net189 clknet_leaf_111_clk hotp.block.sha1.mixer.w\[235\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3907__CLK clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold40 hotp.block.sha1.mixer.w\[474\] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold62 stream.key_buf\[91\] net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold51 hotp.block.sha1.mixer.w\[293\] net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold73 hotp.block.sha1.mixer.w\[107\] net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold84 hotp.block.sha1.mixer.w\[463\] net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold95 hotp.block.sha1.mixer.e\[28\] net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold99_I hotp.block.sha1.mixer.w\[428\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1640_ _1410_ _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_4 net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3310_ _0051_ clknet_leaf_34_clk stream.msg_buf\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4290_ _0191_ clknet_leaf_95_clk hotp.block.mixer.msg\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3241_ _1628_ _1378_ _0397_ _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3172_ _1329_ _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2123_ stream.msg_buf\[36\] stream.msg_buf\[37\] _0561_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2054_ stream.msg_buf\[6\] stream.msg_buf\[7\] _0524_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4212__CLK clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold238_I hotp.block.sha1.mixer.w\[95\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2956_ hotp.block.mixer.msg\[42\] hotp.block.mixer.msg\[43\] _1213_ _1217_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1907_ _1518_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2887_ hotp.block.mixer.msg\[12\] hotp.block.mixer.msg\[13\] _1176_ _1178_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1838_ _1484_ _1493_ _1597_ _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_96_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold510 hotp.block.sha1.mixer.w\[235\] net530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold543 hotp.block.sha1.mixer.w\[454\] net563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1769_ _1529_ _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold521 hotp.block.sha1.mixer.w\[404\] net541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold554 hotp.block.sha1.mixer.w\[409\] net574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold532 hotp.block.sha1.mixer.b\[25\] net552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold565 stream.key_buf\[112\] net585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold587 stream.key_buf\[108\] net607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold576 hotp.block.sha1.mixer.w\[139\] net596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3508_ _0085_ clknet_leaf_45_clk hotp.block.main_in vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3439_ net418 clknet_leaf_31_clk stream.key_buf\[91\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold598 hotp.block.sha1.mixer.w\[273\] net618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_57_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4272__D net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4182__D net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2810_ hotp.digest\[31\] _1119_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3790_ net734 clknet_leaf_103_clk hotp.block.sha1.mixer.w\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2741_ _1070_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2672_ hotp.digest\[19\] _1009_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4411_ _0312_ clknet_leaf_62_clk hotp.block.mixer.msg\[123\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4342_ _0243_ clknet_leaf_83_clk hotp.block.mixer.msg\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4273_ net67 clknet_leaf_12_clk hotp.block.sha1.mixer.w\[500\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3224_ _1369_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
.ends

