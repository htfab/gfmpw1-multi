magic
tech gf180mcuD
magscale 1 10
timestamp 1702452663
<< metal1 >>
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 1344 55466 58576 55500
rect 1344 55414 4478 55466
rect 4530 55414 4582 55466
rect 4634 55414 4686 55466
rect 4738 55414 35198 55466
rect 35250 55414 35302 55466
rect 35354 55414 35406 55466
rect 35458 55414 58576 55466
rect 1344 55380 58576 55414
rect 1344 54458 58576 54492
rect 1344 54406 19838 54458
rect 19890 54406 19942 54458
rect 19994 54406 20046 54458
rect 20098 54406 50558 54458
rect 50610 54406 50662 54458
rect 50714 54406 50766 54458
rect 50818 54406 58576 54458
rect 1344 54372 58576 54406
rect 3838 54178 3890 54190
rect 3838 54114 3890 54126
rect 56030 54178 56082 54190
rect 56030 54114 56082 54126
rect 1344 53450 58576 53484
rect 1344 53398 4478 53450
rect 4530 53398 4582 53450
rect 4634 53398 4686 53450
rect 4738 53398 35198 53450
rect 35250 53398 35302 53450
rect 35354 53398 35406 53450
rect 35458 53398 58576 53450
rect 1344 53364 58576 53398
rect 1344 52442 58576 52476
rect 1344 52390 19838 52442
rect 19890 52390 19942 52442
rect 19994 52390 20046 52442
rect 20098 52390 50558 52442
rect 50610 52390 50662 52442
rect 50714 52390 50766 52442
rect 50818 52390 58576 52442
rect 1344 52356 58576 52390
rect 1344 51434 58576 51468
rect 1344 51382 4478 51434
rect 4530 51382 4582 51434
rect 4634 51382 4686 51434
rect 4738 51382 35198 51434
rect 35250 51382 35302 51434
rect 35354 51382 35406 51434
rect 35458 51382 58576 51434
rect 1344 51348 58576 51382
rect 1344 50426 58576 50460
rect 1344 50374 19838 50426
rect 19890 50374 19942 50426
rect 19994 50374 20046 50426
rect 20098 50374 50558 50426
rect 50610 50374 50662 50426
rect 50714 50374 50766 50426
rect 50818 50374 58576 50426
rect 1344 50340 58576 50374
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 32050 49086 32062 49138
rect 32114 49135 32126 49138
rect 33506 49135 33518 49138
rect 32114 49089 33518 49135
rect 32114 49086 32126 49089
rect 33506 49086 33518 49089
rect 33570 49086 33582 49138
rect 32062 49026 32114 49038
rect 32062 48962 32114 48974
rect 39230 48914 39282 48926
rect 39230 48850 39282 48862
rect 39566 48914 39618 48926
rect 39566 48850 39618 48862
rect 21422 48802 21474 48814
rect 21422 48738 21474 48750
rect 23662 48802 23714 48814
rect 23662 48738 23714 48750
rect 23998 48802 24050 48814
rect 23998 48738 24050 48750
rect 24334 48802 24386 48814
rect 24334 48738 24386 48750
rect 25230 48802 25282 48814
rect 25230 48738 25282 48750
rect 25790 48802 25842 48814
rect 25790 48738 25842 48750
rect 32510 48802 32562 48814
rect 32510 48738 32562 48750
rect 33070 48802 33122 48814
rect 33070 48738 33122 48750
rect 33518 48802 33570 48814
rect 33518 48738 33570 48750
rect 38782 48802 38834 48814
rect 38782 48738 38834 48750
rect 40686 48802 40738 48814
rect 40686 48738 40738 48750
rect 41358 48802 41410 48814
rect 41358 48738 41410 48750
rect 42590 48802 42642 48814
rect 42590 48738 42642 48750
rect 43150 48802 43202 48814
rect 43150 48738 43202 48750
rect 21870 48690 21922 48702
rect 21870 48626 21922 48638
rect 22318 48690 22370 48702
rect 22318 48626 22370 48638
rect 24670 48690 24722 48702
rect 24670 48626 24722 48638
rect 26462 48690 26514 48702
rect 26462 48626 26514 48638
rect 35534 48690 35586 48702
rect 35534 48626 35586 48638
rect 38334 48690 38386 48702
rect 41234 48638 41246 48690
rect 41298 48638 41310 48690
rect 38334 48626 38386 48638
rect 1344 48410 58576 48444
rect 1344 48358 19838 48410
rect 19890 48358 19942 48410
rect 19994 48358 20046 48410
rect 20098 48358 50558 48410
rect 50610 48358 50662 48410
rect 50714 48358 50766 48410
rect 50818 48358 58576 48410
rect 1344 48324 58576 48358
rect 26450 48190 26462 48242
rect 26514 48239 26526 48242
rect 27234 48239 27246 48242
rect 26514 48193 27246 48239
rect 26514 48190 26526 48193
rect 27234 48190 27246 48193
rect 27298 48239 27310 48242
rect 27682 48239 27694 48242
rect 27298 48193 27694 48239
rect 27298 48190 27310 48193
rect 27682 48190 27694 48193
rect 27746 48190 27758 48242
rect 23102 48130 23154 48142
rect 23102 48066 23154 48078
rect 26462 48130 26514 48142
rect 41470 48130 41522 48142
rect 35522 48078 35534 48130
rect 35586 48078 35598 48130
rect 26462 48066 26514 48078
rect 41470 48066 41522 48078
rect 19854 48018 19906 48030
rect 26014 48018 26066 48030
rect 22082 47966 22094 48018
rect 22146 47966 22158 48018
rect 19854 47954 19906 47966
rect 26014 47954 26066 47966
rect 28478 48018 28530 48030
rect 28478 47954 28530 47966
rect 19518 47906 19570 47918
rect 19518 47842 19570 47854
rect 27694 47906 27746 47918
rect 39006 47906 39058 47918
rect 36978 47854 36990 47906
rect 37042 47854 37054 47906
rect 27694 47842 27746 47854
rect 39006 47842 39058 47854
rect 19070 47794 19122 47806
rect 19070 47730 19122 47742
rect 23550 47794 23602 47806
rect 23550 47730 23602 47742
rect 23998 47794 24050 47806
rect 23998 47730 24050 47742
rect 26910 47794 26962 47806
rect 26910 47730 26962 47742
rect 27358 47794 27410 47806
rect 27358 47730 27410 47742
rect 32062 47794 32114 47806
rect 32062 47730 32114 47742
rect 32622 47794 32674 47806
rect 32622 47730 32674 47742
rect 40350 47794 40402 47806
rect 40350 47730 40402 47742
rect 41022 47794 41074 47806
rect 41022 47730 41074 47742
rect 41918 47794 41970 47806
rect 41918 47730 41970 47742
rect 42366 47794 42418 47806
rect 42366 47730 42418 47742
rect 42814 47794 42866 47806
rect 42814 47730 42866 47742
rect 43262 47794 43314 47806
rect 43262 47730 43314 47742
rect 43822 47794 43874 47806
rect 43822 47730 43874 47742
rect 44158 47794 44210 47806
rect 44158 47730 44210 47742
rect 45166 47794 45218 47806
rect 45166 47730 45218 47742
rect 50206 47794 50258 47806
rect 50206 47730 50258 47742
rect 50654 47794 50706 47806
rect 50654 47730 50706 47742
rect 52110 47794 52162 47806
rect 52110 47730 52162 47742
rect 52670 47794 52722 47806
rect 52670 47730 52722 47742
rect 53006 47794 53058 47806
rect 53006 47730 53058 47742
rect 53454 47794 53506 47806
rect 53454 47730 53506 47742
rect 31042 47630 31054 47682
rect 31106 47630 31118 47682
rect 41010 47630 41022 47682
rect 41074 47679 41086 47682
rect 41570 47679 41582 47682
rect 41074 47633 41582 47679
rect 41074 47630 41086 47633
rect 41570 47630 41582 47633
rect 41634 47679 41646 47682
rect 42354 47679 42366 47682
rect 41634 47633 42366 47679
rect 41634 47630 41646 47633
rect 42354 47630 42366 47633
rect 42418 47679 42430 47682
rect 43138 47679 43150 47682
rect 42418 47633 43150 47679
rect 42418 47630 42430 47633
rect 43138 47630 43150 47633
rect 43202 47630 43214 47682
rect 52098 47630 52110 47682
rect 52162 47679 52174 47682
rect 52994 47679 53006 47682
rect 52162 47633 53006 47679
rect 52162 47630 52174 47633
rect 52994 47630 53006 47633
rect 53058 47630 53070 47682
rect 27010 47518 27022 47570
rect 27074 47567 27086 47570
rect 27346 47567 27358 47570
rect 27074 47521 27358 47567
rect 27074 47518 27086 47521
rect 27346 47518 27358 47521
rect 27410 47518 27422 47570
rect 40786 47518 40798 47570
rect 40850 47567 40862 47570
rect 41346 47567 41358 47570
rect 40850 47521 41358 47567
rect 40850 47518 40862 47521
rect 41346 47518 41358 47521
rect 41410 47567 41422 47570
rect 41906 47567 41918 47570
rect 41410 47521 41918 47567
rect 41410 47518 41422 47521
rect 41906 47518 41918 47521
rect 41970 47567 41982 47570
rect 42802 47567 42814 47570
rect 41970 47521 42814 47567
rect 41970 47518 41982 47521
rect 42802 47518 42814 47521
rect 42866 47518 42878 47570
rect 1344 47402 58576 47436
rect 1344 47350 4478 47402
rect 4530 47350 4582 47402
rect 4634 47350 4686 47402
rect 4738 47350 35198 47402
rect 35250 47350 35302 47402
rect 35354 47350 35406 47402
rect 35458 47350 58576 47402
rect 1344 47316 58576 47350
rect 27234 47070 27246 47122
rect 27298 47119 27310 47122
rect 27794 47119 27806 47122
rect 27298 47073 27806 47119
rect 27298 47070 27310 47073
rect 27794 47070 27806 47073
rect 27858 47119 27870 47122
rect 28466 47119 28478 47122
rect 27858 47073 28478 47119
rect 27858 47070 27870 47073
rect 28466 47070 28478 47073
rect 28530 47070 28542 47122
rect 21646 47010 21698 47022
rect 27246 47010 27298 47022
rect 25890 46958 25902 47010
rect 25954 46958 25966 47010
rect 21646 46946 21698 46958
rect 27246 46946 27298 46958
rect 28142 47010 28194 47022
rect 28142 46946 28194 46958
rect 28590 47010 28642 47022
rect 28590 46946 28642 46958
rect 43150 47010 43202 47022
rect 43150 46946 43202 46958
rect 43598 47010 43650 47022
rect 43598 46946 43650 46958
rect 22430 46898 22482 46910
rect 22430 46834 22482 46846
rect 22878 46898 22930 46910
rect 22878 46834 22930 46846
rect 29374 46898 29426 46910
rect 29374 46834 29426 46846
rect 29822 46898 29874 46910
rect 32622 46898 32674 46910
rect 32162 46846 32174 46898
rect 32226 46846 32238 46898
rect 29822 46834 29874 46846
rect 32622 46834 32674 46846
rect 34078 46898 34130 46910
rect 34078 46834 34130 46846
rect 34862 46898 34914 46910
rect 34862 46834 34914 46846
rect 37550 46898 37602 46910
rect 37550 46834 37602 46846
rect 41246 46898 41298 46910
rect 52782 46898 52834 46910
rect 45490 46846 45502 46898
rect 45554 46846 45566 46898
rect 41246 46834 41298 46846
rect 52782 46834 52834 46846
rect 53678 46898 53730 46910
rect 53678 46834 53730 46846
rect 17838 46786 17890 46798
rect 17838 46722 17890 46734
rect 39118 46786 39170 46798
rect 39118 46722 39170 46734
rect 39454 46786 39506 46798
rect 39454 46722 39506 46734
rect 39790 46786 39842 46798
rect 39790 46722 39842 46734
rect 40686 46786 40738 46798
rect 40686 46722 40738 46734
rect 17390 46674 17442 46686
rect 17390 46610 17442 46622
rect 18510 46674 18562 46686
rect 18510 46610 18562 46622
rect 20526 46674 20578 46686
rect 20526 46610 20578 46622
rect 22094 46674 22146 46686
rect 22094 46610 22146 46622
rect 25118 46674 25170 46686
rect 25118 46610 25170 46622
rect 27694 46674 27746 46686
rect 27694 46610 27746 46622
rect 33182 46674 33234 46686
rect 33182 46610 33234 46622
rect 33854 46674 33906 46686
rect 33854 46610 33906 46622
rect 37102 46674 37154 46686
rect 37102 46610 37154 46622
rect 37998 46674 38050 46686
rect 37998 46610 38050 46622
rect 40126 46674 40178 46686
rect 40126 46610 40178 46622
rect 41918 46674 41970 46686
rect 41918 46610 41970 46622
rect 42702 46674 42754 46686
rect 42702 46610 42754 46622
rect 44046 46674 44098 46686
rect 44046 46610 44098 46622
rect 44942 46674 44994 46686
rect 44942 46610 44994 46622
rect 53230 46674 53282 46686
rect 53230 46610 53282 46622
rect 54126 46674 54178 46686
rect 54126 46610 54178 46622
rect 21634 46510 21646 46562
rect 21698 46559 21710 46562
rect 22082 46559 22094 46562
rect 21698 46513 22094 46559
rect 21698 46510 21710 46513
rect 22082 46510 22094 46513
rect 22146 46559 22158 46562
rect 22418 46559 22430 46562
rect 22146 46513 22430 46559
rect 22146 46510 22158 46513
rect 22418 46510 22430 46513
rect 22482 46510 22494 46562
rect 35634 46510 35646 46562
rect 35698 46510 35710 46562
rect 43138 46510 43150 46562
rect 43202 46559 43214 46562
rect 43922 46559 43934 46562
rect 43202 46513 43934 46559
rect 43202 46510 43214 46513
rect 43922 46510 43934 46513
rect 43986 46510 43998 46562
rect 50978 46510 50990 46562
rect 51042 46510 51054 46562
rect 53218 46510 53230 46562
rect 53282 46559 53294 46562
rect 53778 46559 53790 46562
rect 53282 46513 53790 46559
rect 53282 46510 53294 46513
rect 53778 46510 53790 46513
rect 53842 46510 53854 46562
rect 1344 46394 58576 46428
rect 1344 46342 19838 46394
rect 19890 46342 19942 46394
rect 19994 46342 20046 46394
rect 20098 46342 50558 46394
rect 50610 46342 50662 46394
rect 50714 46342 50766 46394
rect 50818 46342 58576 46394
rect 1344 46308 58576 46342
rect 32274 46174 32286 46226
rect 32338 46174 32350 46226
rect 41906 46174 41918 46226
rect 41970 46174 41982 46226
rect 22654 46114 22706 46126
rect 22654 46050 22706 46062
rect 23326 46114 23378 46126
rect 23326 46050 23378 46062
rect 24222 46114 24274 46126
rect 24222 46050 24274 46062
rect 25454 46114 25506 46126
rect 25454 46050 25506 46062
rect 26462 46114 26514 46126
rect 26462 46050 26514 46062
rect 27246 46114 27298 46126
rect 27246 46050 27298 46062
rect 30606 46114 30658 46126
rect 30606 46050 30658 46062
rect 35870 46114 35922 46126
rect 35870 46050 35922 46062
rect 39566 46114 39618 46126
rect 39566 46050 39618 46062
rect 46174 46114 46226 46126
rect 46174 46050 46226 46062
rect 25230 46002 25282 46014
rect 25230 45938 25282 45950
rect 28254 46002 28306 46014
rect 28254 45938 28306 45950
rect 31950 46002 32002 46014
rect 31950 45938 32002 45950
rect 33070 46002 33122 46014
rect 35198 46002 35250 46014
rect 34514 45950 34526 46002
rect 34578 45950 34590 46002
rect 33070 45938 33122 45950
rect 35198 45938 35250 45950
rect 40126 46002 40178 46014
rect 40126 45938 40178 45950
rect 41134 46002 41186 46014
rect 50878 46002 50930 46014
rect 44034 45950 44046 46002
rect 44098 45950 44110 46002
rect 41134 45938 41186 45950
rect 50878 45938 50930 45950
rect 51550 46002 51602 46014
rect 51550 45938 51602 45950
rect 53006 46002 53058 46014
rect 53006 45938 53058 45950
rect 53790 46002 53842 46014
rect 53790 45938 53842 45950
rect 54910 46002 54962 46014
rect 54910 45938 54962 45950
rect 55358 46002 55410 46014
rect 55358 45938 55410 45950
rect 17950 45890 18002 45902
rect 17950 45826 18002 45838
rect 18286 45890 18338 45902
rect 27806 45890 27858 45902
rect 20514 45838 20526 45890
rect 20578 45838 20590 45890
rect 18286 45826 18338 45838
rect 27806 45826 27858 45838
rect 31502 45890 31554 45902
rect 31502 45826 31554 45838
rect 33406 45890 33458 45902
rect 33406 45826 33458 45838
rect 33742 45890 33794 45902
rect 33742 45826 33794 45838
rect 34078 45890 34130 45902
rect 41582 45890 41634 45902
rect 37874 45838 37886 45890
rect 37938 45838 37950 45890
rect 39106 45838 39118 45890
rect 39170 45838 39182 45890
rect 41346 45838 41358 45890
rect 41410 45838 41422 45890
rect 34078 45826 34130 45838
rect 41582 45826 41634 45838
rect 41806 45890 41858 45902
rect 41806 45826 41858 45838
rect 42814 45890 42866 45902
rect 42814 45826 42866 45838
rect 43934 45890 43986 45902
rect 45266 45865 45278 45917
rect 45330 45865 45342 45917
rect 48750 45890 48802 45902
rect 43934 45826 43986 45838
rect 48750 45826 48802 45838
rect 49086 45890 49138 45902
rect 49086 45826 49138 45838
rect 49422 45890 49474 45902
rect 49422 45826 49474 45838
rect 49758 45890 49810 45902
rect 49758 45826 49810 45838
rect 50318 45890 50370 45902
rect 50318 45826 50370 45838
rect 53454 45890 53506 45902
rect 53454 45826 53506 45838
rect 54014 45890 54066 45902
rect 54014 45826 54066 45838
rect 17502 45778 17554 45790
rect 23774 45778 23826 45790
rect 21746 45726 21758 45778
rect 21810 45726 21822 45778
rect 17502 45714 17554 45726
rect 23774 45714 23826 45726
rect 24670 45778 24722 45790
rect 24670 45714 24722 45726
rect 36990 45778 37042 45790
rect 46622 45778 46674 45790
rect 37538 45726 37550 45778
rect 37602 45726 37614 45778
rect 36990 45714 37042 45726
rect 46622 45714 46674 45726
rect 47070 45778 47122 45790
rect 47070 45714 47122 45726
rect 48190 45778 48242 45790
rect 48190 45714 48242 45726
rect 52334 45778 52386 45790
rect 52334 45714 52386 45726
rect 53678 45778 53730 45790
rect 53678 45714 53730 45726
rect 23762 45614 23774 45666
rect 23826 45663 23838 45666
rect 24658 45663 24670 45666
rect 23826 45617 24670 45663
rect 23826 45614 23838 45617
rect 24658 45614 24670 45617
rect 24722 45614 24734 45666
rect 43810 45614 43822 45666
rect 43874 45614 43886 45666
rect 1344 45386 58576 45420
rect 1344 45334 4478 45386
rect 4530 45334 4582 45386
rect 4634 45334 4686 45386
rect 4738 45334 35198 45386
rect 35250 45334 35302 45386
rect 35354 45334 35406 45386
rect 35458 45334 58576 45386
rect 1344 45300 58576 45334
rect 38658 45166 38670 45218
rect 38722 45166 38734 45218
rect 48514 45166 48526 45218
rect 48578 45166 48590 45218
rect 35310 45106 35362 45118
rect 35310 45042 35362 45054
rect 34078 44994 34130 45006
rect 34078 44930 34130 44942
rect 37550 44994 37602 45006
rect 37550 44930 37602 44942
rect 17166 44882 17218 44894
rect 17166 44818 17218 44830
rect 17502 44882 17554 44894
rect 27358 44882 27410 44894
rect 18050 44830 18062 44882
rect 18114 44830 18126 44882
rect 24546 44830 24558 44882
rect 24610 44830 24622 44882
rect 17502 44818 17554 44830
rect 27358 44818 27410 44830
rect 32062 44882 32114 44894
rect 32062 44818 32114 44830
rect 32622 44882 32674 44894
rect 32622 44818 32674 44830
rect 34526 44882 34578 44894
rect 34526 44818 34578 44830
rect 36094 44882 36146 44894
rect 36094 44818 36146 44830
rect 37102 44882 37154 44894
rect 37102 44818 37154 44830
rect 37886 44882 37938 44894
rect 37886 44818 37938 44830
rect 38110 44882 38162 44894
rect 38110 44818 38162 44830
rect 38334 44882 38386 44894
rect 38334 44818 38386 44830
rect 39566 44882 39618 44894
rect 39566 44818 39618 44830
rect 43710 44882 43762 44894
rect 43710 44818 43762 44830
rect 44832 44882 44884 44894
rect 44832 44818 44884 44830
rect 45278 44882 45330 44894
rect 53006 44882 53058 44894
rect 46610 44830 46622 44882
rect 46674 44830 46686 44882
rect 50978 44830 50990 44882
rect 51042 44830 51054 44882
rect 45278 44818 45330 44830
rect 53006 44818 53058 44830
rect 54798 44882 54850 44894
rect 54798 44818 54850 44830
rect 21310 44770 21362 44782
rect 30494 44770 30546 44782
rect 21858 44718 21870 44770
rect 21922 44718 21934 44770
rect 28130 44718 28142 44770
rect 28194 44718 28206 44770
rect 21310 44706 21362 44718
rect 30494 44706 30546 44718
rect 30830 44770 30882 44782
rect 30830 44706 30882 44718
rect 31166 44770 31218 44782
rect 31166 44706 31218 44718
rect 39230 44770 39282 44782
rect 39230 44706 39282 44718
rect 39902 44770 39954 44782
rect 39902 44706 39954 44718
rect 40798 44770 40850 44782
rect 40798 44706 40850 44718
rect 41358 44770 41410 44782
rect 41358 44706 41410 44718
rect 43262 44770 43314 44782
rect 45054 44770 45106 44782
rect 43474 44718 43486 44770
rect 43538 44718 43550 44770
rect 43922 44718 43934 44770
rect 43986 44718 43998 44770
rect 43262 44706 43314 44718
rect 45054 44706 45106 44718
rect 50654 44770 50706 44782
rect 50654 44706 50706 44718
rect 51214 44770 51266 44782
rect 51214 44706 51266 44718
rect 51886 44770 51938 44782
rect 51886 44706 51938 44718
rect 52670 44770 52722 44782
rect 52670 44706 52722 44718
rect 53342 44770 53394 44782
rect 54114 44718 54126 44770
rect 54178 44718 54190 44770
rect 53342 44706 53394 44718
rect 20638 44658 20690 44670
rect 20290 44606 20302 44658
rect 20354 44606 20366 44658
rect 20638 44594 20690 44606
rect 24222 44658 24274 44670
rect 24222 44594 24274 44606
rect 25342 44658 25394 44670
rect 25342 44594 25394 44606
rect 26014 44658 26066 44670
rect 26014 44594 26066 44606
rect 28254 44658 28306 44670
rect 28254 44594 28306 44606
rect 31502 44658 31554 44670
rect 31502 44594 31554 44606
rect 33294 44658 33346 44670
rect 33294 44594 33346 44606
rect 40238 44658 40290 44670
rect 40238 44594 40290 44606
rect 42030 44658 42082 44670
rect 42030 44594 42082 44606
rect 43598 44658 43650 44670
rect 43598 44594 43650 44606
rect 44942 44658 44994 44670
rect 44942 44594 44994 44606
rect 51438 44658 51490 44670
rect 51438 44594 51490 44606
rect 53678 44658 53730 44670
rect 53678 44594 53730 44606
rect 55470 44658 55522 44670
rect 55470 44594 55522 44606
rect 1344 44378 58576 44412
rect 1344 44326 19838 44378
rect 19890 44326 19942 44378
rect 19994 44326 20046 44378
rect 20098 44326 50558 44378
rect 50610 44326 50662 44378
rect 50714 44326 50766 44378
rect 50818 44326 58576 44378
rect 1344 44292 58576 44326
rect 20290 44158 20302 44210
rect 20354 44207 20366 44210
rect 21186 44207 21198 44210
rect 20354 44161 21198 44207
rect 20354 44158 20366 44161
rect 21186 44158 21198 44161
rect 21250 44158 21262 44210
rect 24210 44158 24222 44210
rect 24274 44207 24286 44210
rect 24546 44207 24558 44210
rect 24274 44161 24558 44207
rect 24274 44158 24286 44161
rect 24546 44158 24558 44161
rect 24610 44158 24622 44210
rect 31266 44158 31278 44210
rect 31330 44158 31342 44210
rect 38098 44158 38110 44210
rect 38162 44207 38174 44210
rect 38994 44207 39006 44210
rect 38162 44161 39006 44207
rect 38162 44158 38174 44161
rect 38994 44158 39006 44161
rect 39058 44158 39070 44210
rect 40786 44158 40798 44210
rect 40850 44207 40862 44210
rect 41346 44207 41358 44210
rect 40850 44161 41358 44207
rect 40850 44158 40862 44161
rect 41346 44158 41358 44161
rect 41410 44158 41422 44210
rect 20302 44098 20354 44110
rect 20302 44034 20354 44046
rect 21198 44098 21250 44110
rect 21198 44034 21250 44046
rect 21646 44098 21698 44110
rect 21646 44034 21698 44046
rect 24222 44098 24274 44110
rect 24222 44034 24274 44046
rect 24670 44098 24722 44110
rect 24670 44034 24722 44046
rect 25678 44098 25730 44110
rect 25678 44034 25730 44046
rect 27246 44098 27298 44110
rect 27246 44034 27298 44046
rect 28702 44098 28754 44110
rect 34190 44098 34242 44110
rect 30482 44046 30494 44098
rect 30546 44046 30558 44098
rect 28702 44034 28754 44046
rect 34190 44034 34242 44046
rect 39006 44098 39058 44110
rect 39006 44034 39058 44046
rect 43486 44098 43538 44110
rect 45938 44046 45950 44098
rect 46002 44046 46014 44098
rect 48066 44046 48078 44098
rect 48130 44046 48142 44098
rect 55458 44046 55470 44098
rect 55522 44046 55534 44098
rect 43486 44034 43538 44046
rect 29038 43986 29090 43998
rect 29038 43922 29090 43934
rect 32174 43986 32226 43998
rect 32174 43922 32226 43934
rect 42142 43986 42194 43998
rect 42142 43922 42194 43934
rect 42590 43986 42642 43998
rect 42590 43922 42642 43934
rect 49646 43986 49698 43998
rect 53118 43986 53170 43998
rect 51874 43934 51886 43986
rect 51938 43934 51950 43986
rect 49646 43922 49698 43934
rect 53118 43922 53170 43934
rect 54686 43986 54738 43998
rect 54686 43922 54738 43934
rect 56702 43986 56754 43998
rect 56702 43922 56754 43934
rect 57150 43986 57202 43998
rect 57150 43922 57202 43934
rect 31726 43874 31778 43886
rect 31726 43810 31778 43822
rect 38558 43874 38610 43886
rect 38558 43810 38610 43822
rect 39454 43874 39506 43886
rect 39454 43810 39506 43822
rect 44046 43874 44098 43886
rect 44046 43810 44098 43822
rect 45166 43874 45218 43886
rect 45166 43810 45218 43822
rect 46958 43874 47010 43886
rect 46958 43810 47010 43822
rect 47294 43874 47346 43886
rect 50878 43874 50930 43886
rect 47394 43822 47406 43874
rect 47458 43822 47470 43874
rect 47618 43822 47630 43874
rect 47682 43822 47694 43874
rect 47294 43810 47346 43822
rect 50878 43810 50930 43822
rect 52894 43874 52946 43886
rect 52894 43810 52946 43822
rect 55022 43874 55074 43886
rect 55022 43810 55074 43822
rect 19854 43762 19906 43774
rect 19854 43698 19906 43710
rect 20750 43762 20802 43774
rect 20750 43698 20802 43710
rect 26126 43762 26178 43774
rect 26126 43698 26178 43710
rect 28030 43762 28082 43774
rect 28030 43698 28082 43710
rect 37326 43762 37378 43774
rect 37326 43698 37378 43710
rect 37774 43762 37826 43774
rect 37774 43698 37826 43710
rect 38110 43762 38162 43774
rect 38110 43698 38162 43710
rect 39902 43762 39954 43774
rect 39902 43698 39954 43710
rect 40350 43762 40402 43774
rect 40350 43698 40402 43710
rect 41022 43762 41074 43774
rect 41022 43698 41074 43710
rect 41470 43762 41522 43774
rect 41470 43698 41522 43710
rect 42814 43762 42866 43774
rect 42814 43698 42866 43710
rect 49534 43762 49586 43774
rect 49534 43698 49586 43710
rect 38658 43598 38670 43650
rect 38722 43647 38734 43650
rect 39106 43647 39118 43650
rect 38722 43601 39118 43647
rect 38722 43598 38734 43601
rect 39106 43598 39118 43601
rect 39170 43647 39182 43650
rect 39890 43647 39902 43650
rect 39170 43601 39902 43647
rect 39170 43598 39182 43601
rect 39890 43598 39902 43601
rect 39954 43647 39966 43650
rect 40338 43647 40350 43650
rect 39954 43601 40350 43647
rect 39954 43598 39966 43601
rect 40338 43598 40350 43601
rect 40402 43598 40414 43650
rect 20738 43486 20750 43538
rect 20802 43535 20814 43538
rect 21634 43535 21646 43538
rect 20802 43489 21646 43535
rect 20802 43486 20814 43489
rect 21634 43486 21646 43489
rect 21698 43486 21710 43538
rect 41682 43486 41694 43538
rect 41746 43486 41758 43538
rect 1344 43370 58576 43404
rect 1344 43318 4478 43370
rect 4530 43318 4582 43370
rect 4634 43318 4686 43370
rect 4738 43318 35198 43370
rect 35250 43318 35302 43370
rect 35354 43318 35406 43370
rect 35458 43318 58576 43370
rect 1344 43284 58576 43318
rect 47282 43150 47294 43202
rect 47346 43199 47358 43202
rect 48626 43199 48638 43202
rect 47346 43153 48638 43199
rect 47346 43150 47358 43153
rect 48626 43150 48638 43153
rect 48690 43150 48702 43202
rect 50642 43150 50654 43202
rect 50706 43199 50718 43202
rect 51538 43199 51550 43202
rect 50706 43153 51550 43199
rect 50706 43150 50718 43153
rect 51538 43150 51550 43153
rect 51602 43150 51614 43202
rect 33966 43090 34018 43102
rect 37090 43038 37102 43090
rect 37154 43087 37166 43090
rect 37538 43087 37550 43090
rect 37154 43041 37550 43087
rect 37154 43038 37166 43041
rect 37538 43038 37550 43041
rect 37602 43087 37614 43090
rect 38322 43087 38334 43090
rect 37602 43041 38334 43087
rect 37602 43038 37614 43041
rect 38322 43038 38334 43041
rect 38386 43038 38398 43090
rect 47730 43038 47742 43090
rect 47794 43087 47806 43090
rect 49074 43087 49086 43090
rect 47794 43041 49086 43087
rect 47794 43038 47806 43041
rect 49074 43038 49086 43041
rect 49138 43038 49150 43090
rect 33966 43026 34018 43038
rect 21646 42978 21698 42990
rect 21646 42914 21698 42926
rect 27246 42978 27298 42990
rect 27246 42914 27298 42926
rect 27694 42978 27746 42990
rect 27694 42914 27746 42926
rect 37550 42978 37602 42990
rect 37550 42914 37602 42926
rect 39790 42978 39842 42990
rect 39790 42914 39842 42926
rect 42478 42978 42530 42990
rect 42478 42914 42530 42926
rect 47294 42978 47346 42990
rect 47294 42914 47346 42926
rect 47742 42978 47794 42990
rect 47742 42914 47794 42926
rect 48638 42978 48690 42990
rect 48638 42914 48690 42926
rect 49086 42978 49138 42990
rect 49086 42914 49138 42926
rect 55134 42978 55186 42990
rect 55134 42914 55186 42926
rect 7534 42866 7586 42878
rect 23102 42866 23154 42878
rect 8082 42814 8094 42866
rect 8146 42814 8158 42866
rect 7534 42802 7586 42814
rect 23102 42802 23154 42814
rect 23438 42866 23490 42878
rect 23438 42802 23490 42814
rect 23774 42866 23826 42878
rect 23774 42802 23826 42814
rect 24670 42866 24722 42878
rect 24670 42802 24722 42814
rect 25230 42866 25282 42878
rect 25230 42802 25282 42814
rect 29038 42866 29090 42878
rect 29038 42802 29090 42814
rect 30270 42866 30322 42878
rect 30270 42802 30322 42814
rect 32958 42866 33010 42878
rect 32958 42802 33010 42814
rect 33294 42866 33346 42878
rect 33294 42802 33346 42814
rect 38670 42866 38722 42878
rect 38670 42802 38722 42814
rect 39454 42866 39506 42878
rect 39454 42802 39506 42814
rect 42590 42866 42642 42878
rect 42590 42802 42642 42814
rect 42702 42866 42754 42878
rect 42702 42802 42754 42814
rect 43598 42866 43650 42878
rect 46398 42866 46450 42878
rect 43922 42814 43934 42866
rect 43986 42814 43998 42866
rect 45378 42814 45390 42866
rect 45442 42814 45454 42866
rect 43598 42802 43650 42814
rect 46398 42802 46450 42814
rect 50206 42866 50258 42878
rect 50206 42802 50258 42814
rect 53230 42866 53282 42878
rect 53230 42802 53282 42814
rect 53454 42866 53506 42878
rect 54348 42866 54400 42878
rect 53778 42814 53790 42866
rect 53842 42814 53854 42866
rect 53454 42802 53506 42814
rect 54348 42802 54400 42814
rect 55358 42866 55410 42878
rect 55358 42802 55410 42814
rect 56142 42866 56194 42878
rect 56142 42802 56194 42814
rect 56478 42866 56530 42878
rect 56478 42802 56530 42814
rect 25902 42754 25954 42766
rect 25902 42690 25954 42702
rect 28142 42754 28194 42766
rect 28142 42690 28194 42702
rect 29374 42754 29426 42766
rect 29374 42690 29426 42702
rect 29598 42754 29650 42766
rect 29598 42690 29650 42702
rect 39230 42754 39282 42766
rect 41246 42754 41298 42766
rect 40450 42702 40462 42754
rect 40514 42702 40526 42754
rect 39230 42690 39282 42702
rect 41246 42690 41298 42702
rect 45166 42754 45218 42766
rect 45166 42690 45218 42702
rect 45614 42754 45666 42766
rect 55694 42754 55746 42766
rect 54226 42702 54238 42754
rect 54290 42702 54302 42754
rect 45614 42690 45666 42702
rect 55694 42690 55746 42702
rect 56926 42754 56978 42766
rect 56926 42690 56978 42702
rect 7198 42642 7250 42654
rect 7198 42578 7250 42590
rect 10222 42642 10274 42654
rect 10222 42578 10274 42590
rect 10670 42642 10722 42654
rect 10670 42578 10722 42590
rect 20414 42642 20466 42654
rect 20414 42578 20466 42590
rect 22094 42642 22146 42654
rect 22094 42578 22146 42590
rect 24110 42642 24162 42654
rect 24110 42578 24162 42590
rect 26798 42642 26850 42654
rect 26798 42578 26850 42590
rect 28590 42642 28642 42654
rect 28590 42578 28642 42590
rect 36430 42642 36482 42654
rect 36430 42578 36482 42590
rect 37102 42642 37154 42654
rect 37102 42578 37154 42590
rect 37998 42642 38050 42654
rect 37998 42578 38050 42590
rect 41918 42642 41970 42654
rect 41918 42578 41970 42590
rect 46846 42642 46898 42654
rect 46846 42578 46898 42590
rect 48190 42642 48242 42654
rect 48190 42578 48242 42590
rect 49758 42642 49810 42654
rect 49758 42578 49810 42590
rect 50654 42642 50706 42654
rect 50654 42578 50706 42590
rect 51102 42642 51154 42654
rect 51102 42578 51154 42590
rect 51550 42642 51602 42654
rect 51550 42578 51602 42590
rect 51998 42642 52050 42654
rect 51998 42578 52050 42590
rect 53342 42642 53394 42654
rect 53342 42578 53394 42590
rect 55806 42642 55858 42654
rect 55806 42578 55858 42590
rect 57374 42642 57426 42654
rect 57374 42578 57426 42590
rect 57822 42642 57874 42654
rect 57822 42578 57874 42590
rect 37090 42478 37102 42530
rect 37154 42527 37166 42530
rect 37986 42527 37998 42530
rect 37154 42481 37998 42527
rect 37154 42478 37166 42481
rect 37986 42478 37998 42481
rect 38050 42478 38062 42530
rect 44706 42478 44718 42530
rect 44770 42478 44782 42530
rect 55010 42478 55022 42530
rect 55074 42478 55086 42530
rect 56690 42478 56702 42530
rect 56754 42527 56766 42530
rect 57810 42527 57822 42530
rect 56754 42481 57822 42527
rect 56754 42478 56766 42481
rect 57810 42478 57822 42481
rect 57874 42478 57886 42530
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 35086 42082 35138 42094
rect 6850 42030 6862 42082
rect 6914 42030 6926 42082
rect 35086 42018 35138 42030
rect 44046 42082 44098 42094
rect 44046 42018 44098 42030
rect 48974 42082 49026 42094
rect 48974 42018 49026 42030
rect 50878 42082 50930 42094
rect 50878 42018 50930 42030
rect 52670 42082 52722 42094
rect 52670 42018 52722 42030
rect 56702 42082 56754 42094
rect 56702 42018 56754 42030
rect 9662 41970 9714 41982
rect 9662 41906 9714 41918
rect 9774 41970 9826 41982
rect 9774 41906 9826 41918
rect 19294 41970 19346 41982
rect 19294 41906 19346 41918
rect 19518 41970 19570 41982
rect 19518 41906 19570 41918
rect 21646 41970 21698 41982
rect 25342 41970 25394 41982
rect 22754 41918 22766 41970
rect 22818 41918 22830 41970
rect 21646 41906 21698 41918
rect 25342 41906 25394 41918
rect 27470 41970 27522 41982
rect 27470 41906 27522 41918
rect 27918 41970 27970 41982
rect 27918 41906 27970 41918
rect 30270 41970 30322 41982
rect 30270 41906 30322 41918
rect 30830 41970 30882 41982
rect 30830 41906 30882 41918
rect 34414 41970 34466 41982
rect 34414 41906 34466 41918
rect 36878 41970 36930 41982
rect 36878 41906 36930 41918
rect 39566 41970 39618 41982
rect 39566 41906 39618 41918
rect 41918 41970 41970 41982
rect 41918 41906 41970 41918
rect 42366 41970 42418 41982
rect 42366 41906 42418 41918
rect 43038 41970 43090 41982
rect 43038 41906 43090 41918
rect 43710 41970 43762 41982
rect 43710 41906 43762 41918
rect 45166 41970 45218 41982
rect 45166 41906 45218 41918
rect 45838 41970 45890 41982
rect 45838 41906 45890 41918
rect 52222 41970 52274 41982
rect 52222 41906 52274 41918
rect 53790 41970 53842 41982
rect 53790 41906 53842 41918
rect 54798 41970 54850 41982
rect 55682 41918 55694 41970
rect 55746 41918 55758 41970
rect 54798 41906 54850 41918
rect 4062 41858 4114 41870
rect 25566 41858 25618 41870
rect 4610 41806 4622 41858
rect 4674 41806 4686 41858
rect 10994 41806 11006 41858
rect 11058 41806 11070 41858
rect 4062 41794 4114 41806
rect 25566 41794 25618 41806
rect 26798 41858 26850 41870
rect 26798 41794 26850 41806
rect 33966 41858 34018 41870
rect 33966 41794 34018 41806
rect 36318 41858 36370 41870
rect 39902 41858 39954 41870
rect 43374 41858 43426 41870
rect 36418 41806 36430 41858
rect 36482 41806 36494 41858
rect 37762 41806 37774 41858
rect 37826 41806 37838 41858
rect 42130 41806 42142 41858
rect 42194 41806 42206 41858
rect 36318 41794 36370 41806
rect 39902 41794 39954 41806
rect 43374 41794 43426 41806
rect 44606 41858 44658 41870
rect 44606 41794 44658 41806
rect 46622 41858 46674 41870
rect 46622 41794 46674 41806
rect 52334 41858 52386 41870
rect 52334 41794 52386 41806
rect 56030 41858 56082 41870
rect 56030 41794 56082 41806
rect 1822 41746 1874 41758
rect 1822 41682 1874 41694
rect 3726 41746 3778 41758
rect 3726 41682 3778 41694
rect 24670 41746 24722 41758
rect 24670 41682 24722 41694
rect 28142 41746 28194 41758
rect 28142 41682 28194 41694
rect 28814 41746 28866 41758
rect 28814 41682 28866 41694
rect 30942 41746 30994 41758
rect 30942 41682 30994 41694
rect 31502 41746 31554 41758
rect 31502 41682 31554 41694
rect 33406 41746 33458 41758
rect 33406 41682 33458 41694
rect 40350 41746 40402 41758
rect 40350 41682 40402 41694
rect 41358 41746 41410 41758
rect 41358 41682 41410 41694
rect 49422 41746 49474 41758
rect 49422 41682 49474 41694
rect 49870 41746 49922 41758
rect 49870 41682 49922 41694
rect 50430 41746 50482 41758
rect 50430 41682 50482 41694
rect 51326 41746 51378 41758
rect 51326 41682 51378 41694
rect 57150 41746 57202 41758
rect 57150 41682 57202 41694
rect 57598 41746 57650 41758
rect 57598 41682 57650 41694
rect 37214 41634 37266 41646
rect 7186 41582 7198 41634
rect 7250 41582 7262 41634
rect 23874 41582 23886 41634
rect 23938 41582 23950 41634
rect 49410 41582 49422 41634
rect 49474 41631 49486 41634
rect 50418 41631 50430 41634
rect 49474 41585 50430 41631
rect 49474 41582 49486 41585
rect 50418 41582 50430 41585
rect 50482 41582 50494 41634
rect 55458 41582 55470 41634
rect 55522 41582 55534 41634
rect 37214 41570 37266 41582
rect 10882 41470 10894 41522
rect 10946 41470 10958 41522
rect 21522 41470 21534 41522
rect 21586 41470 21598 41522
rect 27010 41470 27022 41522
rect 27074 41470 27086 41522
rect 29810 41470 29822 41522
rect 29874 41470 29886 41522
rect 41458 41470 41470 41522
rect 41522 41470 41534 41522
rect 49858 41470 49870 41522
rect 49922 41519 49934 41522
rect 50866 41519 50878 41522
rect 49922 41473 50878 41519
rect 49922 41470 49934 41473
rect 50866 41470 50878 41473
rect 50930 41519 50942 41522
rect 51090 41519 51102 41522
rect 50930 41473 51102 41519
rect 50930 41470 50942 41473
rect 51090 41470 51102 41473
rect 51154 41519 51166 41522
rect 51314 41519 51326 41522
rect 51154 41473 51326 41519
rect 51154 41470 51166 41473
rect 51314 41470 51326 41473
rect 51378 41470 51390 41522
rect 1344 41354 58576 41388
rect 1344 41302 4478 41354
rect 4530 41302 4582 41354
rect 4634 41302 4686 41354
rect 4738 41302 35198 41354
rect 35250 41302 35302 41354
rect 35354 41302 35406 41354
rect 35458 41302 58576 41354
rect 1344 41268 58576 41302
rect 6178 41134 6190 41186
rect 6242 41134 6254 41186
rect 42690 41134 42702 41186
rect 42754 41183 42766 41186
rect 43362 41183 43374 41186
rect 42754 41137 43374 41183
rect 42754 41134 42766 41137
rect 43362 41134 43374 41137
rect 43426 41134 43438 41186
rect 55906 41134 55918 41186
rect 55970 41183 55982 41186
rect 56242 41183 56254 41186
rect 55970 41137 56254 41183
rect 55970 41134 55982 41137
rect 56242 41134 56254 41137
rect 56306 41134 56318 41186
rect 12114 41022 12126 41074
rect 12178 41022 12190 41074
rect 19854 40962 19906 40974
rect 19854 40898 19906 40910
rect 20302 40962 20354 40974
rect 20302 40898 20354 40910
rect 27134 40962 27186 40974
rect 27134 40898 27186 40910
rect 34638 40962 34690 40974
rect 34638 40898 34690 40910
rect 35534 40962 35586 40974
rect 35534 40898 35586 40910
rect 41918 40962 41970 40974
rect 41918 40898 41970 40910
rect 43150 40962 43202 40974
rect 43150 40898 43202 40910
rect 43598 40962 43650 40974
rect 43598 40898 43650 40910
rect 51214 40962 51266 40974
rect 51214 40898 51266 40910
rect 51998 40962 52050 40974
rect 51998 40898 52050 40910
rect 56254 40962 56306 40974
rect 56254 40898 56306 40910
rect 1822 40850 1874 40862
rect 8990 40850 9042 40862
rect 16606 40850 16658 40862
rect 2370 40798 2382 40850
rect 2434 40798 2446 40850
rect 6290 40798 6302 40850
rect 6354 40798 6366 40850
rect 9538 40798 9550 40850
rect 9602 40798 9614 40850
rect 1822 40786 1874 40798
rect 8990 40786 9042 40798
rect 16606 40786 16658 40798
rect 19294 40850 19346 40862
rect 19294 40786 19346 40798
rect 22766 40850 22818 40862
rect 22766 40786 22818 40798
rect 25454 40850 25506 40862
rect 25454 40786 25506 40798
rect 25790 40850 25842 40862
rect 36430 40850 36482 40862
rect 31826 40798 31838 40850
rect 31890 40798 31902 40850
rect 25790 40786 25842 40798
rect 36430 40786 36482 40798
rect 38446 40850 38498 40862
rect 52670 40850 52722 40862
rect 38882 40798 38894 40850
rect 38946 40798 38958 40850
rect 47954 40798 47966 40850
rect 48018 40798 48030 40850
rect 38446 40786 38498 40798
rect 52670 40786 52722 40798
rect 53006 40850 53058 40862
rect 53006 40786 53058 40798
rect 53342 40850 53394 40862
rect 53342 40786 53394 40798
rect 54798 40850 54850 40862
rect 54798 40786 54850 40798
rect 20750 40738 20802 40750
rect 20750 40674 20802 40686
rect 21534 40738 21586 40750
rect 21534 40674 21586 40686
rect 21870 40738 21922 40750
rect 21870 40674 21922 40686
rect 22318 40738 22370 40750
rect 22318 40674 22370 40686
rect 35982 40738 36034 40750
rect 35982 40674 36034 40686
rect 37886 40738 37938 40750
rect 37886 40674 37938 40686
rect 39678 40738 39730 40750
rect 39678 40674 39730 40686
rect 47070 40738 47122 40750
rect 47070 40674 47122 40686
rect 47742 40738 47794 40750
rect 47742 40674 47794 40686
rect 48302 40738 48354 40750
rect 48302 40674 48354 40686
rect 49534 40738 49586 40750
rect 49534 40674 49586 40686
rect 49982 40738 50034 40750
rect 49982 40674 50034 40686
rect 50542 40738 50594 40750
rect 50542 40674 50594 40686
rect 50654 40738 50706 40750
rect 50654 40674 50706 40686
rect 54238 40738 54290 40750
rect 54238 40674 54290 40686
rect 55470 40738 55522 40750
rect 55470 40674 55522 40686
rect 4958 40626 5010 40638
rect 4610 40574 4622 40626
rect 4674 40574 4686 40626
rect 4958 40562 5010 40574
rect 5742 40626 5794 40638
rect 5742 40562 5794 40574
rect 7982 40626 8034 40638
rect 7982 40562 8034 40574
rect 8654 40626 8706 40638
rect 8654 40562 8706 40574
rect 11678 40626 11730 40638
rect 11678 40562 11730 40574
rect 16158 40626 16210 40638
rect 16158 40562 16210 40574
rect 17278 40626 17330 40638
rect 17278 40562 17330 40574
rect 31278 40626 31330 40638
rect 35086 40626 35138 40638
rect 33170 40574 33182 40626
rect 33234 40574 33246 40626
rect 31278 40562 31330 40574
rect 35086 40562 35138 40574
rect 39566 40626 39618 40638
rect 39566 40562 39618 40574
rect 42702 40626 42754 40638
rect 42702 40562 42754 40574
rect 45390 40626 45442 40638
rect 45390 40562 45442 40574
rect 49198 40626 49250 40638
rect 49198 40562 49250 40574
rect 53678 40626 53730 40638
rect 53678 40562 53730 40574
rect 5618 40462 5630 40514
rect 5682 40462 5694 40514
rect 7858 40462 7870 40514
rect 7922 40462 7934 40514
rect 26562 40462 26574 40514
rect 26626 40462 26638 40514
rect 47282 40462 47294 40514
rect 47346 40462 47358 40514
rect 1344 40346 58576 40380
rect 1344 40294 19838 40346
rect 19890 40294 19942 40346
rect 19994 40294 20046 40346
rect 20098 40294 50558 40346
rect 50610 40294 50662 40346
rect 50714 40294 50766 40346
rect 50818 40294 58576 40346
rect 1344 40260 58576 40294
rect 30370 40126 30382 40178
rect 30434 40126 30446 40178
rect 48626 40126 48638 40178
rect 48690 40126 48702 40178
rect 1822 40066 1874 40078
rect 1822 40002 1874 40014
rect 4846 40066 4898 40078
rect 4846 40002 4898 40014
rect 5294 40066 5346 40078
rect 8878 40066 8930 40078
rect 21310 40066 21362 40078
rect 24670 40066 24722 40078
rect 8530 40014 8542 40066
rect 8594 40014 8606 40066
rect 12562 40014 12574 40066
rect 12626 40014 12638 40066
rect 23650 40014 23662 40066
rect 23714 40014 23726 40066
rect 5294 40002 5346 40014
rect 8878 40002 8930 40014
rect 21310 40002 21362 40014
rect 24670 40002 24722 40014
rect 35086 40066 35138 40078
rect 35086 40002 35138 40014
rect 41022 40066 41074 40078
rect 41022 40002 41074 40014
rect 44494 40066 44546 40078
rect 44494 40002 44546 40014
rect 44942 40066 44994 40078
rect 44942 40002 44994 40014
rect 45390 40066 45442 40078
rect 45390 40002 45442 40014
rect 46398 40066 46450 40078
rect 46398 40002 46450 40014
rect 53902 40066 53954 40078
rect 53902 40002 53954 40014
rect 18174 39954 18226 39966
rect 18174 39890 18226 39902
rect 20862 39954 20914 39966
rect 20862 39890 20914 39902
rect 22542 39954 22594 39966
rect 22542 39890 22594 39902
rect 26350 39954 26402 39966
rect 26350 39890 26402 39902
rect 33406 39954 33458 39966
rect 33406 39890 33458 39902
rect 33854 39954 33906 39966
rect 38446 39954 38498 39966
rect 36530 39902 36542 39954
rect 36594 39902 36606 39954
rect 37538 39902 37550 39954
rect 37602 39902 37614 39954
rect 33854 39890 33906 39902
rect 38446 39890 38498 39902
rect 45726 39954 45778 39966
rect 45726 39890 45778 39902
rect 49086 39954 49138 39966
rect 49086 39890 49138 39902
rect 49646 39954 49698 39966
rect 49646 39890 49698 39902
rect 50206 39954 50258 39966
rect 50206 39890 50258 39902
rect 51102 39954 51154 39966
rect 55694 39954 55746 39966
rect 54338 39902 54350 39954
rect 54402 39902 54414 39954
rect 51102 39890 51154 39902
rect 55694 39890 55746 39902
rect 2158 39842 2210 39854
rect 5742 39842 5794 39854
rect 9774 39842 9826 39854
rect 12910 39842 12962 39854
rect 17502 39842 17554 39854
rect 2706 39790 2718 39842
rect 2770 39790 2782 39842
rect 6290 39790 6302 39842
rect 6354 39790 6366 39842
rect 10322 39790 10334 39842
rect 10386 39790 10398 39842
rect 13458 39790 13470 39842
rect 13522 39790 13534 39842
rect 2158 39778 2210 39790
rect 5742 39778 5794 39790
rect 9774 39778 9826 39790
rect 12910 39778 12962 39790
rect 17502 39778 17554 39790
rect 20190 39842 20242 39854
rect 20190 39778 20242 39790
rect 21646 39842 21698 39854
rect 21646 39778 21698 39790
rect 30718 39842 30770 39854
rect 30718 39778 30770 39790
rect 32062 39842 32114 39854
rect 32062 39778 32114 39790
rect 35758 39842 35810 39854
rect 35758 39778 35810 39790
rect 37998 39842 38050 39854
rect 37998 39778 38050 39790
rect 38782 39842 38834 39854
rect 38782 39778 38834 39790
rect 41470 39842 41522 39854
rect 41470 39778 41522 39790
rect 41918 39842 41970 39854
rect 41918 39778 41970 39790
rect 48190 39842 48242 39854
rect 50430 39842 50482 39854
rect 49410 39790 49422 39842
rect 49474 39790 49486 39842
rect 48190 39778 48242 39790
rect 50430 39778 50482 39790
rect 50654 39848 50706 39860
rect 50654 39784 50706 39796
rect 50878 39842 50930 39854
rect 50878 39778 50930 39790
rect 51774 39842 51826 39854
rect 51774 39778 51826 39790
rect 52110 39842 52162 39854
rect 52110 39778 52162 39790
rect 52446 39842 52498 39854
rect 52446 39778 52498 39790
rect 52894 39842 52946 39854
rect 52894 39778 52946 39790
rect 53230 39842 53282 39854
rect 53230 39778 53282 39790
rect 53566 39842 53618 39854
rect 53566 39778 53618 39790
rect 55022 39842 55074 39854
rect 55022 39778 55074 39790
rect 57262 39842 57314 39854
rect 57262 39778 57314 39790
rect 16830 39730 16882 39742
rect 16830 39666 16882 39678
rect 25454 39730 25506 39742
rect 25454 39666 25506 39678
rect 31166 39730 31218 39742
rect 31166 39666 31218 39678
rect 31726 39730 31778 39742
rect 31726 39666 31778 39678
rect 34078 39730 34130 39742
rect 34078 39666 34130 39678
rect 39790 39730 39842 39742
rect 39790 39666 39842 39678
rect 40238 39730 40290 39742
rect 40238 39666 40290 39678
rect 44046 39730 44098 39742
rect 44046 39666 44098 39678
rect 13358 39618 13410 39630
rect 13358 39554 13410 39566
rect 32398 39618 32450 39630
rect 47518 39618 47570 39630
rect 41010 39566 41022 39618
rect 41074 39615 41086 39618
rect 41794 39615 41806 39618
rect 41074 39569 41806 39615
rect 41074 39566 41086 39569
rect 41794 39566 41806 39569
rect 41858 39566 41870 39618
rect 32398 39554 32450 39566
rect 47518 39554 47570 39566
rect 32946 39454 32958 39506
rect 33010 39454 33022 39506
rect 51202 39454 51214 39506
rect 51266 39454 51278 39506
rect 56802 39454 56814 39506
rect 56866 39454 56878 39506
rect 1344 39338 58576 39372
rect 1344 39286 4478 39338
rect 4530 39286 4582 39338
rect 4634 39286 4686 39338
rect 4738 39286 35198 39338
rect 35250 39286 35302 39338
rect 35354 39286 35406 39338
rect 35458 39286 58576 39338
rect 1344 39252 58576 39286
rect 6066 39118 6078 39170
rect 6130 39118 6142 39170
rect 52546 39118 52558 39170
rect 52610 39167 52622 39170
rect 53218 39167 53230 39170
rect 52610 39121 53230 39167
rect 52610 39118 52622 39121
rect 53218 39118 53230 39121
rect 53282 39118 53294 39170
rect 55794 39118 55806 39170
rect 55858 39167 55870 39170
rect 56802 39167 56814 39170
rect 55858 39121 56814 39167
rect 55858 39118 55870 39121
rect 56802 39118 56814 39121
rect 56866 39118 56878 39170
rect 53454 39058 53506 39070
rect 17154 39006 17166 39058
rect 17218 39006 17230 39058
rect 34626 39006 34638 39058
rect 34690 39055 34702 39058
rect 35074 39055 35086 39058
rect 34690 39009 35086 39055
rect 34690 39006 34702 39009
rect 35074 39006 35086 39009
rect 35138 39006 35150 39058
rect 55346 39006 55358 39058
rect 55410 39006 55422 39058
rect 53454 38994 53506 39006
rect 5630 38946 5682 38958
rect 5630 38882 5682 38894
rect 13470 38946 13522 38958
rect 13470 38882 13522 38894
rect 34862 38946 34914 38958
rect 34862 38882 34914 38894
rect 35310 38946 35362 38958
rect 35310 38882 35362 38894
rect 44270 38946 44322 38958
rect 44270 38882 44322 38894
rect 52782 38946 52834 38958
rect 52782 38882 52834 38894
rect 53230 38946 53282 38958
rect 53230 38882 53282 38894
rect 53566 38946 53618 38958
rect 56478 38946 56530 38958
rect 53778 38894 53790 38946
rect 53842 38943 53854 38946
rect 54114 38943 54126 38946
rect 53842 38897 54126 38943
rect 53842 38894 53854 38897
rect 54114 38894 54126 38897
rect 54178 38894 54190 38946
rect 53566 38882 53618 38894
rect 56478 38882 56530 38894
rect 56926 38946 56978 38958
rect 56926 38882 56978 38894
rect 1822 38834 1874 38846
rect 9662 38834 9714 38846
rect 19854 38834 19906 38846
rect 2370 38782 2382 38834
rect 2434 38782 2446 38834
rect 6178 38782 6190 38834
rect 6242 38782 6254 38834
rect 10210 38782 10222 38834
rect 10274 38782 10286 38834
rect 1822 38770 1874 38782
rect 9662 38770 9714 38782
rect 19854 38770 19906 38782
rect 23774 38834 23826 38846
rect 23774 38770 23826 38782
rect 24110 38834 24162 38846
rect 24110 38770 24162 38782
rect 24446 38834 24498 38846
rect 24446 38770 24498 38782
rect 24782 38834 24834 38846
rect 24782 38770 24834 38782
rect 25902 38834 25954 38846
rect 25902 38770 25954 38782
rect 36990 38834 37042 38846
rect 36990 38770 37042 38782
rect 37326 38834 37378 38846
rect 37326 38770 37378 38782
rect 37662 38834 37714 38846
rect 37662 38770 37714 38782
rect 38558 38834 38610 38846
rect 38558 38770 38610 38782
rect 39118 38834 39170 38846
rect 39118 38770 39170 38782
rect 42030 38834 42082 38846
rect 47630 38834 47682 38846
rect 45378 38782 45390 38834
rect 45442 38782 45454 38834
rect 42030 38770 42082 38782
rect 47630 38770 47682 38782
rect 48974 38834 49026 38846
rect 48974 38770 49026 38782
rect 49310 38834 49362 38846
rect 49310 38770 49362 38782
rect 49646 38834 49698 38846
rect 49646 38770 49698 38782
rect 54238 38834 54290 38846
rect 55570 38782 55582 38834
rect 55634 38782 55646 38834
rect 54238 38770 54290 38782
rect 4958 38722 5010 38734
rect 4958 38658 5010 38670
rect 5742 38722 5794 38734
rect 5742 38658 5794 38670
rect 12798 38722 12850 38734
rect 12798 38658 12850 38670
rect 13582 38722 13634 38734
rect 13582 38658 13634 38670
rect 20638 38722 20690 38734
rect 20638 38658 20690 38670
rect 25342 38722 25394 38734
rect 25342 38658 25394 38670
rect 26574 38722 26626 38734
rect 26574 38658 26626 38670
rect 27358 38722 27410 38734
rect 27358 38658 27410 38670
rect 30158 38722 30210 38734
rect 30158 38658 30210 38670
rect 30606 38722 30658 38734
rect 30606 38658 30658 38670
rect 36430 38722 36482 38734
rect 36430 38658 36482 38670
rect 39790 38722 39842 38734
rect 39790 38658 39842 38670
rect 40462 38722 40514 38734
rect 40462 38658 40514 38670
rect 40798 38722 40850 38734
rect 40798 38658 40850 38670
rect 41134 38722 41186 38734
rect 41134 38658 41186 38670
rect 42590 38722 42642 38734
rect 42590 38658 42642 38670
rect 43262 38722 43314 38734
rect 43262 38658 43314 38670
rect 44942 38722 44994 38734
rect 48190 38722 48242 38734
rect 46722 38670 46734 38722
rect 46786 38670 46798 38722
rect 44942 38658 44994 38670
rect 48190 38658 48242 38670
rect 48638 38722 48690 38734
rect 50766 38722 50818 38734
rect 50082 38670 50094 38722
rect 50146 38670 50158 38722
rect 48638 38658 48690 38670
rect 50766 38658 50818 38670
rect 51438 38722 51490 38734
rect 51438 38658 51490 38670
rect 53790 38722 53842 38734
rect 53790 38658 53842 38670
rect 54686 38722 54738 38734
rect 54686 38658 54738 38670
rect 56030 38722 56082 38734
rect 56030 38658 56082 38670
rect 6638 38610 6690 38622
rect 4610 38558 4622 38610
rect 4674 38558 4686 38610
rect 6638 38546 6690 38558
rect 8878 38610 8930 38622
rect 8878 38546 8930 38558
rect 9326 38610 9378 38622
rect 16830 38610 16882 38622
rect 12450 38558 12462 38610
rect 12514 38558 12526 38610
rect 9326 38546 9378 38558
rect 16830 38546 16882 38558
rect 19182 38610 19234 38622
rect 19182 38546 19234 38558
rect 33854 38610 33906 38622
rect 33854 38546 33906 38558
rect 37998 38610 38050 38622
rect 37998 38546 38050 38558
rect 41470 38610 41522 38622
rect 41470 38546 41522 38558
rect 1344 38330 58576 38364
rect 1344 38278 19838 38330
rect 19890 38278 19942 38330
rect 19994 38278 20046 38330
rect 20098 38278 50558 38330
rect 50610 38278 50662 38330
rect 50714 38278 50766 38330
rect 50818 38278 58576 38330
rect 1344 38244 58576 38278
rect 40226 38110 40238 38162
rect 40290 38110 40302 38162
rect 47618 38110 47630 38162
rect 47682 38159 47694 38162
rect 48178 38159 48190 38162
rect 47682 38113 48190 38159
rect 47682 38110 47694 38113
rect 48178 38110 48190 38113
rect 48242 38110 48254 38162
rect 1822 38050 1874 38062
rect 1822 37986 1874 37998
rect 2270 38050 2322 38062
rect 2270 37986 2322 37998
rect 5742 38050 5794 38062
rect 20862 38050 20914 38062
rect 13010 37998 13022 38050
rect 13074 37998 13086 38050
rect 5742 37986 5794 37998
rect 20862 37986 20914 37998
rect 23102 38050 23154 38062
rect 23102 37986 23154 37998
rect 23774 38050 23826 38062
rect 23774 37986 23826 37998
rect 33182 38050 33234 38062
rect 33182 37986 33234 37998
rect 47742 38050 47794 38062
rect 47742 37986 47794 37998
rect 48190 38050 48242 38062
rect 48190 37986 48242 37998
rect 49758 38050 49810 38062
rect 49758 37986 49810 37998
rect 55806 38050 55858 38062
rect 55806 37986 55858 37998
rect 18398 37938 18450 37950
rect 18398 37874 18450 37886
rect 25230 37938 25282 37950
rect 25230 37874 25282 37886
rect 27358 37938 27410 37950
rect 27358 37874 27410 37886
rect 31726 37938 31778 37950
rect 31726 37874 31778 37886
rect 32174 37938 32226 37950
rect 32174 37874 32226 37886
rect 38894 37938 38946 37950
rect 38894 37874 38946 37886
rect 42030 37938 42082 37950
rect 42030 37874 42082 37886
rect 43262 37938 43314 37950
rect 43262 37874 43314 37886
rect 44606 37938 44658 37950
rect 44606 37874 44658 37886
rect 46510 37938 46562 37950
rect 46510 37874 46562 37886
rect 49086 37938 49138 37950
rect 49086 37874 49138 37886
rect 53790 37938 53842 37950
rect 53790 37874 53842 37886
rect 55022 37938 55074 37950
rect 55022 37874 55074 37886
rect 3054 37826 3106 37838
rect 10222 37826 10274 37838
rect 13358 37826 13410 37838
rect 17614 37826 17666 37838
rect 2594 37774 2606 37826
rect 2658 37774 2670 37826
rect 3602 37774 3614 37826
rect 3666 37774 3678 37826
rect 10770 37774 10782 37826
rect 10834 37774 10846 37826
rect 13906 37774 13918 37826
rect 13970 37774 13982 37826
rect 3054 37762 3106 37774
rect 10222 37762 10274 37774
rect 13358 37762 13410 37774
rect 17614 37762 17666 37774
rect 25566 37826 25618 37838
rect 38222 37826 38274 37838
rect 31826 37774 31838 37826
rect 31890 37774 31902 37826
rect 33506 37774 33518 37826
rect 33570 37774 33582 37826
rect 25566 37762 25618 37774
rect 38222 37762 38274 37774
rect 41358 37826 41410 37838
rect 41358 37762 41410 37774
rect 41582 37826 41634 37838
rect 41582 37762 41634 37774
rect 41806 37826 41858 37838
rect 41806 37762 41858 37774
rect 42366 37826 42418 37838
rect 42366 37762 42418 37774
rect 42590 37826 42642 37838
rect 51550 37826 51602 37838
rect 46274 37774 46286 37826
rect 46338 37774 46350 37826
rect 42590 37762 42642 37774
rect 51550 37762 51602 37774
rect 52222 37826 52274 37838
rect 52222 37762 52274 37774
rect 52558 37826 52610 37838
rect 52558 37762 52610 37774
rect 52894 37826 52946 37838
rect 52894 37762 52946 37774
rect 53230 37826 53282 37838
rect 53230 37762 53282 37774
rect 54350 37826 54402 37838
rect 54350 37762 54402 37774
rect 9886 37714 9938 37726
rect 2594 37711 2606 37714
rect 2385 37665 2606 37711
rect 1922 37550 1934 37602
rect 1986 37599 1998 37602
rect 2385 37599 2431 37665
rect 2594 37662 2606 37665
rect 2658 37662 2670 37714
rect 9886 37650 9938 37662
rect 16830 37714 16882 37726
rect 16830 37650 16882 37662
rect 21422 37714 21474 37726
rect 21422 37650 21474 37662
rect 21870 37714 21922 37726
rect 21870 37650 21922 37662
rect 24222 37714 24274 37726
rect 24222 37650 24274 37662
rect 24670 37714 24722 37726
rect 24670 37650 24722 37662
rect 31054 37714 31106 37726
rect 31054 37650 31106 37662
rect 36654 37714 36706 37726
rect 36654 37650 36706 37662
rect 37102 37714 37154 37726
rect 37102 37650 37154 37662
rect 37662 37714 37714 37726
rect 37662 37650 37714 37662
rect 13806 37602 13858 37614
rect 1986 37553 2431 37599
rect 1986 37550 1998 37553
rect 6178 37550 6190 37602
rect 6242 37550 6254 37602
rect 20402 37550 20414 37602
rect 20466 37550 20478 37602
rect 41906 37550 41918 37602
rect 41970 37550 41982 37602
rect 13806 37538 13858 37550
rect 2706 37438 2718 37490
rect 2770 37438 2782 37490
rect 28354 37438 28366 37490
rect 28418 37438 28430 37490
rect 32610 37438 32622 37490
rect 32674 37438 32686 37490
rect 1344 37322 58576 37356
rect 1344 37270 4478 37322
rect 4530 37270 4582 37322
rect 4634 37270 4686 37322
rect 4738 37270 35198 37322
rect 35250 37270 35302 37322
rect 35354 37270 35406 37322
rect 35458 37270 58576 37322
rect 1344 37236 58576 37270
rect 52210 37102 52222 37154
rect 52274 37102 52286 37154
rect 43934 37042 43986 37054
rect 1922 36990 1934 37042
rect 1986 36990 1998 37042
rect 43934 36978 43986 36990
rect 50318 37042 50370 37054
rect 55122 36990 55134 37042
rect 55186 36990 55198 37042
rect 50318 36978 50370 36990
rect 6078 36930 6130 36942
rect 6078 36866 6130 36878
rect 9326 36930 9378 36942
rect 9326 36866 9378 36878
rect 16718 36930 16770 36942
rect 16718 36866 16770 36878
rect 20190 36930 20242 36942
rect 20190 36866 20242 36878
rect 23102 36930 23154 36942
rect 23102 36866 23154 36878
rect 24222 36930 24274 36942
rect 24222 36866 24274 36878
rect 32062 36930 32114 36942
rect 32062 36866 32114 36878
rect 36430 36930 36482 36942
rect 36430 36866 36482 36878
rect 43150 36930 43202 36942
rect 43150 36866 43202 36878
rect 49534 36930 49586 36942
rect 49534 36866 49586 36878
rect 53118 36930 53170 36942
rect 54114 36878 54126 36930
rect 54178 36878 54190 36930
rect 53118 36866 53170 36878
rect 5070 36818 5122 36830
rect 9662 36818 9714 36830
rect 19518 36818 19570 36830
rect 4498 36766 4510 36818
rect 4562 36766 4574 36818
rect 6178 36766 6190 36818
rect 6242 36766 6254 36818
rect 10210 36766 10222 36818
rect 10274 36766 10286 36818
rect 5070 36754 5122 36766
rect 9662 36754 9714 36766
rect 19518 36754 19570 36766
rect 21646 36818 21698 36830
rect 23886 36818 23938 36830
rect 38334 36818 38386 36830
rect 21858 36766 21870 36818
rect 21922 36766 21934 36818
rect 28354 36766 28366 36818
rect 28418 36766 28430 36818
rect 34066 36766 34078 36818
rect 34130 36766 34142 36818
rect 21646 36754 21698 36766
rect 23886 36754 23938 36766
rect 38334 36754 38386 36766
rect 39454 36818 39506 36830
rect 39454 36754 39506 36766
rect 42702 36818 42754 36830
rect 51774 36818 51826 36830
rect 57486 36818 57538 36830
rect 45938 36766 45950 36818
rect 46002 36766 46014 36818
rect 48178 36766 48190 36818
rect 48242 36766 48254 36818
rect 56018 36766 56030 36818
rect 56082 36766 56094 36818
rect 42702 36754 42754 36766
rect 51774 36754 51826 36766
rect 57486 36754 57538 36766
rect 5630 36706 5682 36718
rect 5630 36642 5682 36654
rect 22094 36706 22146 36718
rect 22094 36642 22146 36654
rect 26014 36706 26066 36718
rect 26014 36642 26066 36654
rect 37550 36706 37602 36718
rect 37550 36642 37602 36654
rect 37774 36706 37826 36718
rect 37774 36642 37826 36654
rect 38670 36706 38722 36718
rect 38670 36642 38722 36654
rect 39118 36706 39170 36718
rect 39118 36642 39170 36654
rect 39790 36706 39842 36718
rect 41246 36706 41298 36718
rect 40562 36654 40574 36706
rect 40626 36654 40638 36706
rect 39790 36642 39842 36654
rect 41246 36642 41298 36654
rect 41918 36706 41970 36718
rect 41918 36642 41970 36654
rect 44270 36706 44322 36718
rect 44270 36642 44322 36654
rect 45166 36706 45218 36718
rect 45166 36642 45218 36654
rect 47854 36706 47906 36718
rect 47854 36642 47906 36654
rect 49870 36706 49922 36718
rect 49870 36642 49922 36654
rect 50654 36706 50706 36718
rect 50654 36642 50706 36654
rect 51102 36706 51154 36718
rect 51102 36642 51154 36654
rect 51326 36706 51378 36718
rect 51326 36642 51378 36654
rect 52782 36706 52834 36718
rect 52782 36642 52834 36654
rect 54574 36706 54626 36718
rect 54574 36642 54626 36654
rect 57598 36706 57650 36718
rect 57598 36642 57650 36654
rect 5742 36594 5794 36606
rect 12798 36594 12850 36606
rect 2258 36542 2270 36594
rect 2322 36542 2334 36594
rect 12450 36542 12462 36594
rect 12514 36542 12526 36594
rect 5742 36530 5794 36542
rect 12798 36530 12850 36542
rect 13582 36594 13634 36606
rect 13582 36530 13634 36542
rect 16382 36594 16434 36606
rect 16382 36530 16434 36542
rect 18734 36594 18786 36606
rect 18734 36530 18786 36542
rect 20638 36594 20690 36606
rect 20638 36530 20690 36542
rect 21198 36594 21250 36606
rect 21198 36530 21250 36542
rect 23550 36594 23602 36606
rect 23550 36530 23602 36542
rect 27358 36594 27410 36606
rect 27358 36530 27410 36542
rect 29262 36594 29314 36606
rect 29262 36530 29314 36542
rect 31502 36594 31554 36606
rect 31502 36530 31554 36542
rect 37102 36594 37154 36606
rect 37102 36530 37154 36542
rect 40126 36594 40178 36606
rect 40126 36530 40178 36542
rect 43598 36594 43650 36606
rect 43598 36530 43650 36542
rect 49086 36594 49138 36606
rect 49086 36530 49138 36542
rect 13458 36430 13470 36482
rect 13522 36430 13534 36482
rect 27906 36430 27918 36482
rect 27970 36430 27982 36482
rect 42690 36430 42702 36482
rect 42754 36479 42766 36482
rect 43586 36479 43598 36482
rect 42754 36433 43598 36479
rect 42754 36430 42766 36433
rect 43586 36430 43598 36433
rect 43650 36430 43662 36482
rect 1344 36314 58576 36348
rect 1344 36262 19838 36314
rect 19890 36262 19942 36314
rect 19994 36262 20046 36314
rect 20098 36262 50558 36314
rect 50610 36262 50662 36314
rect 50714 36262 50766 36314
rect 50818 36262 58576 36314
rect 1344 36228 58576 36262
rect 17714 36094 17726 36146
rect 17778 36094 17790 36146
rect 19170 36094 19182 36146
rect 19234 36094 19246 36146
rect 20738 36094 20750 36146
rect 20802 36094 20814 36146
rect 36642 36094 36654 36146
rect 36706 36143 36718 36146
rect 37090 36143 37102 36146
rect 36706 36097 37102 36143
rect 36706 36094 36718 36097
rect 37090 36094 37102 36097
rect 37154 36094 37166 36146
rect 1822 36034 1874 36046
rect 1822 35970 1874 35982
rect 3054 36034 3106 36046
rect 36206 36034 36258 36046
rect 6178 35982 6190 36034
rect 6242 35982 6254 36034
rect 14130 35982 14142 36034
rect 14194 35982 14206 36034
rect 3054 35970 3106 35982
rect 36206 35970 36258 35982
rect 36654 36034 36706 36046
rect 36654 35970 36706 35982
rect 39678 36034 39730 36046
rect 39678 35970 39730 35982
rect 55694 36034 55746 36046
rect 55694 35970 55746 35982
rect 56702 36034 56754 36046
rect 56702 35970 56754 35982
rect 11006 35922 11058 35934
rect 11006 35858 11058 35870
rect 18174 35922 18226 35934
rect 18174 35858 18226 35870
rect 18622 35922 18674 35934
rect 18622 35858 18674 35870
rect 18846 35922 18898 35934
rect 18846 35858 18898 35870
rect 20190 35922 20242 35934
rect 20190 35858 20242 35870
rect 23886 35922 23938 35934
rect 23886 35858 23938 35870
rect 25902 35922 25954 35934
rect 25902 35858 25954 35870
rect 26462 35922 26514 35934
rect 26462 35858 26514 35870
rect 27806 35922 27858 35934
rect 27806 35858 27858 35870
rect 37102 35922 37154 35934
rect 37102 35858 37154 35870
rect 43038 35922 43090 35934
rect 43038 35858 43090 35870
rect 49422 35922 49474 35934
rect 49422 35858 49474 35870
rect 50206 35922 50258 35934
rect 54338 35870 54350 35922
rect 54402 35870 54414 35922
rect 50206 35858 50258 35870
rect 3390 35810 3442 35822
rect 6526 35810 6578 35822
rect 3938 35758 3950 35810
rect 4002 35758 4014 35810
rect 3390 35746 3442 35758
rect 6526 35746 6578 35758
rect 11342 35810 11394 35822
rect 19630 35810 19682 35822
rect 11890 35758 11902 35810
rect 11954 35758 11966 35810
rect 11342 35746 11394 35758
rect 19630 35746 19682 35758
rect 20302 35810 20354 35822
rect 20302 35746 20354 35758
rect 21086 35810 21138 35822
rect 21086 35746 21138 35758
rect 21870 35810 21922 35822
rect 21870 35746 21922 35758
rect 24558 35810 24610 35822
rect 24558 35746 24610 35758
rect 27022 35810 27074 35822
rect 27022 35746 27074 35758
rect 29822 35810 29874 35822
rect 29822 35746 29874 35758
rect 31838 35810 31890 35822
rect 37662 35810 37714 35822
rect 33506 35758 33518 35810
rect 33570 35758 33582 35810
rect 31838 35746 31890 35758
rect 37662 35746 37714 35758
rect 37886 35810 37938 35822
rect 37886 35746 37938 35758
rect 38334 35810 38386 35822
rect 38334 35746 38386 35758
rect 40350 35810 40402 35822
rect 40350 35746 40402 35758
rect 41246 35810 41298 35822
rect 41246 35746 41298 35758
rect 42814 35810 42866 35822
rect 42814 35746 42866 35758
rect 44046 35810 44098 35822
rect 50654 35810 50706 35822
rect 44370 35758 44382 35810
rect 44434 35758 44446 35810
rect 44046 35746 44098 35758
rect 50654 35746 50706 35758
rect 51102 35810 51154 35822
rect 52894 35810 52946 35822
rect 52098 35758 52110 35810
rect 52162 35758 52174 35810
rect 52322 35758 52334 35810
rect 52386 35807 52398 35810
rect 52386 35761 52607 35807
rect 52386 35758 52398 35761
rect 51102 35746 51154 35758
rect 16382 35698 16434 35710
rect 16382 35634 16434 35646
rect 16830 35698 16882 35710
rect 16830 35634 16882 35646
rect 17614 35698 17666 35710
rect 17614 35634 17666 35646
rect 21534 35698 21586 35710
rect 21534 35634 21586 35646
rect 26574 35698 26626 35710
rect 26574 35634 26626 35646
rect 33182 35698 33234 35710
rect 33182 35634 33234 35646
rect 34078 35698 34130 35710
rect 34078 35634 34130 35646
rect 41694 35698 41746 35710
rect 41694 35634 41746 35646
rect 44494 35698 44546 35710
rect 44494 35634 44546 35646
rect 44942 35698 44994 35710
rect 44942 35634 44994 35646
rect 45390 35698 45442 35710
rect 45390 35634 45442 35646
rect 48974 35698 49026 35710
rect 50082 35646 50094 35698
rect 50146 35646 50158 35698
rect 52561 35695 52607 35761
rect 52894 35746 52946 35758
rect 53230 35810 53282 35822
rect 53230 35746 53282 35758
rect 53566 35810 53618 35822
rect 53566 35746 53618 35758
rect 53902 35810 53954 35822
rect 53902 35746 53954 35758
rect 55022 35810 55074 35822
rect 55022 35746 55074 35758
rect 57150 35810 57202 35822
rect 57150 35746 57202 35758
rect 52882 35695 52894 35698
rect 52561 35649 52894 35695
rect 52882 35646 52894 35649
rect 52946 35646 52958 35698
rect 56802 35646 56814 35698
rect 56866 35646 56878 35698
rect 48974 35634 49026 35646
rect 31502 35586 31554 35598
rect 14466 35534 14478 35586
rect 14530 35534 14542 35586
rect 31502 35522 31554 35534
rect 40014 35586 40066 35598
rect 40014 35522 40066 35534
rect 40910 35586 40962 35598
rect 43362 35534 43374 35586
rect 43426 35534 43438 35586
rect 40910 35522 40962 35534
rect 25442 35422 25454 35474
rect 25506 35422 25518 35474
rect 33618 35422 33630 35474
rect 33682 35422 33694 35474
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 5618 35086 5630 35138
rect 5682 35086 5694 35138
rect 13458 35086 13470 35138
rect 13522 35086 13534 35138
rect 17266 35086 17278 35138
rect 17330 35086 17342 35138
rect 17714 35086 17726 35138
rect 17778 35135 17790 35138
rect 18162 35135 18174 35138
rect 17778 35089 18174 35135
rect 17778 35086 17790 35089
rect 18162 35086 18174 35089
rect 18226 35086 18238 35138
rect 18722 35086 18734 35138
rect 18786 35086 18798 35138
rect 27122 35086 27134 35138
rect 27186 35086 27198 35138
rect 35298 35086 35310 35138
rect 35362 35086 35374 35138
rect 50754 35086 50766 35138
rect 50818 35135 50830 35138
rect 51090 35135 51102 35138
rect 50818 35089 51102 35135
rect 50818 35086 50830 35089
rect 51090 35086 51102 35089
rect 51154 35086 51166 35138
rect 20750 35026 20802 35038
rect 20750 34962 20802 34974
rect 39678 35026 39730 35038
rect 39678 34962 39730 34974
rect 51886 35026 51938 35038
rect 56130 34974 56142 35026
rect 56194 35023 56206 35026
rect 56690 35023 56702 35026
rect 56194 34977 56702 35023
rect 56194 34974 56206 34977
rect 56690 34974 56702 34977
rect 56754 34974 56766 35026
rect 51886 34962 51938 34974
rect 18398 34914 18450 34926
rect 18398 34850 18450 34862
rect 19854 34914 19906 34926
rect 19854 34850 19906 34862
rect 21422 34914 21474 34926
rect 21422 34850 21474 34862
rect 30606 34914 30658 34926
rect 30606 34850 30658 34862
rect 44046 34914 44098 34926
rect 44046 34850 44098 34862
rect 44942 34914 44994 34926
rect 44942 34850 44994 34862
rect 49422 34914 49474 34926
rect 49422 34850 49474 34862
rect 50766 34914 50818 34926
rect 50766 34850 50818 34862
rect 51214 34914 51266 34926
rect 51214 34850 51266 34862
rect 54686 34914 54738 34926
rect 54686 34850 54738 34862
rect 56142 34914 56194 34926
rect 56142 34850 56194 34862
rect 20414 34802 20466 34814
rect 20414 34738 20466 34750
rect 21310 34802 21362 34814
rect 21310 34738 21362 34750
rect 21534 34802 21586 34814
rect 23326 34802 23378 34814
rect 22866 34750 22878 34802
rect 22930 34750 22942 34802
rect 21534 34738 21586 34750
rect 23326 34738 23378 34750
rect 24894 34802 24946 34814
rect 24894 34738 24946 34750
rect 25678 34802 25730 34814
rect 25678 34738 25730 34750
rect 26686 34802 26738 34814
rect 26686 34738 26738 34750
rect 27806 34802 27858 34814
rect 30942 34802 30994 34814
rect 28018 34750 28030 34802
rect 28082 34750 28094 34802
rect 29474 34750 29486 34802
rect 29538 34750 29550 34802
rect 27806 34738 27858 34750
rect 30942 34738 30994 34750
rect 33742 34802 33794 34814
rect 36990 34802 37042 34814
rect 35186 34750 35198 34802
rect 35250 34750 35262 34802
rect 33742 34738 33794 34750
rect 36990 34738 37042 34750
rect 37214 34802 37266 34814
rect 37214 34738 37266 34750
rect 38110 34802 38162 34814
rect 38110 34738 38162 34750
rect 38334 34802 38386 34814
rect 38334 34738 38386 34750
rect 38670 34802 38722 34814
rect 38670 34738 38722 34750
rect 38894 34802 38946 34814
rect 38894 34738 38946 34750
rect 49870 34802 49922 34814
rect 49870 34738 49922 34750
rect 52782 34802 52834 34814
rect 54910 34802 54962 34814
rect 52994 34750 53006 34802
rect 53058 34750 53070 34802
rect 52782 34738 52834 34750
rect 54910 34738 54962 34750
rect 16606 34690 16658 34702
rect 16606 34626 16658 34638
rect 17726 34690 17778 34702
rect 17726 34626 17778 34638
rect 18174 34690 18226 34702
rect 18174 34626 18226 34638
rect 19182 34690 19234 34702
rect 19182 34626 19234 34638
rect 19630 34690 19682 34702
rect 19630 34626 19682 34638
rect 21758 34690 21810 34702
rect 21758 34626 21810 34638
rect 21982 34690 22034 34702
rect 21982 34626 22034 34638
rect 22430 34690 22482 34702
rect 22430 34626 22482 34638
rect 23774 34690 23826 34702
rect 23774 34626 23826 34638
rect 25118 34690 25170 34702
rect 25118 34626 25170 34638
rect 26014 34690 26066 34702
rect 26014 34626 26066 34638
rect 26126 34690 26178 34702
rect 26126 34626 26178 34638
rect 28366 34690 28418 34702
rect 28366 34626 28418 34638
rect 33966 34690 34018 34702
rect 40014 34690 40066 34702
rect 34850 34638 34862 34690
rect 34914 34638 34926 34690
rect 33966 34626 34018 34638
rect 40014 34626 40066 34638
rect 42814 34690 42866 34702
rect 42814 34626 42866 34638
rect 51550 34690 51602 34702
rect 51550 34626 51602 34638
rect 55694 34690 55746 34702
rect 55694 34626 55746 34638
rect 56590 34690 56642 34702
rect 56590 34626 56642 34638
rect 5742 34578 5794 34590
rect 5742 34514 5794 34526
rect 13582 34578 13634 34590
rect 13582 34514 13634 34526
rect 16270 34578 16322 34590
rect 16270 34514 16322 34526
rect 17054 34578 17106 34590
rect 17054 34514 17106 34526
rect 22318 34578 22370 34590
rect 22318 34514 22370 34526
rect 22766 34578 22818 34590
rect 22766 34514 22818 34526
rect 24670 34578 24722 34590
rect 24670 34514 24722 34526
rect 25230 34578 25282 34590
rect 29374 34578 29426 34590
rect 25442 34526 25454 34578
rect 25506 34526 25518 34578
rect 25230 34514 25282 34526
rect 29374 34514 29426 34526
rect 31726 34578 31778 34590
rect 40686 34578 40738 34590
rect 38658 34526 38670 34578
rect 38722 34526 38734 34578
rect 31726 34514 31778 34526
rect 40686 34514 40738 34526
rect 41358 34578 41410 34590
rect 41358 34514 41410 34526
rect 41806 34578 41858 34590
rect 41806 34514 41858 34526
rect 42254 34578 42306 34590
rect 42254 34514 42306 34526
rect 43150 34578 43202 34590
rect 43150 34514 43202 34526
rect 45390 34578 45442 34590
rect 45390 34514 45442 34526
rect 45838 34578 45890 34590
rect 45838 34514 45890 34526
rect 46286 34578 46338 34590
rect 46286 34514 46338 34526
rect 50318 34578 50370 34590
rect 50318 34514 50370 34526
rect 54014 34578 54066 34590
rect 54014 34514 54066 34526
rect 55246 34578 55298 34590
rect 55246 34514 55298 34526
rect 27346 34414 27358 34466
rect 27410 34414 27422 34466
rect 37314 34414 37326 34466
rect 37378 34414 37390 34466
rect 37986 34414 37998 34466
rect 38050 34414 38062 34466
rect 1344 34298 58576 34332
rect 1344 34246 19838 34298
rect 19890 34246 19942 34298
rect 19994 34246 20046 34298
rect 20098 34246 50558 34298
rect 50610 34246 50662 34298
rect 50714 34246 50766 34298
rect 50818 34246 58576 34298
rect 1344 34212 58576 34246
rect 23426 34078 23438 34130
rect 23490 34078 23502 34130
rect 32274 34078 32286 34130
rect 32338 34078 32350 34130
rect 50194 34078 50206 34130
rect 50258 34127 50270 34130
rect 51090 34127 51102 34130
rect 50258 34081 51102 34127
rect 50258 34078 50270 34081
rect 51090 34078 51102 34081
rect 51154 34078 51166 34130
rect 3278 34018 3330 34030
rect 3278 33954 3330 33966
rect 3726 34018 3778 34030
rect 16830 34018 16882 34030
rect 4050 33966 4062 34018
rect 4114 33966 4126 34018
rect 3726 33954 3778 33966
rect 16830 33954 16882 33966
rect 19854 34018 19906 34030
rect 19854 33954 19906 33966
rect 20862 34018 20914 34030
rect 26462 34018 26514 34030
rect 25330 33966 25342 34018
rect 25394 33966 25406 34018
rect 20862 33954 20914 33966
rect 26462 33954 26514 33966
rect 27022 34018 27074 34030
rect 27022 33954 27074 33966
rect 28814 34018 28866 34030
rect 28814 33954 28866 33966
rect 30270 34018 30322 34030
rect 30270 33954 30322 33966
rect 36542 34018 36594 34030
rect 36542 33954 36594 33966
rect 37214 34018 37266 34030
rect 37214 33954 37266 33966
rect 40350 34018 40402 34030
rect 44718 34018 44770 34030
rect 42130 33966 42142 34018
rect 42194 33966 42206 34018
rect 40350 33954 40402 33966
rect 44718 33954 44770 33966
rect 47182 34018 47234 34030
rect 47182 33954 47234 33966
rect 48190 34018 48242 34030
rect 48190 33954 48242 33966
rect 50206 34018 50258 34030
rect 50206 33954 50258 33966
rect 50654 34018 50706 34030
rect 50654 33954 50706 33966
rect 51102 34018 51154 34030
rect 51102 33954 51154 33966
rect 51550 34018 51602 34030
rect 51550 33954 51602 33966
rect 51998 34018 52050 34030
rect 51998 33954 52050 33966
rect 55022 34018 55074 34030
rect 55022 33954 55074 33966
rect 11902 33906 11954 33918
rect 11902 33842 11954 33854
rect 16382 33906 16434 33918
rect 16382 33842 16434 33854
rect 18846 33906 18898 33918
rect 18846 33842 18898 33854
rect 20974 33906 21026 33918
rect 20974 33842 21026 33854
rect 21310 33906 21362 33918
rect 21310 33842 21362 33854
rect 21982 33906 22034 33918
rect 21982 33842 22034 33854
rect 22430 33906 22482 33918
rect 22430 33842 22482 33854
rect 22654 33906 22706 33918
rect 22654 33842 22706 33854
rect 23886 33906 23938 33918
rect 23886 33842 23938 33854
rect 24334 33906 24386 33918
rect 24334 33842 24386 33854
rect 25790 33906 25842 33918
rect 31278 33906 31330 33918
rect 27346 33854 27358 33906
rect 27410 33854 27422 33906
rect 25790 33842 25842 33854
rect 31278 33842 31330 33854
rect 31838 33906 31890 33918
rect 31838 33842 31890 33854
rect 33630 33906 33682 33918
rect 33630 33842 33682 33854
rect 34190 33906 34242 33918
rect 34190 33842 34242 33854
rect 35534 33906 35586 33918
rect 35534 33842 35586 33854
rect 36206 33906 36258 33918
rect 36206 33842 36258 33854
rect 36878 33906 36930 33918
rect 36878 33842 36930 33854
rect 42366 33906 42418 33918
rect 42366 33842 42418 33854
rect 53118 33906 53170 33918
rect 53118 33842 53170 33854
rect 54350 33906 54402 33918
rect 54350 33842 54402 33854
rect 6862 33794 6914 33806
rect 6290 33742 6302 33794
rect 6354 33742 6366 33794
rect 6862 33730 6914 33742
rect 18286 33794 18338 33806
rect 18286 33730 18338 33742
rect 20190 33794 20242 33806
rect 25118 33794 25170 33806
rect 22194 33742 22206 33794
rect 22258 33742 22270 33794
rect 24098 33742 24110 33794
rect 24162 33742 24174 33794
rect 20190 33730 20242 33742
rect 25118 33730 25170 33742
rect 26014 33794 26066 33806
rect 26014 33730 26066 33742
rect 26686 33794 26738 33806
rect 26686 33730 26738 33742
rect 27582 33794 27634 33806
rect 27582 33730 27634 33742
rect 30718 33794 30770 33806
rect 30718 33730 30770 33742
rect 35086 33794 35138 33806
rect 42254 33794 42306 33806
rect 35298 33742 35310 33794
rect 35362 33742 35374 33794
rect 35086 33730 35138 33742
rect 42254 33730 42306 33742
rect 44270 33794 44322 33806
rect 52670 33794 52722 33806
rect 45714 33742 45726 33794
rect 45778 33742 45790 33794
rect 52882 33742 52894 33794
rect 52946 33742 52958 33794
rect 44270 33730 44322 33742
rect 52670 33730 52722 33742
rect 12126 33682 12178 33694
rect 12126 33618 12178 33630
rect 17726 33682 17778 33694
rect 17726 33618 17778 33630
rect 18958 33682 19010 33694
rect 18958 33618 19010 33630
rect 23214 33682 23266 33694
rect 23214 33618 23266 33630
rect 25566 33682 25618 33694
rect 31166 33682 31218 33694
rect 27234 33630 27246 33682
rect 27298 33630 27310 33682
rect 25566 33618 25618 33630
rect 31166 33618 31218 33630
rect 34302 33682 34354 33694
rect 34302 33618 34354 33630
rect 37998 33682 38050 33694
rect 37998 33618 38050 33630
rect 41022 33682 41074 33694
rect 41022 33618 41074 33630
rect 43822 33682 43874 33694
rect 43822 33618 43874 33630
rect 45390 33682 45442 33694
rect 46734 33682 46786 33694
rect 46050 33630 46062 33682
rect 46114 33630 46126 33682
rect 45390 33618 45442 33630
rect 46734 33618 46786 33630
rect 53902 33682 53954 33694
rect 53902 33618 53954 33630
rect 55806 33682 55858 33694
rect 55806 33618 55858 33630
rect 12238 33570 12290 33582
rect 12238 33506 12290 33518
rect 17838 33570 17890 33582
rect 17838 33506 17890 33518
rect 21646 33570 21698 33582
rect 22194 33518 22206 33570
rect 22258 33518 22270 33570
rect 46050 33518 46062 33570
rect 46114 33518 46126 33570
rect 21646 33506 21698 33518
rect 33170 33406 33182 33458
rect 33234 33406 33246 33458
rect 34626 33406 34638 33458
rect 34690 33406 34702 33458
rect 46065 33455 46111 33518
rect 46834 33455 46846 33458
rect 46065 33409 46846 33455
rect 46834 33406 46846 33409
rect 46898 33406 46910 33458
rect 50642 33406 50654 33458
rect 50706 33455 50718 33458
rect 51538 33455 51550 33458
rect 50706 33409 51550 33455
rect 50706 33406 50718 33409
rect 51538 33406 51550 33409
rect 51602 33406 51614 33458
rect 52210 33406 52222 33458
rect 52274 33406 52286 33458
rect 1344 33290 58576 33324
rect 1344 33238 4478 33290
rect 4530 33238 4582 33290
rect 4634 33238 4686 33290
rect 4738 33238 35198 33290
rect 35250 33238 35302 33290
rect 35354 33238 35406 33290
rect 35458 33238 58576 33290
rect 1344 33204 58576 33238
rect 5730 33070 5742 33122
rect 5794 33070 5806 33122
rect 34414 33010 34466 33022
rect 12898 32958 12910 33010
rect 12962 32958 12974 33010
rect 34414 32946 34466 32958
rect 34750 33010 34802 33022
rect 34750 32946 34802 32958
rect 19742 32898 19794 32910
rect 19742 32834 19794 32846
rect 21758 32898 21810 32910
rect 21758 32834 21810 32846
rect 28590 32898 28642 32910
rect 28590 32834 28642 32846
rect 43486 32898 43538 32910
rect 43486 32834 43538 32846
rect 43934 32898 43986 32910
rect 43934 32834 43986 32846
rect 45054 32898 45106 32910
rect 45054 32834 45106 32846
rect 50654 32898 50706 32910
rect 50654 32834 50706 32846
rect 9774 32786 9826 32798
rect 9774 32722 9826 32734
rect 10110 32786 10162 32798
rect 15262 32786 15314 32798
rect 14018 32734 14030 32786
rect 14082 32734 14094 32786
rect 10110 32722 10162 32734
rect 15262 32722 15314 32734
rect 15710 32786 15762 32798
rect 15710 32722 15762 32734
rect 18398 32786 18450 32798
rect 18398 32722 18450 32734
rect 20190 32786 20242 32798
rect 20190 32722 20242 32734
rect 20638 32786 20690 32798
rect 20638 32722 20690 32734
rect 22094 32786 22146 32798
rect 24334 32786 24386 32798
rect 23538 32734 23550 32786
rect 23602 32734 23614 32786
rect 22094 32722 22146 32734
rect 24334 32722 24386 32734
rect 24446 32786 24498 32798
rect 24446 32722 24498 32734
rect 25342 32786 25394 32798
rect 30830 32786 30882 32798
rect 29810 32734 29822 32786
rect 29874 32734 29886 32786
rect 25342 32722 25394 32734
rect 30830 32722 30882 32734
rect 33518 32786 33570 32798
rect 38222 32786 38274 32798
rect 34066 32734 34078 32786
rect 34130 32734 34142 32786
rect 33518 32722 33570 32734
rect 38222 32722 38274 32734
rect 38334 32786 38386 32798
rect 38334 32722 38386 32734
rect 39790 32786 39842 32798
rect 39790 32722 39842 32734
rect 44270 32786 44322 32798
rect 44270 32722 44322 32734
rect 45390 32786 45442 32798
rect 45390 32722 45442 32734
rect 45726 32786 45778 32798
rect 46062 32786 46114 32798
rect 45826 32734 45838 32786
rect 45890 32734 45902 32786
rect 45726 32722 45778 32734
rect 46062 32722 46114 32734
rect 46846 32786 46898 32798
rect 46846 32722 46898 32734
rect 47070 32786 47122 32798
rect 47070 32722 47122 32734
rect 47294 32786 47346 32798
rect 53230 32786 53282 32798
rect 51874 32734 51886 32786
rect 51938 32734 51950 32786
rect 52882 32734 52894 32786
rect 52946 32734 52958 32786
rect 47294 32722 47346 32734
rect 53230 32722 53282 32734
rect 54014 32786 54066 32798
rect 54014 32722 54066 32734
rect 54126 32786 54178 32798
rect 56578 32734 56590 32786
rect 56642 32734 56654 32786
rect 54126 32722 54178 32734
rect 16382 32674 16434 32686
rect 16382 32610 16434 32622
rect 19070 32674 19122 32686
rect 19070 32610 19122 32622
rect 19518 32674 19570 32686
rect 19518 32610 19570 32622
rect 20302 32674 20354 32686
rect 20302 32610 20354 32622
rect 20414 32674 20466 32686
rect 25902 32674 25954 32686
rect 23650 32622 23662 32674
rect 23714 32622 23726 32674
rect 20414 32610 20466 32622
rect 25902 32610 25954 32622
rect 29486 32674 29538 32686
rect 29486 32610 29538 32622
rect 30046 32674 30098 32686
rect 30046 32610 30098 32622
rect 30494 32674 30546 32686
rect 30494 32610 30546 32622
rect 31502 32674 31554 32686
rect 31502 32610 31554 32622
rect 35086 32674 35138 32686
rect 35086 32610 35138 32622
rect 35534 32674 35586 32686
rect 35534 32610 35586 32622
rect 37102 32674 37154 32686
rect 37102 32610 37154 32622
rect 39118 32674 39170 32686
rect 39118 32610 39170 32622
rect 39454 32674 39506 32686
rect 39454 32610 39506 32622
rect 40126 32674 40178 32686
rect 40126 32610 40178 32622
rect 41022 32674 41074 32686
rect 41022 32610 41074 32622
rect 41582 32674 41634 32686
rect 41582 32610 41634 32622
rect 42254 32674 42306 32686
rect 42254 32610 42306 32622
rect 46622 32674 46674 32686
rect 46622 32610 46674 32622
rect 47966 32674 48018 32686
rect 47966 32610 48018 32622
rect 48414 32674 48466 32686
rect 48414 32610 48466 32622
rect 48974 32674 49026 32686
rect 48974 32610 49026 32622
rect 49758 32674 49810 32686
rect 49758 32610 49810 32622
rect 51326 32674 51378 32686
rect 51326 32610 51378 32622
rect 51774 32674 51826 32686
rect 51774 32610 51826 32622
rect 55022 32674 55074 32686
rect 55022 32610 55074 32622
rect 5630 32562 5682 32574
rect 5630 32498 5682 32510
rect 6078 32562 6130 32574
rect 6078 32498 6130 32510
rect 10894 32562 10946 32574
rect 10894 32498 10946 32510
rect 13470 32562 13522 32574
rect 13470 32498 13522 32510
rect 13582 32562 13634 32574
rect 13582 32498 13634 32510
rect 23214 32562 23266 32574
rect 23214 32498 23266 32510
rect 23886 32562 23938 32574
rect 23886 32498 23938 32510
rect 24110 32562 24162 32574
rect 24894 32562 24946 32574
rect 24658 32510 24670 32562
rect 24722 32510 24734 32562
rect 24110 32498 24162 32510
rect 24894 32498 24946 32510
rect 25118 32562 25170 32574
rect 25118 32498 25170 32510
rect 25566 32562 25618 32574
rect 25566 32498 25618 32510
rect 37550 32562 37602 32574
rect 37550 32498 37602 32510
rect 40462 32562 40514 32574
rect 40462 32498 40514 32510
rect 43038 32562 43090 32574
rect 47630 32562 47682 32574
rect 46834 32510 46846 32562
rect 46898 32510 46910 32562
rect 43038 32498 43090 32510
rect 47630 32498 47682 32510
rect 50206 32562 50258 32574
rect 50206 32498 50258 32510
rect 52894 32562 52946 32574
rect 52894 32498 52946 32510
rect 57038 32562 57090 32574
rect 57038 32498 57090 32510
rect 6178 32398 6190 32450
rect 6242 32398 6254 32450
rect 13906 32398 13918 32450
rect 13970 32398 13982 32450
rect 18610 32398 18622 32450
rect 18674 32398 18686 32450
rect 49298 32398 49310 32450
rect 49362 32398 49374 32450
rect 50866 32398 50878 32450
rect 50930 32398 50942 32450
rect 54674 32398 54686 32450
rect 54738 32398 54750 32450
rect 55570 32398 55582 32450
rect 55634 32398 55646 32450
rect 1344 32282 58576 32316
rect 1344 32230 19838 32282
rect 19890 32230 19942 32282
rect 19994 32230 20046 32282
rect 20098 32230 50558 32282
rect 50610 32230 50662 32282
rect 50714 32230 50766 32282
rect 50818 32230 58576 32282
rect 1344 32196 58576 32230
rect 41682 32062 41694 32114
rect 41746 32062 41758 32114
rect 8878 32002 8930 32014
rect 4162 31950 4174 32002
rect 4226 31950 4238 32002
rect 8878 31938 8930 31950
rect 9886 32002 9938 32014
rect 9886 31938 9938 31950
rect 14142 32002 14194 32014
rect 14142 31938 14194 31950
rect 16942 32002 16994 32014
rect 16942 31938 16994 31950
rect 18174 32002 18226 32014
rect 18174 31938 18226 31950
rect 26014 32002 26066 32014
rect 26014 31938 26066 31950
rect 30494 32002 30546 32014
rect 56814 32002 56866 32014
rect 44370 31950 44382 32002
rect 44434 31950 44446 32002
rect 52546 31950 52558 32002
rect 52610 31950 52622 32002
rect 30494 31938 30546 31950
rect 56814 31938 56866 31950
rect 57150 32002 57202 32014
rect 57150 31938 57202 31950
rect 3838 31890 3890 31902
rect 3838 31826 3890 31838
rect 10334 31890 10386 31902
rect 12238 31890 12290 31902
rect 10434 31838 10446 31890
rect 10498 31838 10510 31890
rect 10334 31826 10386 31838
rect 12238 31826 12290 31838
rect 13806 31890 13858 31902
rect 13806 31826 13858 31838
rect 14814 31890 14866 31902
rect 14814 31826 14866 31838
rect 15374 31890 15426 31902
rect 15374 31826 15426 31838
rect 21310 31890 21362 31902
rect 21310 31826 21362 31838
rect 24222 31890 24274 31902
rect 24222 31826 24274 31838
rect 29374 31890 29426 31902
rect 29374 31826 29426 31838
rect 34078 31890 34130 31902
rect 34078 31826 34130 31838
rect 37326 31890 37378 31902
rect 37326 31826 37378 31838
rect 40126 31890 40178 31902
rect 40126 31826 40178 31838
rect 42814 31890 42866 31902
rect 42814 31826 42866 31838
rect 45054 31890 45106 31902
rect 45054 31826 45106 31838
rect 45726 31890 45778 31902
rect 45726 31826 45778 31838
rect 47854 31890 47906 31902
rect 47854 31826 47906 31838
rect 48862 31890 48914 31902
rect 48862 31826 48914 31838
rect 49870 31890 49922 31902
rect 49870 31826 49922 31838
rect 50430 31890 50482 31902
rect 50430 31826 50482 31838
rect 51998 31890 52050 31902
rect 51998 31826 52050 31838
rect 52894 31890 52946 31902
rect 52894 31826 52946 31838
rect 53230 31890 53282 31902
rect 55694 31890 55746 31902
rect 54338 31838 54350 31890
rect 54402 31838 54414 31890
rect 53230 31826 53282 31838
rect 55694 31826 55746 31838
rect 58158 31890 58210 31902
rect 58158 31826 58210 31838
rect 3390 31778 3442 31790
rect 6974 31778 7026 31790
rect 16382 31778 16434 31790
rect 6402 31726 6414 31778
rect 6466 31726 6478 31778
rect 7410 31726 7422 31778
rect 7474 31726 7486 31778
rect 15138 31726 15150 31778
rect 15202 31726 15214 31778
rect 3390 31714 3442 31726
rect 6974 31714 7026 31726
rect 16382 31714 16434 31726
rect 17390 31778 17442 31790
rect 17390 31714 17442 31726
rect 20862 31778 20914 31790
rect 25230 31778 25282 31790
rect 21410 31726 21422 31778
rect 21474 31726 21486 31778
rect 24658 31726 24670 31778
rect 24722 31726 24734 31778
rect 20862 31714 20914 31726
rect 25230 31714 25282 31726
rect 29710 31778 29762 31790
rect 29710 31714 29762 31726
rect 33854 31778 33906 31790
rect 33854 31714 33906 31726
rect 34302 31778 34354 31790
rect 34302 31714 34354 31726
rect 36654 31778 36706 31790
rect 36654 31714 36706 31726
rect 37102 31778 37154 31790
rect 37102 31714 37154 31726
rect 39006 31778 39058 31790
rect 39006 31714 39058 31726
rect 41134 31778 41186 31790
rect 41134 31714 41186 31726
rect 41358 31778 41410 31790
rect 41358 31714 41410 31726
rect 43038 31778 43090 31790
rect 43038 31714 43090 31726
rect 45390 31778 45442 31790
rect 45390 31714 45442 31726
rect 46062 31778 46114 31790
rect 46062 31714 46114 31726
rect 46622 31778 46674 31790
rect 46622 31714 46674 31726
rect 47182 31778 47234 31790
rect 47182 31714 47234 31726
rect 49086 31778 49138 31790
rect 51326 31778 51378 31790
rect 50082 31726 50094 31778
rect 50146 31726 50158 31778
rect 49086 31714 49138 31726
rect 51326 31714 51378 31726
rect 51550 31778 51602 31790
rect 51550 31714 51602 31726
rect 51774 31778 51826 31790
rect 51774 31714 51826 31726
rect 52446 31778 52498 31790
rect 52446 31714 52498 31726
rect 53566 31778 53618 31790
rect 53566 31714 53618 31726
rect 53902 31778 53954 31790
rect 53902 31714 53954 31726
rect 55022 31778 55074 31790
rect 55022 31714 55074 31726
rect 56478 31778 56530 31790
rect 56478 31714 56530 31726
rect 57374 31778 57426 31790
rect 57374 31714 57426 31726
rect 8542 31666 8594 31678
rect 8542 31602 8594 31614
rect 14366 31666 14418 31678
rect 14366 31602 14418 31614
rect 20190 31666 20242 31678
rect 20190 31602 20242 31614
rect 22206 31666 22258 31678
rect 22206 31602 22258 31614
rect 34750 31666 34802 31678
rect 34750 31602 34802 31614
rect 35982 31666 36034 31678
rect 37774 31666 37826 31678
rect 52222 31666 52274 31678
rect 57710 31666 57762 31678
rect 37314 31614 37326 31666
rect 37378 31663 37390 31666
rect 37378 31617 37599 31663
rect 37378 31614 37390 31617
rect 35982 31602 36034 31614
rect 36990 31554 37042 31566
rect 12898 31502 12910 31554
rect 12962 31502 12974 31554
rect 28018 31502 28030 31554
rect 28082 31502 28094 31554
rect 32498 31502 32510 31554
rect 32562 31502 32574 31554
rect 37553 31551 37599 31617
rect 38546 31614 38558 31666
rect 38610 31614 38622 31666
rect 42914 31614 42926 31666
rect 42978 31614 42990 31666
rect 48738 31614 48750 31666
rect 48802 31614 48814 31666
rect 56802 31614 56814 31666
rect 56866 31614 56878 31666
rect 37774 31602 37826 31614
rect 52222 31602 52274 31614
rect 57710 31602 57762 31614
rect 37553 31505 37711 31551
rect 36990 31490 37042 31502
rect 37665 31442 37711 31505
rect 7298 31390 7310 31442
rect 7362 31390 7374 31442
rect 8978 31390 8990 31442
rect 9042 31390 9054 31442
rect 20402 31390 20414 31442
rect 20466 31390 20478 31442
rect 24546 31390 24558 31442
rect 24610 31390 24622 31442
rect 33954 31390 33966 31442
rect 34018 31390 34030 31442
rect 37650 31390 37662 31442
rect 37714 31439 37726 31442
rect 38098 31439 38110 31442
rect 37714 31393 38110 31439
rect 37714 31390 37726 31393
rect 38098 31390 38110 31393
rect 38162 31390 38174 31442
rect 49410 31390 49422 31442
rect 49474 31390 49486 31442
rect 1344 31274 58576 31308
rect 1344 31222 4478 31274
rect 4530 31222 4582 31274
rect 4634 31222 4686 31274
rect 4738 31222 35198 31274
rect 35250 31222 35302 31274
rect 35354 31222 35406 31274
rect 35458 31222 58576 31274
rect 1344 31188 58576 31222
rect 28466 31054 28478 31106
rect 28530 31054 28542 31106
rect 38782 30994 38834 31006
rect 8754 30942 8766 30994
rect 8818 30942 8830 30994
rect 26002 30942 26014 30994
rect 26066 30942 26078 30994
rect 38782 30930 38834 30942
rect 14926 30882 14978 30894
rect 14926 30818 14978 30830
rect 22878 30882 22930 30894
rect 32062 30882 32114 30894
rect 31154 30830 31166 30882
rect 31218 30830 31230 30882
rect 22878 30818 22930 30830
rect 32062 30818 32114 30830
rect 33742 30882 33794 30894
rect 33742 30818 33794 30830
rect 36990 30882 37042 30894
rect 36990 30818 37042 30830
rect 37662 30882 37714 30894
rect 37662 30818 37714 30830
rect 38222 30882 38274 30894
rect 38222 30818 38274 30830
rect 50206 30882 50258 30894
rect 50206 30818 50258 30830
rect 51214 30882 51266 30894
rect 51214 30818 51266 30830
rect 51550 30882 51602 30894
rect 51550 30818 51602 30830
rect 1822 30770 1874 30782
rect 5630 30770 5682 30782
rect 9886 30770 9938 30782
rect 2370 30718 2382 30770
rect 2434 30718 2446 30770
rect 6178 30718 6190 30770
rect 6242 30718 6254 30770
rect 1822 30706 1874 30718
rect 5630 30706 5682 30718
rect 9886 30706 9938 30718
rect 12462 30770 12514 30782
rect 12462 30706 12514 30718
rect 17950 30770 18002 30782
rect 17950 30706 18002 30718
rect 18622 30770 18674 30782
rect 18622 30706 18674 30718
rect 23214 30770 23266 30782
rect 27458 30718 27470 30770
rect 27522 30718 27534 30770
rect 28578 30718 28590 30770
rect 28642 30718 28654 30770
rect 30158 30764 30210 30776
rect 23214 30706 23266 30718
rect 30158 30700 30210 30712
rect 30828 30770 30880 30782
rect 30828 30706 30880 30718
rect 31502 30770 31554 30782
rect 31502 30706 31554 30718
rect 32622 30770 32674 30782
rect 32622 30706 32674 30718
rect 33070 30770 33122 30782
rect 33070 30706 33122 30718
rect 33406 30770 33458 30782
rect 33406 30706 33458 30718
rect 33854 30770 33906 30782
rect 33854 30706 33906 30718
rect 34974 30770 35026 30782
rect 34974 30706 35026 30718
rect 35198 30770 35250 30782
rect 35198 30706 35250 30718
rect 35422 30770 35474 30782
rect 35422 30706 35474 30718
rect 35646 30770 35698 30782
rect 35646 30706 35698 30718
rect 37326 30770 37378 30782
rect 37326 30706 37378 30718
rect 38446 30770 38498 30782
rect 42366 30770 42418 30782
rect 42130 30718 42142 30770
rect 42194 30718 42206 30770
rect 38446 30706 38498 30718
rect 42366 30706 42418 30718
rect 43374 30770 43426 30782
rect 50990 30770 51042 30782
rect 45938 30718 45950 30770
rect 46002 30718 46014 30770
rect 46498 30718 46510 30770
rect 46562 30718 46574 30770
rect 43374 30706 43426 30718
rect 50990 30706 51042 30718
rect 52670 30770 52722 30782
rect 56142 30770 56194 30782
rect 54002 30718 54014 30770
rect 54066 30718 54078 30770
rect 57586 30718 57598 30770
rect 57650 30718 57662 30770
rect 52670 30706 52722 30718
rect 56142 30706 56194 30718
rect 14030 30658 14082 30670
rect 14030 30594 14082 30606
rect 14702 30658 14754 30670
rect 14702 30594 14754 30606
rect 17614 30658 17666 30670
rect 17614 30594 17666 30606
rect 18286 30658 18338 30670
rect 19742 30658 19794 30670
rect 19058 30606 19070 30658
rect 19122 30606 19134 30658
rect 18286 30594 18338 30606
rect 19742 30594 19794 30606
rect 23998 30658 24050 30670
rect 23998 30594 24050 30606
rect 26686 30658 26738 30670
rect 26686 30594 26738 30606
rect 27022 30658 27074 30670
rect 27022 30594 27074 30606
rect 28142 30658 28194 30670
rect 28142 30594 28194 30606
rect 29150 30658 29202 30670
rect 29150 30594 29202 30606
rect 29934 30658 29986 30670
rect 29934 30594 29986 30606
rect 30606 30658 30658 30670
rect 30606 30594 30658 30606
rect 31278 30658 31330 30670
rect 31278 30594 31330 30606
rect 32846 30658 32898 30670
rect 32846 30594 32898 30606
rect 33630 30658 33682 30670
rect 33630 30594 33682 30606
rect 34638 30658 34690 30670
rect 34638 30594 34690 30606
rect 36430 30658 36482 30670
rect 36430 30594 36482 30606
rect 37886 30658 37938 30670
rect 37886 30594 37938 30606
rect 39118 30658 39170 30670
rect 39118 30594 39170 30606
rect 39454 30658 39506 30670
rect 39454 30594 39506 30606
rect 40798 30658 40850 30670
rect 40798 30594 40850 30606
rect 45166 30658 45218 30670
rect 49758 30658 49810 30670
rect 54462 30658 54514 30670
rect 48738 30606 48750 30658
rect 48802 30606 48814 30658
rect 51314 30606 51326 30658
rect 51378 30606 51390 30658
rect 45166 30594 45218 30606
rect 49758 30594 49810 30606
rect 54462 30594 54514 30606
rect 57262 30658 57314 30670
rect 57262 30594 57314 30606
rect 4958 30546 5010 30558
rect 4610 30494 4622 30546
rect 4674 30494 4686 30546
rect 4958 30482 5010 30494
rect 8318 30546 8370 30558
rect 8318 30482 8370 30494
rect 10558 30546 10610 30558
rect 10558 30482 10610 30494
rect 12126 30546 12178 30558
rect 12126 30482 12178 30494
rect 14366 30546 14418 30558
rect 14366 30482 14418 30494
rect 20414 30546 20466 30558
rect 27806 30546 27858 30558
rect 27234 30494 27246 30546
rect 27298 30494 27310 30546
rect 20414 30482 20466 30494
rect 27806 30482 27858 30494
rect 29486 30546 29538 30558
rect 29486 30482 29538 30494
rect 32958 30546 33010 30558
rect 32958 30482 33010 30494
rect 34302 30546 34354 30558
rect 34302 30482 34354 30494
rect 35086 30546 35138 30558
rect 35086 30482 35138 30494
rect 36094 30546 36146 30558
rect 36094 30482 36146 30494
rect 37550 30546 37602 30558
rect 37550 30482 37602 30494
rect 39790 30546 39842 30558
rect 39790 30482 39842 30494
rect 40462 30546 40514 30558
rect 40462 30482 40514 30494
rect 41134 30546 41186 30558
rect 41134 30482 41186 30494
rect 44382 30546 44434 30558
rect 44382 30482 44434 30494
rect 45502 30546 45554 30558
rect 45502 30482 45554 30494
rect 52110 30546 52162 30558
rect 55010 30494 55022 30546
rect 55074 30494 55086 30546
rect 52110 30482 52162 30494
rect 11666 30382 11678 30434
rect 11730 30382 11742 30434
rect 15026 30382 15038 30434
rect 15090 30382 15102 30434
rect 27010 30382 27022 30434
rect 27074 30382 27086 30434
rect 30034 30382 30046 30434
rect 30098 30382 30110 30434
rect 30706 30382 30718 30434
rect 30770 30382 30782 30434
rect 38098 30382 38110 30434
rect 38162 30382 38174 30434
rect 47618 30382 47630 30434
rect 47682 30382 47694 30434
rect 50642 30382 50654 30434
rect 50706 30382 50718 30434
rect 52994 30382 53006 30434
rect 53058 30382 53070 30434
rect 1344 30266 58576 30300
rect 1344 30214 19838 30266
rect 19890 30214 19942 30266
rect 19994 30214 20046 30266
rect 20098 30214 50558 30266
rect 50610 30214 50662 30266
rect 50714 30214 50766 30266
rect 50818 30214 58576 30266
rect 1344 30180 58576 30214
rect 11778 30046 11790 30098
rect 11842 30046 11854 30098
rect 12114 30046 12126 30098
rect 12178 30046 12190 30098
rect 21410 30046 21422 30098
rect 21474 30046 21486 30098
rect 27122 30046 27134 30098
rect 27186 30046 27198 30098
rect 39890 30046 39902 30098
rect 39954 30095 39966 30098
rect 40450 30095 40462 30098
rect 39954 30049 40462 30095
rect 39954 30046 39966 30049
rect 40450 30046 40462 30049
rect 40514 30046 40526 30098
rect 41682 30046 41694 30098
rect 41746 30095 41758 30098
rect 42130 30095 42142 30098
rect 41746 30049 42142 30095
rect 41746 30046 41758 30049
rect 42130 30046 42142 30049
rect 42194 30095 42206 30098
rect 42578 30095 42590 30098
rect 42194 30049 42590 30095
rect 42194 30046 42206 30049
rect 42578 30046 42590 30049
rect 42642 30046 42654 30098
rect 1822 29986 1874 29998
rect 1822 29922 1874 29934
rect 2830 29986 2882 29998
rect 2830 29922 2882 29934
rect 3726 29986 3778 29998
rect 7310 29986 7362 29998
rect 4050 29934 4062 29986
rect 4114 29934 4126 29986
rect 3726 29922 3778 29934
rect 7310 29922 7362 29934
rect 11678 29986 11730 29998
rect 11678 29922 11730 29934
rect 16270 29986 16322 29998
rect 16270 29922 16322 29934
rect 20414 29986 20466 29998
rect 20414 29922 20466 29934
rect 25678 29986 25730 29998
rect 25678 29922 25730 29934
rect 28478 29986 28530 29998
rect 28478 29922 28530 29934
rect 28814 29986 28866 29998
rect 28814 29922 28866 29934
rect 30494 29986 30546 29998
rect 30494 29922 30546 29934
rect 31838 29986 31890 29998
rect 31838 29922 31890 29934
rect 34750 29986 34802 29998
rect 34750 29922 34802 29934
rect 35086 29986 35138 29998
rect 35086 29922 35138 29934
rect 38222 29986 38274 29998
rect 38222 29922 38274 29934
rect 39230 29986 39282 29998
rect 39230 29922 39282 29934
rect 41246 29986 41298 29998
rect 41246 29922 41298 29934
rect 41694 29986 41746 29998
rect 41694 29922 41746 29934
rect 42590 29986 42642 29998
rect 42590 29922 42642 29934
rect 45726 29986 45778 29998
rect 45726 29922 45778 29934
rect 50318 29986 50370 29998
rect 50318 29922 50370 29934
rect 51662 29986 51714 29998
rect 51662 29922 51714 29934
rect 53902 29986 53954 29998
rect 53902 29922 53954 29934
rect 55694 29986 55746 29998
rect 55694 29922 55746 29934
rect 12574 29874 12626 29886
rect 12574 29810 12626 29822
rect 13134 29874 13186 29886
rect 13134 29810 13186 29822
rect 13246 29874 13298 29886
rect 13246 29810 13298 29822
rect 14926 29874 14978 29886
rect 14926 29810 14978 29822
rect 16158 29874 16210 29886
rect 16158 29810 16210 29822
rect 21870 29874 21922 29886
rect 21870 29810 21922 29822
rect 22318 29874 22370 29886
rect 22318 29810 22370 29822
rect 25902 29874 25954 29886
rect 25902 29810 25954 29822
rect 26574 29874 26626 29886
rect 26574 29810 26626 29822
rect 27022 29874 27074 29886
rect 27022 29810 27074 29822
rect 27134 29874 27186 29886
rect 27134 29810 27186 29822
rect 27470 29874 27522 29886
rect 27470 29810 27522 29822
rect 28142 29874 28194 29886
rect 28142 29810 28194 29822
rect 29150 29874 29202 29886
rect 38334 29874 38386 29886
rect 33506 29822 33518 29874
rect 33570 29822 33582 29874
rect 33842 29822 33854 29874
rect 33906 29822 33918 29874
rect 29150 29810 29202 29822
rect 38334 29810 38386 29822
rect 40910 29874 40962 29886
rect 40910 29810 40962 29822
rect 44718 29874 44770 29886
rect 44718 29810 44770 29822
rect 45390 29874 45442 29886
rect 45390 29810 45442 29822
rect 46286 29874 46338 29886
rect 46286 29810 46338 29822
rect 46846 29874 46898 29886
rect 46846 29810 46898 29822
rect 47518 29874 47570 29886
rect 47518 29810 47570 29822
rect 52894 29874 52946 29886
rect 52894 29810 52946 29822
rect 53230 29874 53282 29886
rect 53230 29810 53282 29822
rect 6862 29762 6914 29774
rect 3266 29710 3278 29762
rect 3330 29710 3342 29762
rect 6290 29710 6302 29762
rect 6354 29710 6366 29762
rect 6862 29698 6914 29710
rect 11118 29762 11170 29774
rect 11118 29698 11170 29710
rect 11230 29762 11282 29774
rect 11230 29698 11282 29710
rect 14366 29762 14418 29774
rect 14366 29698 14418 29710
rect 15934 29762 15986 29774
rect 15934 29698 15986 29710
rect 16382 29762 16434 29774
rect 16382 29698 16434 29710
rect 21086 29762 21138 29774
rect 23102 29762 23154 29774
rect 24446 29762 24498 29774
rect 22082 29710 22094 29762
rect 22146 29710 22158 29762
rect 22978 29710 22990 29762
rect 23042 29710 23054 29762
rect 24210 29710 24222 29762
rect 24274 29710 24286 29762
rect 21086 29698 21138 29710
rect 23102 29698 23154 29710
rect 24446 29698 24498 29710
rect 24670 29762 24722 29774
rect 34190 29762 34242 29774
rect 26114 29710 26126 29762
rect 26178 29710 26190 29762
rect 26338 29710 26350 29762
rect 26402 29710 26414 29762
rect 24670 29698 24722 29710
rect 34190 29698 34242 29710
rect 35422 29762 35474 29774
rect 35422 29698 35474 29710
rect 35646 29762 35698 29774
rect 35646 29698 35698 29710
rect 35870 29768 35922 29780
rect 35870 29704 35922 29716
rect 36094 29762 36146 29774
rect 36094 29698 36146 29710
rect 36654 29762 36706 29774
rect 36654 29698 36706 29710
rect 36878 29762 36930 29774
rect 36878 29698 36930 29710
rect 37102 29762 37154 29774
rect 37102 29698 37154 29710
rect 37326 29762 37378 29774
rect 37326 29698 37378 29710
rect 37886 29762 37938 29774
rect 37886 29698 37938 29710
rect 45054 29762 45106 29774
rect 45054 29698 45106 29710
rect 53566 29762 53618 29774
rect 53566 29698 53618 29710
rect 54462 29762 54514 29774
rect 54462 29698 54514 29710
rect 55022 29762 55074 29774
rect 55022 29698 55074 29710
rect 10446 29650 10498 29662
rect 10446 29586 10498 29598
rect 15038 29650 15090 29662
rect 15038 29586 15090 29598
rect 18062 29650 18114 29662
rect 33182 29650 33234 29662
rect 25666 29598 25678 29650
rect 25730 29647 25742 29650
rect 26674 29647 26686 29650
rect 25730 29601 26686 29647
rect 25730 29598 25742 29601
rect 26674 29598 26686 29601
rect 26738 29598 26750 29650
rect 18062 29586 18114 29598
rect 33182 29586 33234 29598
rect 33854 29650 33906 29662
rect 33854 29586 33906 29598
rect 36766 29650 36818 29662
rect 36766 29586 36818 29598
rect 39902 29650 39954 29662
rect 39902 29586 39954 29598
rect 40350 29650 40402 29662
rect 40350 29586 40402 29598
rect 42142 29650 42194 29662
rect 42142 29586 42194 29598
rect 44382 29650 44434 29662
rect 44382 29586 44434 29598
rect 48862 29650 48914 29662
rect 48862 29586 48914 29598
rect 49870 29650 49922 29662
rect 49870 29586 49922 29598
rect 50766 29650 50818 29662
rect 50766 29586 50818 29598
rect 51214 29650 51266 29662
rect 51214 29586 51266 29598
rect 52334 29650 52386 29662
rect 52334 29586 52386 29598
rect 18386 29486 18398 29538
rect 18450 29486 18462 29538
rect 49858 29486 49870 29538
rect 49922 29535 49934 29538
rect 50866 29535 50878 29538
rect 49922 29489 50878 29535
rect 49922 29486 49934 29489
rect 50866 29486 50878 29489
rect 50930 29535 50942 29538
rect 51314 29535 51326 29538
rect 50930 29489 51326 29535
rect 50930 29486 50942 29489
rect 51314 29486 51326 29489
rect 51378 29486 51390 29538
rect 3154 29374 3166 29426
rect 3218 29374 3230 29426
rect 13906 29374 13918 29426
rect 13970 29374 13982 29426
rect 24098 29374 24110 29426
rect 24162 29374 24174 29426
rect 25218 29374 25230 29426
rect 25282 29374 25294 29426
rect 34962 29374 34974 29426
rect 35026 29374 35038 29426
rect 36194 29374 36206 29426
rect 36258 29374 36270 29426
rect 50978 29374 50990 29426
rect 51042 29423 51054 29426
rect 51202 29423 51214 29426
rect 51042 29377 51214 29423
rect 51042 29374 51054 29377
rect 51202 29374 51214 29377
rect 51266 29374 51278 29426
rect 1344 29258 58576 29292
rect 1344 29206 4478 29258
rect 4530 29206 4582 29258
rect 4634 29206 4686 29258
rect 4738 29206 35198 29258
rect 35250 29206 35302 29258
rect 35354 29206 35406 29258
rect 35458 29206 58576 29258
rect 1344 29172 58576 29206
rect 5618 29038 5630 29090
rect 5682 29038 5694 29090
rect 15474 29038 15486 29090
rect 15538 29038 15550 29090
rect 18722 29038 18734 29090
rect 18786 29038 18798 29090
rect 21634 29038 21646 29090
rect 21698 29038 21710 29090
rect 26338 29038 26350 29090
rect 26402 29038 26414 29090
rect 41234 29038 41246 29090
rect 41298 29087 41310 29090
rect 43026 29087 43038 29090
rect 41298 29041 43038 29087
rect 41298 29038 41310 29041
rect 43026 29038 43038 29041
rect 43090 29038 43102 29090
rect 53778 29038 53790 29090
rect 53842 29038 53854 29090
rect 55570 29038 55582 29090
rect 55634 29038 55646 29090
rect 16942 28978 16994 28990
rect 16942 28914 16994 28926
rect 20638 28978 20690 28990
rect 20638 28914 20690 28926
rect 35086 28978 35138 28990
rect 38434 28926 38446 28978
rect 38498 28975 38510 28978
rect 38498 28929 38663 28975
rect 38498 28926 38510 28929
rect 35086 28914 35138 28926
rect 15150 28866 15202 28878
rect 15150 28802 15202 28814
rect 16606 28866 16658 28878
rect 16606 28802 16658 28814
rect 19854 28866 19906 28878
rect 19854 28802 19906 28814
rect 29150 28866 29202 28878
rect 29150 28802 29202 28814
rect 31166 28866 31218 28878
rect 31166 28802 31218 28814
rect 31614 28866 31666 28878
rect 31614 28802 31666 28814
rect 36430 28866 36482 28878
rect 36430 28802 36482 28814
rect 37102 28866 37154 28878
rect 37102 28802 37154 28814
rect 38446 28866 38498 28878
rect 38446 28802 38498 28814
rect 1822 28754 1874 28766
rect 14030 28754 14082 28766
rect 2370 28702 2382 28754
rect 2434 28702 2446 28754
rect 5730 28702 5742 28754
rect 5794 28702 5806 28754
rect 12338 28702 12350 28754
rect 12402 28702 12414 28754
rect 12898 28702 12910 28754
rect 12962 28702 12974 28754
rect 1822 28690 1874 28702
rect 14030 28690 14082 28702
rect 17390 28754 17442 28766
rect 20302 28754 20354 28766
rect 17714 28702 17726 28754
rect 17778 28702 17790 28754
rect 17390 28690 17442 28702
rect 20302 28690 20354 28702
rect 21310 28754 21362 28766
rect 21310 28690 21362 28702
rect 21758 28754 21810 28766
rect 24670 28754 24722 28766
rect 24434 28702 24446 28754
rect 24498 28702 24510 28754
rect 21758 28690 21810 28702
rect 24670 28690 24722 28702
rect 24894 28754 24946 28766
rect 24894 28690 24946 28702
rect 26462 28754 26514 28766
rect 26462 28690 26514 28702
rect 26686 28754 26738 28766
rect 26686 28690 26738 28702
rect 26910 28754 26962 28766
rect 26910 28690 26962 28702
rect 27134 28754 27186 28766
rect 27134 28690 27186 28702
rect 29486 28754 29538 28766
rect 29486 28690 29538 28702
rect 29934 28754 29986 28766
rect 33742 28754 33794 28766
rect 33282 28702 33294 28754
rect 33346 28702 33358 28754
rect 29934 28690 29986 28702
rect 33742 28690 33794 28702
rect 34302 28754 34354 28766
rect 34302 28690 34354 28702
rect 34526 28754 34578 28766
rect 34526 28690 34578 28702
rect 34750 28754 34802 28766
rect 34750 28690 34802 28702
rect 34974 28754 35026 28766
rect 34974 28690 35026 28702
rect 35310 28754 35362 28766
rect 36878 28754 36930 28766
rect 35634 28702 35646 28754
rect 35698 28702 35710 28754
rect 37202 28702 37214 28754
rect 37266 28702 37278 28754
rect 35310 28690 35362 28702
rect 36878 28690 36930 28702
rect 4958 28642 5010 28654
rect 4958 28578 5010 28590
rect 6078 28642 6130 28654
rect 6078 28578 6130 28590
rect 6190 28642 6242 28654
rect 6190 28578 6242 28590
rect 12238 28642 12290 28654
rect 12238 28578 12290 28590
rect 13470 28642 13522 28654
rect 13470 28578 13522 28590
rect 14478 28642 14530 28654
rect 14478 28578 14530 28590
rect 15038 28642 15090 28654
rect 15038 28578 15090 28590
rect 15934 28642 15986 28654
rect 15934 28578 15986 28590
rect 16494 28642 16546 28654
rect 16494 28578 16546 28590
rect 17950 28642 18002 28654
rect 17950 28578 18002 28590
rect 19182 28642 19234 28654
rect 19182 28578 19234 28590
rect 19630 28642 19682 28654
rect 19630 28578 19682 28590
rect 21534 28642 21586 28654
rect 21534 28578 21586 28590
rect 25118 28642 25170 28654
rect 25118 28578 25170 28590
rect 25790 28642 25842 28654
rect 25790 28578 25842 28590
rect 26014 28642 26066 28654
rect 26014 28578 26066 28590
rect 27358 28642 27410 28654
rect 27358 28578 27410 28590
rect 28030 28642 28082 28654
rect 28030 28578 28082 28590
rect 28254 28642 28306 28654
rect 28254 28578 28306 28590
rect 30718 28642 30770 28654
rect 30718 28578 30770 28590
rect 32398 28642 32450 28654
rect 32398 28578 32450 28590
rect 35534 28642 35586 28654
rect 37438 28642 37490 28654
rect 35970 28590 35982 28642
rect 36034 28590 36046 28642
rect 35534 28578 35586 28590
rect 37438 28578 37490 28590
rect 4510 28530 4562 28542
rect 4510 28466 4562 28478
rect 13582 28530 13634 28542
rect 25566 28530 25618 28542
rect 24322 28478 24334 28530
rect 24386 28478 24398 28530
rect 13582 28466 13634 28478
rect 25566 28466 25618 28478
rect 27806 28530 27858 28542
rect 27806 28466 27858 28478
rect 30382 28530 30434 28542
rect 30382 28466 30434 28478
rect 32062 28530 32114 28542
rect 32062 28466 32114 28478
rect 32734 28530 32786 28542
rect 32734 28466 32786 28478
rect 33070 28530 33122 28542
rect 33070 28466 33122 28478
rect 37998 28530 38050 28542
rect 38617 28527 38663 28929
rect 45938 28926 45950 28978
rect 46002 28975 46014 28978
rect 46498 28975 46510 28978
rect 46002 28929 46510 28975
rect 46002 28926 46014 28929
rect 46498 28926 46510 28929
rect 46562 28975 46574 28978
rect 46834 28975 46846 28978
rect 46562 28929 46846 28975
rect 46562 28926 46574 28929
rect 46834 28926 46846 28929
rect 46898 28926 46910 28978
rect 42142 28866 42194 28878
rect 42142 28802 42194 28814
rect 43038 28866 43090 28878
rect 43038 28802 43090 28814
rect 45950 28866 46002 28878
rect 45950 28802 46002 28814
rect 46398 28866 46450 28878
rect 46398 28802 46450 28814
rect 50542 28866 50594 28878
rect 50542 28802 50594 28814
rect 52782 28866 52834 28878
rect 52782 28802 52834 28814
rect 53230 28866 53282 28878
rect 54114 28814 54126 28866
rect 54178 28814 54190 28866
rect 53230 28802 53282 28814
rect 39342 28754 39394 28766
rect 39342 28690 39394 28702
rect 40238 28754 40290 28766
rect 40238 28690 40290 28702
rect 41246 28754 41298 28766
rect 41246 28690 41298 28702
rect 47070 28754 47122 28766
rect 47070 28690 47122 28702
rect 47630 28754 47682 28766
rect 47630 28690 47682 28702
rect 48078 28754 48130 28766
rect 48290 28702 48302 28754
rect 48354 28702 48366 28754
rect 55682 28702 55694 28754
rect 55746 28702 55758 28754
rect 48078 28690 48130 28702
rect 42590 28642 42642 28654
rect 54562 28590 54574 28642
rect 54626 28590 54638 28642
rect 42590 28578 42642 28590
rect 38894 28530 38946 28542
rect 38617 28481 38831 28527
rect 37998 28466 38050 28478
rect 12786 28366 12798 28418
rect 12850 28366 12862 28418
rect 25330 28366 25342 28418
rect 25394 28366 25406 28418
rect 27570 28366 27582 28418
rect 27634 28366 27646 28418
rect 38785 28415 38831 28481
rect 38894 28466 38946 28478
rect 41694 28530 41746 28542
rect 41694 28466 41746 28478
rect 45054 28530 45106 28542
rect 45054 28466 45106 28478
rect 45502 28530 45554 28542
rect 45502 28466 45554 28478
rect 48974 28530 49026 28542
rect 48974 28466 49026 28478
rect 50094 28530 50146 28542
rect 50094 28466 50146 28478
rect 50990 28530 51042 28542
rect 50990 28466 51042 28478
rect 51662 28530 51714 28542
rect 51662 28466 51714 28478
rect 52110 28530 52162 28542
rect 52110 28466 52162 28478
rect 56702 28530 56754 28542
rect 56702 28466 56754 28478
rect 39218 28415 39230 28418
rect 38785 28369 39230 28415
rect 39218 28366 39230 28369
rect 39282 28366 39294 28418
rect 39890 28366 39902 28418
rect 39954 28366 39966 28418
rect 40898 28366 40910 28418
rect 40962 28366 40974 28418
rect 47506 28366 47518 28418
rect 47570 28366 47582 28418
rect 50082 28366 50094 28418
rect 50146 28415 50158 28418
rect 50978 28415 50990 28418
rect 50146 28369 50990 28415
rect 50146 28366 50158 28369
rect 50978 28366 50990 28369
rect 51042 28366 51054 28418
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 1810 28030 1822 28082
rect 1874 28079 1886 28082
rect 2370 28079 2382 28082
rect 1874 28033 2382 28079
rect 1874 28030 1886 28033
rect 2370 28030 2382 28033
rect 2434 28030 2446 28082
rect 2594 28030 2606 28082
rect 2658 28030 2670 28082
rect 18498 28030 18510 28082
rect 18562 28030 18574 28082
rect 25330 28030 25342 28082
rect 25394 28030 25406 28082
rect 27010 28030 27022 28082
rect 27074 28030 27086 28082
rect 31154 28030 31166 28082
rect 31218 28030 31230 28082
rect 33506 28030 33518 28082
rect 33570 28030 33582 28082
rect 36194 28030 36206 28082
rect 36258 28030 36270 28082
rect 48850 28030 48862 28082
rect 48914 28079 48926 28082
rect 50194 28079 50206 28082
rect 48914 28033 50206 28079
rect 48914 28030 48926 28033
rect 50194 28030 50206 28033
rect 50258 28030 50270 28082
rect 3166 27970 3218 27982
rect 3166 27906 3218 27918
rect 3614 27970 3666 27982
rect 3614 27906 3666 27918
rect 14254 27970 14306 27982
rect 14254 27906 14306 27918
rect 14702 27970 14754 27982
rect 27806 27970 27858 27982
rect 26898 27918 26910 27970
rect 26962 27918 26974 27970
rect 14702 27906 14754 27918
rect 27806 27906 27858 27918
rect 28478 27970 28530 27982
rect 28478 27906 28530 27918
rect 29710 27970 29762 27982
rect 29710 27906 29762 27918
rect 30718 27970 30770 27982
rect 30718 27906 30770 27918
rect 34414 27970 34466 27982
rect 34414 27906 34466 27918
rect 37886 27970 37938 27982
rect 37886 27906 37938 27918
rect 39230 27970 39282 27982
rect 39230 27906 39282 27918
rect 42142 27970 42194 27982
rect 42142 27906 42194 27918
rect 42814 27970 42866 27982
rect 42814 27906 42866 27918
rect 43262 27970 43314 27982
rect 43262 27906 43314 27918
rect 44718 27970 44770 27982
rect 44718 27906 44770 27918
rect 45166 27970 45218 27982
rect 45166 27906 45218 27918
rect 45614 27970 45666 27982
rect 45614 27906 45666 27918
rect 46062 27970 46114 27982
rect 46062 27906 46114 27918
rect 46846 27970 46898 27982
rect 46846 27906 46898 27918
rect 48862 27970 48914 27982
rect 48862 27906 48914 27918
rect 49310 27970 49362 27982
rect 49310 27906 49362 27918
rect 50206 27970 50258 27982
rect 50206 27906 50258 27918
rect 50654 27970 50706 27982
rect 50654 27906 50706 27918
rect 53118 27970 53170 27982
rect 54786 27918 54798 27970
rect 54850 27918 54862 27970
rect 55346 27918 55358 27970
rect 55410 27918 55422 27970
rect 53118 27906 53170 27918
rect 1822 27858 1874 27870
rect 1822 27794 1874 27806
rect 2270 27858 2322 27870
rect 2270 27794 2322 27806
rect 16046 27858 16098 27870
rect 16046 27794 16098 27806
rect 18958 27858 19010 27870
rect 18958 27794 19010 27806
rect 19406 27858 19458 27870
rect 19406 27794 19458 27806
rect 25902 27858 25954 27870
rect 25902 27794 25954 27806
rect 26126 27858 26178 27870
rect 26126 27794 26178 27806
rect 27134 27858 27186 27870
rect 27134 27794 27186 27806
rect 27358 27858 27410 27870
rect 27358 27794 27410 27806
rect 28142 27858 28194 27870
rect 28142 27794 28194 27806
rect 28814 27858 28866 27870
rect 28814 27794 28866 27806
rect 30046 27858 30098 27870
rect 30046 27794 30098 27806
rect 30382 27858 30434 27870
rect 30382 27794 30434 27806
rect 31502 27858 31554 27870
rect 31502 27794 31554 27806
rect 32062 27858 32114 27870
rect 32062 27794 32114 27806
rect 33070 27858 33122 27870
rect 33070 27794 33122 27806
rect 33406 27858 33458 27870
rect 33406 27794 33458 27806
rect 33518 27858 33570 27870
rect 33518 27794 33570 27806
rect 33854 27858 33906 27870
rect 35982 27858 36034 27870
rect 36542 27858 36594 27870
rect 35522 27806 35534 27858
rect 35586 27806 35598 27858
rect 36306 27806 36318 27858
rect 36370 27806 36382 27858
rect 33854 27794 33906 27806
rect 35982 27794 36034 27806
rect 36542 27794 36594 27806
rect 36766 27858 36818 27870
rect 40014 27858 40066 27870
rect 39666 27806 39678 27858
rect 39730 27806 39742 27858
rect 36766 27794 36818 27806
rect 40014 27794 40066 27806
rect 41358 27858 41410 27870
rect 47182 27858 47234 27870
rect 46498 27806 46510 27858
rect 46562 27806 46574 27858
rect 41358 27794 41410 27806
rect 47182 27794 47234 27806
rect 48190 27858 48242 27870
rect 48190 27794 48242 27806
rect 51102 27858 51154 27870
rect 51102 27794 51154 27806
rect 51662 27858 51714 27870
rect 51662 27794 51714 27806
rect 52110 27858 52162 27870
rect 52110 27794 52162 27806
rect 52334 27858 52386 27870
rect 52334 27794 52386 27806
rect 53454 27858 53506 27870
rect 53454 27794 53506 27806
rect 54350 27858 54402 27870
rect 54898 27806 54910 27858
rect 54962 27806 54974 27858
rect 55794 27806 55806 27858
rect 55858 27806 55870 27858
rect 54350 27794 54402 27806
rect 6302 27746 6354 27758
rect 2706 27694 2718 27746
rect 2770 27694 2782 27746
rect 5730 27694 5742 27746
rect 5794 27694 5806 27746
rect 6302 27682 6354 27694
rect 11566 27746 11618 27758
rect 15486 27746 15538 27758
rect 25678 27746 25730 27758
rect 12114 27694 12126 27746
rect 12178 27694 12190 27746
rect 15698 27694 15710 27746
rect 15762 27694 15774 27746
rect 19506 27694 19518 27746
rect 19570 27694 19582 27746
rect 11566 27682 11618 27694
rect 15486 27682 15538 27694
rect 25678 27682 25730 27694
rect 26350 27746 26402 27758
rect 26350 27682 26402 27694
rect 26574 27746 26626 27758
rect 37326 27746 37378 27758
rect 34178 27694 34190 27746
rect 34242 27694 34254 27746
rect 26574 27682 26626 27694
rect 37326 27682 37378 27694
rect 37550 27746 37602 27758
rect 37550 27682 37602 27694
rect 37774 27746 37826 27758
rect 37774 27682 37826 27694
rect 37998 27746 38050 27758
rect 39790 27746 39842 27758
rect 39106 27694 39118 27746
rect 39170 27694 39182 27746
rect 37998 27682 38050 27694
rect 39790 27682 39842 27694
rect 40910 27746 40962 27758
rect 53342 27746 53394 27758
rect 42242 27694 42254 27746
rect 42306 27694 42318 27746
rect 51874 27694 51886 27746
rect 51938 27694 51950 27746
rect 40910 27682 40962 27694
rect 53342 27682 53394 27694
rect 11230 27634 11282 27646
rect 11230 27570 11282 27582
rect 25454 27634 25506 27646
rect 25454 27570 25506 27582
rect 29262 27634 29314 27646
rect 29262 27570 29314 27582
rect 31838 27634 31890 27646
rect 31838 27570 31890 27582
rect 32510 27634 32562 27646
rect 32510 27570 32562 27582
rect 38446 27634 38498 27646
rect 38446 27570 38498 27582
rect 40238 27634 40290 27646
rect 43710 27634 43762 27646
rect 40338 27582 40350 27634
rect 40402 27582 40414 27634
rect 40238 27570 40290 27582
rect 43710 27570 43762 27582
rect 46286 27634 46338 27646
rect 46286 27570 46338 27582
rect 49758 27634 49810 27646
rect 56702 27634 56754 27646
rect 51874 27631 51886 27634
rect 49758 27570 49810 27582
rect 51441 27585 51886 27631
rect 31726 27522 31778 27534
rect 31726 27458 31778 27470
rect 41022 27522 41074 27534
rect 41022 27458 41074 27470
rect 47854 27522 47906 27534
rect 48962 27470 48974 27522
rect 49026 27519 49038 27522
rect 49858 27519 49870 27522
rect 49026 27473 49870 27519
rect 49026 27470 49038 27473
rect 49858 27470 49870 27473
rect 49922 27519 49934 27522
rect 50082 27519 50094 27522
rect 49922 27473 50094 27519
rect 49922 27470 49934 27473
rect 50082 27470 50094 27473
rect 50146 27519 50158 27522
rect 51441 27519 51487 27585
rect 51874 27582 51886 27585
rect 51938 27582 51950 27634
rect 56702 27570 56754 27582
rect 50146 27473 51487 27519
rect 51998 27522 52050 27534
rect 50146 27470 50158 27473
rect 47854 27458 47906 27470
rect 51998 27458 52050 27470
rect 15026 27358 15038 27410
rect 15090 27358 15102 27410
rect 1344 27242 58576 27276
rect 1344 27190 4478 27242
rect 4530 27190 4582 27242
rect 4634 27190 4686 27242
rect 4738 27190 35198 27242
rect 35250 27190 35302 27242
rect 35354 27190 35406 27242
rect 35458 27190 58576 27242
rect 1344 27156 58576 27190
rect 37426 27022 37438 27074
rect 37490 27022 37502 27074
rect 35298 26910 35310 26962
rect 35362 26910 35374 26962
rect 4958 26850 5010 26862
rect 4958 26786 5010 26798
rect 9326 26850 9378 26862
rect 9326 26786 9378 26798
rect 23438 26850 23490 26862
rect 23438 26786 23490 26798
rect 24558 26850 24610 26862
rect 24558 26786 24610 26798
rect 26126 26850 26178 26862
rect 33518 26850 33570 26862
rect 39006 26850 39058 26862
rect 28130 26798 28142 26850
rect 28194 26798 28206 26850
rect 36306 26798 36318 26850
rect 36370 26798 36382 26850
rect 26126 26786 26178 26798
rect 33518 26786 33570 26798
rect 39006 26786 39058 26798
rect 43374 26850 43426 26862
rect 43374 26786 43426 26798
rect 44270 26850 44322 26862
rect 44270 26786 44322 26798
rect 44718 26850 44770 26862
rect 44718 26786 44770 26798
rect 46398 26850 46450 26862
rect 46398 26786 46450 26798
rect 50654 26850 50706 26862
rect 50654 26786 50706 26798
rect 1822 26738 1874 26750
rect 12910 26738 12962 26750
rect 2370 26686 2382 26738
rect 2434 26686 2446 26738
rect 12338 26686 12350 26738
rect 12402 26686 12414 26738
rect 1822 26674 1874 26686
rect 12910 26674 12962 26686
rect 13470 26738 13522 26750
rect 28478 26738 28530 26750
rect 14018 26686 14030 26738
rect 14082 26686 14094 26738
rect 13470 26674 13522 26686
rect 28478 26674 28530 26686
rect 30830 26738 30882 26750
rect 30830 26674 30882 26686
rect 33070 26738 33122 26750
rect 34190 26738 34242 26750
rect 33730 26686 33742 26738
rect 33794 26686 33806 26738
rect 33070 26674 33122 26686
rect 34190 26674 34242 26686
rect 34750 26738 34802 26750
rect 35646 26738 35698 26750
rect 35074 26686 35086 26738
rect 35138 26686 35150 26738
rect 34750 26674 34802 26686
rect 35646 26674 35698 26686
rect 37102 26738 37154 26750
rect 37102 26674 37154 26686
rect 37326 26738 37378 26750
rect 37326 26674 37378 26686
rect 37550 26738 37602 26750
rect 37550 26674 37602 26686
rect 37774 26738 37826 26750
rect 37774 26674 37826 26686
rect 38894 26738 38946 26750
rect 38894 26674 38946 26686
rect 39342 26738 39394 26750
rect 39342 26674 39394 26686
rect 39790 26738 39842 26750
rect 39790 26674 39842 26686
rect 40238 26738 40290 26750
rect 49758 26738 49810 26750
rect 40562 26686 40574 26738
rect 40626 26686 40638 26738
rect 42130 26686 42142 26738
rect 42194 26686 42206 26738
rect 45490 26686 45502 26738
rect 45554 26686 45566 26738
rect 46834 26686 46846 26738
rect 46898 26686 46910 26738
rect 40238 26674 40290 26686
rect 49758 26674 49810 26686
rect 51326 26738 51378 26750
rect 52670 26738 52722 26750
rect 51538 26686 51550 26738
rect 51602 26686 51614 26738
rect 51326 26674 51378 26686
rect 52670 26674 52722 26686
rect 53006 26738 53058 26750
rect 53006 26674 53058 26686
rect 53678 26738 53730 26750
rect 53678 26674 53730 26686
rect 54238 26738 54290 26750
rect 54238 26674 54290 26686
rect 54798 26738 54850 26750
rect 54798 26674 54850 26686
rect 9774 26626 9826 26638
rect 9774 26562 9826 26574
rect 23550 26626 23602 26638
rect 23550 26562 23602 26574
rect 24110 26626 24162 26638
rect 24110 26562 24162 26574
rect 26686 26626 26738 26638
rect 26686 26562 26738 26574
rect 27022 26626 27074 26638
rect 27022 26562 27074 26574
rect 27358 26626 27410 26638
rect 27358 26562 27410 26574
rect 27918 26626 27970 26638
rect 27918 26562 27970 26574
rect 28254 26626 28306 26638
rect 39118 26626 39170 26638
rect 31266 26574 31278 26626
rect 31330 26574 31342 26626
rect 31602 26574 31614 26626
rect 31666 26574 31678 26626
rect 35970 26574 35982 26626
rect 36034 26574 36046 26626
rect 28254 26562 28306 26574
rect 39118 26562 39170 26574
rect 40798 26626 40850 26638
rect 40798 26562 40850 26574
rect 41694 26626 41746 26638
rect 41694 26562 41746 26574
rect 42254 26626 42306 26638
rect 42254 26562 42306 26574
rect 42926 26626 42978 26638
rect 42926 26562 42978 26574
rect 45166 26626 45218 26638
rect 45166 26562 45218 26574
rect 45614 26626 45666 26638
rect 45614 26562 45666 26574
rect 50878 26626 50930 26638
rect 50878 26562 50930 26574
rect 51886 26626 51938 26638
rect 51886 26562 51938 26574
rect 53342 26626 53394 26638
rect 53342 26562 53394 26574
rect 4510 26514 4562 26526
rect 16158 26514 16210 26526
rect 10098 26462 10110 26514
rect 10162 26462 10174 26514
rect 4510 26450 4562 26462
rect 16158 26450 16210 26462
rect 16606 26514 16658 26526
rect 16606 26450 16658 26462
rect 20750 26514 20802 26526
rect 20750 26450 20802 26462
rect 21422 26514 21474 26526
rect 21422 26450 21474 26462
rect 21870 26514 21922 26526
rect 21870 26450 21922 26462
rect 24894 26514 24946 26526
rect 24894 26450 24946 26462
rect 26350 26514 26402 26526
rect 26350 26450 26402 26462
rect 27470 26514 27522 26526
rect 27470 26450 27522 26462
rect 29598 26514 29650 26526
rect 29598 26450 29650 26462
rect 30046 26514 30098 26526
rect 30046 26450 30098 26462
rect 30494 26514 30546 26526
rect 38334 26514 38386 26526
rect 30930 26462 30942 26514
rect 30994 26462 31006 26514
rect 30494 26450 30546 26462
rect 38334 26450 38386 26462
rect 43934 26514 43986 26526
rect 50206 26514 50258 26526
rect 46274 26462 46286 26514
rect 46338 26462 46350 26514
rect 43934 26450 43986 26462
rect 27346 26350 27358 26402
rect 27410 26350 27422 26402
rect 41234 26350 41246 26402
rect 41298 26350 41310 26402
rect 46289 26399 46335 26462
rect 50206 26450 50258 26462
rect 55470 26514 55522 26526
rect 55470 26450 55522 26462
rect 46498 26399 46510 26402
rect 46289 26353 46510 26399
rect 46498 26350 46510 26353
rect 46562 26350 46574 26402
rect 47282 26350 47294 26402
rect 47346 26350 47358 26402
rect 49634 26350 49646 26402
rect 49698 26399 49710 26402
rect 50642 26399 50654 26402
rect 49698 26353 50654 26399
rect 49698 26350 49710 26353
rect 50642 26350 50654 26353
rect 50706 26350 50718 26402
rect 1344 26234 58576 26268
rect 1344 26182 19838 26234
rect 19890 26182 19942 26234
rect 19994 26182 20046 26234
rect 20098 26182 50558 26234
rect 50610 26182 50662 26234
rect 50714 26182 50766 26234
rect 50818 26182 58576 26234
rect 1344 26148 58576 26182
rect 30258 26014 30270 26066
rect 30322 26063 30334 26066
rect 30818 26063 30830 26066
rect 30322 26017 30830 26063
rect 30322 26014 30334 26017
rect 30818 26014 30830 26017
rect 30882 26014 30894 26066
rect 35746 26014 35758 26066
rect 35810 26014 35822 26066
rect 44818 26014 44830 26066
rect 44882 26014 44894 26066
rect 1822 25954 1874 25966
rect 1822 25890 1874 25902
rect 2718 25954 2770 25966
rect 10558 25954 10610 25966
rect 4946 25902 4958 25954
rect 5010 25902 5022 25954
rect 2718 25890 2770 25902
rect 10558 25890 10610 25902
rect 11006 25954 11058 25966
rect 11006 25890 11058 25902
rect 11454 25954 11506 25966
rect 14926 25954 14978 25966
rect 14578 25902 14590 25954
rect 14642 25902 14654 25954
rect 11454 25890 11506 25902
rect 14926 25890 14978 25902
rect 22206 25954 22258 25966
rect 22206 25890 22258 25902
rect 25566 25954 25618 25966
rect 25566 25890 25618 25902
rect 25902 25954 25954 25966
rect 25902 25890 25954 25902
rect 30270 25954 30322 25966
rect 30270 25890 30322 25902
rect 37886 25954 37938 25966
rect 37886 25890 37938 25902
rect 38782 25954 38834 25966
rect 42142 25954 42194 25966
rect 55358 25954 55410 25966
rect 41458 25902 41470 25954
rect 41522 25902 41534 25954
rect 53330 25902 53342 25954
rect 53394 25902 53406 25954
rect 38782 25890 38834 25902
rect 42142 25890 42194 25902
rect 55358 25890 55410 25902
rect 55806 25954 55858 25966
rect 55806 25890 55858 25902
rect 56702 25954 56754 25966
rect 56702 25890 56754 25902
rect 23998 25842 24050 25854
rect 23998 25778 24050 25790
rect 29710 25842 29762 25854
rect 32510 25842 32562 25854
rect 31378 25790 31390 25842
rect 31442 25790 31454 25842
rect 29710 25778 29762 25790
rect 32510 25778 32562 25790
rect 33294 25842 33346 25854
rect 35758 25842 35810 25854
rect 35522 25790 35534 25842
rect 35586 25790 35598 25842
rect 33294 25778 33346 25790
rect 35758 25778 35810 25790
rect 35982 25842 36034 25854
rect 35982 25778 36034 25790
rect 36766 25842 36818 25854
rect 36766 25778 36818 25790
rect 37550 25842 37602 25854
rect 37550 25778 37602 25790
rect 38670 25842 38722 25854
rect 38670 25778 38722 25790
rect 40126 25842 40178 25854
rect 43822 25842 43874 25854
rect 42354 25790 42366 25842
rect 42418 25790 42430 25842
rect 40126 25778 40178 25790
rect 43822 25778 43874 25790
rect 45390 25842 45442 25854
rect 45390 25778 45442 25790
rect 45726 25842 45778 25854
rect 47182 25842 47234 25854
rect 46498 25790 46510 25842
rect 46562 25790 46574 25842
rect 45726 25778 45778 25790
rect 47182 25778 47234 25790
rect 47854 25842 47906 25854
rect 53902 25842 53954 25854
rect 49634 25790 49646 25842
rect 49698 25790 49710 25842
rect 47854 25778 47906 25790
rect 53902 25778 53954 25790
rect 7758 25730 7810 25742
rect 11790 25730 11842 25742
rect 17838 25730 17890 25742
rect 3042 25678 3054 25730
rect 3106 25678 3118 25730
rect 3602 25678 3614 25730
rect 3666 25678 3678 25730
rect 4050 25678 4062 25730
rect 4114 25678 4126 25730
rect 7186 25678 7198 25730
rect 7250 25678 7262 25730
rect 8194 25678 8206 25730
rect 8258 25678 8270 25730
rect 8754 25678 8766 25730
rect 8818 25678 8830 25730
rect 12338 25678 12350 25730
rect 12402 25678 12414 25730
rect 17490 25678 17502 25730
rect 17554 25678 17566 25730
rect 7758 25666 7810 25678
rect 11790 25666 11842 25678
rect 17838 25666 17890 25678
rect 19966 25730 20018 25742
rect 19966 25666 20018 25678
rect 20750 25730 20802 25742
rect 20750 25666 20802 25678
rect 21198 25730 21250 25742
rect 21198 25666 21250 25678
rect 21534 25730 21586 25742
rect 21534 25666 21586 25678
rect 21870 25730 21922 25742
rect 21870 25666 21922 25678
rect 22766 25730 22818 25742
rect 22766 25666 22818 25678
rect 23326 25730 23378 25742
rect 23326 25666 23378 25678
rect 26238 25730 26290 25742
rect 26238 25666 26290 25678
rect 26462 25730 26514 25742
rect 28366 25741 28418 25753
rect 27010 25678 27022 25730
rect 27074 25678 27086 25730
rect 26462 25666 26514 25678
rect 28366 25677 28418 25689
rect 28590 25730 28642 25742
rect 28590 25666 28642 25678
rect 28814 25730 28866 25742
rect 28814 25666 28866 25678
rect 29038 25730 29090 25742
rect 29038 25666 29090 25678
rect 29486 25730 29538 25742
rect 29486 25666 29538 25678
rect 29598 25730 29650 25742
rect 29598 25666 29650 25678
rect 30718 25730 30770 25742
rect 30718 25666 30770 25678
rect 31166 25730 31218 25742
rect 31166 25666 31218 25678
rect 31726 25730 31778 25742
rect 31726 25666 31778 25678
rect 32174 25730 32226 25742
rect 32174 25666 32226 25678
rect 32286 25730 32338 25742
rect 32286 25666 32338 25678
rect 34078 25730 34130 25742
rect 34526 25730 34578 25742
rect 34178 25678 34190 25730
rect 34242 25678 34254 25730
rect 34078 25666 34130 25678
rect 34526 25666 34578 25678
rect 34862 25730 34914 25742
rect 34862 25666 34914 25678
rect 35198 25730 35250 25742
rect 35198 25666 35250 25678
rect 36542 25730 36594 25742
rect 36542 25666 36594 25678
rect 36654 25730 36706 25742
rect 36654 25666 36706 25678
rect 36990 25730 37042 25742
rect 36990 25666 37042 25678
rect 37214 25730 37266 25742
rect 37214 25666 37266 25678
rect 38446 25730 38498 25742
rect 38446 25666 38498 25678
rect 38894 25730 38946 25742
rect 38894 25666 38946 25678
rect 39566 25730 39618 25742
rect 44382 25730 44434 25742
rect 41234 25678 41246 25730
rect 41298 25678 41310 25730
rect 42018 25678 42030 25730
rect 42082 25678 42094 25730
rect 39566 25666 39618 25678
rect 44382 25666 44434 25678
rect 45054 25730 45106 25742
rect 45054 25666 45106 25678
rect 46062 25730 46114 25742
rect 46062 25666 46114 25678
rect 49086 25730 49138 25742
rect 49086 25666 49138 25678
rect 50990 25730 51042 25742
rect 54910 25730 54962 25742
rect 52210 25678 52222 25730
rect 52274 25678 52286 25730
rect 53218 25678 53230 25730
rect 53282 25678 53294 25730
rect 50990 25666 51042 25678
rect 54910 25666 54962 25678
rect 3950 25618 4002 25630
rect 3950 25554 4002 25566
rect 16830 25618 16882 25630
rect 16830 25554 16882 25566
rect 28030 25618 28082 25630
rect 28030 25554 28082 25566
rect 31390 25618 31442 25630
rect 31390 25554 31442 25566
rect 40238 25618 40290 25630
rect 43710 25618 43762 25630
rect 41682 25566 41694 25618
rect 41746 25566 41758 25618
rect 40238 25554 40290 25566
rect 43710 25554 43762 25566
rect 57150 25618 57202 25630
rect 57150 25554 57202 25566
rect 26910 25506 26962 25518
rect 4610 25454 4622 25506
rect 4674 25454 4686 25506
rect 26910 25442 26962 25454
rect 33630 25506 33682 25518
rect 33630 25442 33682 25454
rect 3154 25342 3166 25394
rect 3218 25342 3230 25394
rect 3490 25342 3502 25394
rect 3554 25342 3566 25394
rect 8082 25342 8094 25394
rect 8146 25342 8158 25394
rect 8866 25342 8878 25394
rect 8930 25342 8942 25394
rect 10882 25342 10894 25394
rect 10946 25342 10958 25394
rect 11330 25342 11342 25394
rect 11394 25342 11406 25394
rect 28690 25342 28702 25394
rect 28754 25342 28766 25394
rect 39106 25342 39118 25394
rect 39170 25342 39182 25394
rect 1344 25226 58576 25260
rect 1344 25174 4478 25226
rect 4530 25174 4582 25226
rect 4634 25174 4686 25226
rect 4738 25174 35198 25226
rect 35250 25174 35302 25226
rect 35354 25174 35406 25226
rect 35458 25174 58576 25226
rect 1344 25140 58576 25174
rect 5730 25006 5742 25058
rect 5794 25006 5806 25058
rect 13458 25006 13470 25058
rect 13522 25006 13534 25058
rect 32498 25006 32510 25058
rect 32562 25006 32574 25058
rect 53218 25006 53230 25058
rect 53282 25055 53294 25058
rect 53778 25055 53790 25058
rect 53282 25009 53790 25055
rect 53282 25006 53294 25009
rect 53778 25006 53790 25009
rect 53842 25006 53854 25058
rect 4946 24894 4958 24946
rect 5010 24894 5022 24946
rect 6178 24894 6190 24946
rect 6242 24894 6254 24946
rect 12786 24894 12798 24946
rect 12850 24894 12862 24946
rect 20514 24894 20526 24946
rect 20578 24894 20590 24946
rect 19406 24834 19458 24846
rect 27022 24834 27074 24846
rect 24098 24782 24110 24834
rect 24162 24782 24174 24834
rect 19406 24770 19458 24782
rect 27022 24770 27074 24782
rect 28142 24834 28194 24846
rect 28142 24770 28194 24782
rect 29486 24834 29538 24846
rect 29486 24770 29538 24782
rect 31614 24834 31666 24846
rect 31614 24770 31666 24782
rect 34190 24834 34242 24846
rect 34190 24770 34242 24782
rect 45278 24834 45330 24846
rect 1822 24722 1874 24734
rect 9326 24722 9378 24734
rect 2370 24670 2382 24722
rect 2434 24670 2446 24722
rect 5618 24670 5630 24722
rect 5682 24670 5694 24722
rect 8754 24670 8766 24722
rect 8818 24670 8830 24722
rect 1822 24658 1874 24670
rect 9326 24658 9378 24670
rect 9662 24722 9714 24734
rect 16270 24722 16322 24734
rect 19070 24722 19122 24734
rect 10210 24670 10222 24722
rect 10274 24670 10286 24722
rect 13570 24670 13582 24722
rect 13634 24670 13646 24722
rect 16706 24670 16718 24722
rect 16770 24670 16782 24722
rect 9662 24658 9714 24670
rect 16270 24658 16322 24670
rect 19070 24658 19122 24670
rect 21422 24722 21474 24734
rect 21422 24658 21474 24670
rect 21982 24722 22034 24734
rect 21982 24658 22034 24670
rect 25566 24722 25618 24734
rect 25566 24658 25618 24670
rect 27694 24722 27746 24734
rect 29822 24722 29874 24734
rect 29138 24670 29150 24722
rect 29202 24670 29214 24722
rect 27694 24658 27746 24670
rect 29822 24658 29874 24670
rect 32398 24722 32450 24734
rect 32398 24658 32450 24670
rect 32622 24722 32674 24734
rect 35646 24722 35698 24734
rect 35186 24670 35198 24722
rect 35250 24670 35262 24722
rect 32622 24658 32674 24670
rect 35646 24658 35698 24670
rect 35870 24722 35922 24734
rect 35870 24658 35922 24670
rect 36878 24722 36930 24734
rect 36878 24658 36930 24670
rect 39118 24722 39170 24734
rect 39118 24658 39170 24670
rect 39230 24722 39282 24734
rect 39230 24658 39282 24670
rect 39566 24722 39618 24734
rect 39566 24658 39618 24670
rect 41694 24722 41746 24734
rect 42354 24726 42366 24778
rect 42418 24726 42430 24778
rect 45278 24770 45330 24782
rect 45726 24834 45778 24846
rect 52782 24834 52834 24846
rect 47842 24782 47854 24834
rect 47906 24782 47918 24834
rect 45726 24770 45778 24782
rect 52782 24770 52834 24782
rect 53230 24834 53282 24846
rect 53230 24770 53282 24782
rect 53678 24834 53730 24846
rect 55346 24782 55358 24834
rect 55410 24782 55422 24834
rect 53678 24770 53730 24782
rect 56702 24722 56754 24734
rect 49522 24670 49534 24722
rect 49586 24670 49598 24722
rect 54450 24670 54462 24722
rect 54514 24670 54526 24722
rect 55794 24670 55806 24722
rect 55858 24670 55870 24722
rect 41694 24658 41746 24670
rect 24894 24610 24946 24622
rect 24894 24546 24946 24558
rect 25006 24610 25058 24622
rect 25006 24546 25058 24558
rect 26238 24610 26290 24622
rect 26238 24546 26290 24558
rect 27470 24610 27522 24622
rect 27470 24546 27522 24558
rect 34862 24610 34914 24622
rect 34862 24546 34914 24558
rect 37550 24610 37602 24622
rect 37550 24546 37602 24558
rect 37774 24610 37826 24622
rect 37774 24546 37826 24558
rect 38446 24610 38498 24622
rect 38446 24546 38498 24558
rect 39342 24610 39394 24622
rect 39342 24546 39394 24558
rect 41246 24610 41298 24622
rect 41246 24546 41298 24558
rect 42814 24610 42866 24622
rect 50642 24614 50654 24666
rect 50706 24614 50718 24666
rect 56702 24658 56754 24670
rect 57822 24722 57874 24734
rect 57822 24658 57874 24670
rect 58046 24710 58098 24722
rect 58046 24646 58098 24658
rect 42814 24546 42866 24558
rect 57598 24610 57650 24622
rect 57598 24546 57650 24558
rect 12350 24498 12402 24510
rect 4610 24446 4622 24498
rect 4674 24446 4686 24498
rect 6514 24446 6526 24498
rect 6578 24446 6590 24498
rect 12350 24434 12402 24446
rect 14030 24498 14082 24510
rect 14030 24434 14082 24446
rect 26574 24498 26626 24510
rect 29710 24498 29762 24510
rect 29250 24446 29262 24498
rect 29314 24446 29326 24498
rect 26574 24434 26626 24446
rect 29710 24434 29762 24446
rect 32062 24498 32114 24510
rect 32062 24434 32114 24446
rect 32846 24498 32898 24510
rect 32846 24434 32898 24446
rect 33294 24498 33346 24510
rect 33294 24434 33346 24446
rect 33742 24498 33794 24510
rect 33742 24434 33794 24446
rect 34526 24498 34578 24510
rect 38110 24498 38162 24510
rect 36194 24446 36206 24498
rect 36258 24446 36270 24498
rect 37202 24446 37214 24498
rect 37266 24446 37278 24498
rect 34526 24434 34578 24446
rect 38110 24434 38162 24446
rect 40126 24498 40178 24510
rect 51214 24498 51266 24510
rect 40562 24446 40574 24498
rect 40626 24446 40638 24498
rect 40126 24434 40178 24446
rect 51214 24434 51266 24446
rect 51886 24498 51938 24510
rect 51886 24434 51938 24446
rect 2482 24334 2494 24386
rect 2546 24383 2558 24386
rect 3042 24383 3054 24386
rect 2546 24337 3054 24383
rect 2546 24334 2558 24337
rect 3042 24334 3054 24337
rect 3106 24334 3118 24386
rect 26002 24334 26014 24386
rect 26066 24334 26078 24386
rect 27570 24334 27582 24386
rect 27634 24334 27646 24386
rect 37426 24334 37438 24386
rect 37490 24334 37502 24386
rect 52546 24334 52558 24386
rect 52610 24383 52622 24386
rect 53554 24383 53566 24386
rect 52610 24337 53566 24383
rect 52610 24334 52622 24337
rect 53554 24334 53566 24337
rect 53618 24334 53630 24386
rect 54114 24334 54126 24386
rect 54178 24334 54190 24386
rect 57474 24334 57486 24386
rect 57538 24334 57550 24386
rect 1344 24218 58576 24252
rect 1344 24166 19838 24218
rect 19890 24166 19942 24218
rect 19994 24166 20046 24218
rect 20098 24166 50558 24218
rect 50610 24166 50662 24218
rect 50714 24166 50766 24218
rect 50818 24166 58576 24218
rect 1344 24132 58576 24166
rect 22082 23998 22094 24050
rect 22146 24047 22158 24050
rect 22978 24047 22990 24050
rect 22146 24001 22990 24047
rect 22146 23998 22158 24001
rect 22978 23998 22990 24001
rect 23042 23998 23054 24050
rect 32050 23998 32062 24050
rect 32114 23998 32126 24050
rect 36082 23998 36094 24050
rect 36146 23998 36158 24050
rect 36978 23998 36990 24050
rect 37042 23998 37054 24050
rect 39218 23998 39230 24050
rect 39282 24047 39294 24050
rect 39282 24001 40063 24047
rect 39282 23998 39294 24001
rect 1822 23938 1874 23950
rect 1822 23874 1874 23886
rect 2270 23938 2322 23950
rect 5854 23938 5906 23950
rect 9662 23938 9714 23950
rect 2594 23886 2606 23938
rect 2658 23886 2670 23938
rect 6178 23886 6190 23938
rect 6242 23886 6254 23938
rect 2270 23874 2322 23886
rect 5854 23874 5906 23886
rect 9662 23874 9714 23886
rect 21422 23938 21474 23950
rect 21422 23874 21474 23886
rect 22094 23938 22146 23950
rect 22094 23874 22146 23886
rect 22990 23938 23042 23950
rect 22990 23874 23042 23886
rect 24558 23938 24610 23950
rect 24558 23874 24610 23886
rect 25566 23938 25618 23950
rect 25566 23874 25618 23886
rect 26574 23938 26626 23950
rect 26574 23874 26626 23886
rect 26686 23938 26738 23950
rect 26686 23874 26738 23886
rect 28254 23938 28306 23950
rect 28254 23874 28306 23886
rect 33182 23938 33234 23950
rect 33182 23874 33234 23886
rect 34190 23938 34242 23950
rect 34190 23874 34242 23886
rect 34302 23938 34354 23950
rect 34302 23874 34354 23886
rect 35086 23938 35138 23950
rect 35086 23874 35138 23886
rect 35870 23938 35922 23950
rect 37662 23938 37714 23950
rect 36754 23886 36766 23938
rect 36818 23886 36830 23938
rect 35870 23874 35922 23886
rect 37662 23874 37714 23886
rect 38558 23938 38610 23950
rect 38558 23874 38610 23886
rect 39342 23938 39394 23950
rect 39342 23874 39394 23886
rect 39790 23938 39842 23950
rect 40017 23938 40063 24001
rect 40238 23938 40290 23950
rect 40002 23886 40014 23938
rect 40066 23886 40078 23938
rect 39790 23874 39842 23886
rect 40238 23874 40290 23886
rect 43934 23938 43986 23950
rect 43934 23874 43986 23886
rect 44382 23938 44434 23950
rect 47630 23938 47682 23950
rect 45042 23886 45054 23938
rect 45106 23886 45118 23938
rect 44382 23874 44434 23886
rect 47630 23874 47682 23886
rect 48078 23938 48130 23950
rect 48078 23874 48130 23886
rect 49982 23938 50034 23950
rect 49982 23874 50034 23886
rect 53902 23938 53954 23950
rect 53902 23874 53954 23886
rect 55694 23938 55746 23950
rect 55694 23874 55746 23886
rect 57150 23938 57202 23950
rect 57150 23874 57202 23886
rect 17614 23826 17666 23838
rect 17614 23762 17666 23774
rect 25342 23826 25394 23838
rect 26350 23826 26402 23838
rect 25778 23774 25790 23826
rect 25842 23774 25854 23826
rect 25342 23762 25394 23774
rect 26350 23762 26402 23774
rect 28702 23826 28754 23838
rect 28702 23762 28754 23774
rect 28926 23826 28978 23838
rect 28926 23762 28978 23774
rect 30942 23826 30994 23838
rect 30942 23762 30994 23774
rect 35422 23826 35474 23838
rect 35422 23762 35474 23774
rect 35758 23826 35810 23838
rect 35758 23762 35810 23774
rect 36542 23826 36594 23838
rect 36542 23762 36594 23774
rect 37102 23826 37154 23838
rect 37102 23762 37154 23774
rect 37326 23826 37378 23838
rect 37326 23762 37378 23774
rect 38894 23826 38946 23838
rect 42478 23826 42530 23838
rect 48862 23826 48914 23838
rect 42242 23774 42254 23826
rect 42306 23774 42318 23826
rect 46050 23774 46062 23826
rect 46114 23774 46126 23826
rect 46386 23774 46398 23826
rect 46450 23774 46462 23826
rect 38894 23762 38946 23774
rect 42478 23762 42530 23774
rect 48862 23762 48914 23774
rect 50654 23826 50706 23838
rect 50654 23762 50706 23774
rect 52894 23826 52946 23838
rect 52894 23762 52946 23774
rect 53230 23826 53282 23838
rect 53230 23762 53282 23774
rect 53566 23826 53618 23838
rect 54338 23774 54350 23826
rect 54402 23774 54414 23826
rect 53566 23762 53618 23774
rect 5406 23714 5458 23726
rect 8990 23714 9042 23726
rect 4834 23662 4846 23714
rect 4898 23662 4910 23714
rect 8418 23662 8430 23714
rect 8482 23662 8494 23714
rect 5406 23650 5458 23662
rect 8990 23650 9042 23662
rect 17950 23714 18002 23726
rect 18846 23714 18898 23726
rect 18498 23662 18510 23714
rect 18562 23662 18574 23714
rect 17950 23650 18002 23662
rect 18846 23650 18898 23662
rect 25118 23714 25170 23726
rect 25118 23650 25170 23662
rect 26014 23714 26066 23726
rect 26014 23650 26066 23662
rect 26126 23714 26178 23726
rect 29038 23714 29090 23726
rect 26898 23662 26910 23714
rect 26962 23662 26974 23714
rect 26126 23650 26178 23662
rect 29038 23650 29090 23662
rect 33742 23714 33794 23726
rect 33742 23650 33794 23662
rect 33966 23714 34018 23726
rect 33966 23650 34018 23662
rect 34414 23714 34466 23726
rect 34414 23650 34466 23662
rect 34750 23714 34802 23726
rect 34750 23650 34802 23662
rect 36318 23714 36370 23726
rect 38222 23714 38274 23726
rect 49534 23714 49586 23726
rect 37874 23662 37886 23714
rect 37938 23662 37950 23714
rect 41570 23662 41582 23714
rect 41634 23662 41646 23714
rect 42130 23662 42142 23714
rect 42194 23662 42206 23714
rect 36318 23650 36370 23662
rect 38222 23650 38274 23662
rect 16830 23602 16882 23614
rect 16830 23538 16882 23550
rect 22542 23602 22594 23614
rect 22542 23538 22594 23550
rect 23438 23602 23490 23614
rect 23438 23538 23490 23550
rect 24110 23602 24162 23614
rect 24110 23538 24162 23550
rect 27806 23602 27858 23614
rect 45714 23606 45726 23658
rect 45778 23606 45790 23658
rect 49534 23650 49586 23662
rect 51774 23714 51826 23726
rect 51774 23650 51826 23662
rect 55022 23714 55074 23726
rect 55022 23650 55074 23662
rect 27806 23538 27858 23550
rect 50430 23602 50482 23614
rect 56702 23602 56754 23614
rect 52546 23550 52558 23602
rect 52610 23550 52622 23602
rect 50430 23538 50482 23550
rect 56702 23538 56754 23550
rect 27682 23438 27694 23490
rect 27746 23487 27758 23490
rect 28466 23487 28478 23490
rect 27746 23441 28478 23487
rect 27746 23438 27758 23441
rect 28466 23438 28478 23441
rect 28530 23438 28542 23490
rect 39106 23438 39118 23490
rect 39170 23487 39182 23490
rect 39778 23487 39790 23490
rect 39170 23441 39790 23487
rect 39170 23438 39182 23441
rect 39778 23438 39790 23441
rect 39842 23487 39854 23490
rect 40226 23487 40238 23490
rect 39842 23441 40238 23487
rect 39842 23438 39854 23441
rect 40226 23438 40238 23441
rect 40290 23438 40302 23490
rect 1344 23210 58576 23244
rect 1344 23158 4478 23210
rect 4530 23158 4582 23210
rect 4634 23158 4686 23210
rect 4738 23158 35198 23210
rect 35250 23158 35302 23210
rect 35354 23158 35406 23210
rect 35458 23158 58576 23210
rect 1344 23124 58576 23158
rect 33618 22990 33630 23042
rect 33682 23039 33694 23042
rect 34402 23039 34414 23042
rect 33682 22993 34414 23039
rect 33682 22990 33694 22993
rect 34402 22990 34414 22993
rect 34466 22990 34478 23042
rect 35634 22990 35646 23042
rect 35698 23039 35710 23042
rect 35858 23039 35870 23042
rect 35698 22993 35870 23039
rect 35698 22990 35710 22993
rect 35858 22990 35870 22993
rect 35922 22990 35934 23042
rect 40338 22990 40350 23042
rect 40402 23039 40414 23042
rect 41234 23039 41246 23042
rect 40402 22993 41246 23039
rect 40402 22990 40414 22993
rect 41234 22990 41246 22993
rect 41298 22990 41310 23042
rect 4946 22878 4958 22930
rect 5010 22878 5022 22930
rect 28354 22878 28366 22930
rect 28418 22878 28430 22930
rect 36978 22878 36990 22930
rect 37042 22878 37054 22930
rect 37874 22878 37886 22930
rect 37938 22878 37950 22930
rect 41682 22878 41694 22930
rect 41746 22878 41758 22930
rect 5742 22818 5794 22830
rect 5742 22754 5794 22766
rect 6190 22818 6242 22830
rect 6190 22754 6242 22766
rect 20750 22818 20802 22830
rect 32958 22818 33010 22830
rect 25218 22766 25230 22818
rect 25282 22766 25294 22818
rect 20750 22754 20802 22766
rect 32958 22754 33010 22766
rect 34078 22818 34130 22830
rect 34078 22754 34130 22766
rect 39118 22818 39170 22830
rect 39118 22754 39170 22766
rect 39902 22818 39954 22830
rect 39902 22754 39954 22766
rect 40350 22818 40402 22830
rect 40350 22754 40402 22766
rect 40798 22818 40850 22830
rect 40798 22754 40850 22766
rect 41246 22818 41298 22830
rect 41246 22754 41298 22766
rect 41918 22818 41970 22830
rect 41918 22754 41970 22766
rect 42590 22818 42642 22830
rect 42590 22754 42642 22766
rect 43038 22818 43090 22830
rect 43038 22754 43090 22766
rect 43486 22818 43538 22830
rect 43486 22754 43538 22766
rect 44270 22818 44322 22830
rect 44270 22754 44322 22766
rect 49534 22818 49586 22830
rect 49534 22754 49586 22766
rect 49982 22818 50034 22830
rect 49982 22754 50034 22766
rect 51662 22818 51714 22830
rect 51662 22754 51714 22766
rect 52110 22818 52162 22830
rect 57698 22766 57710 22818
rect 57762 22766 57774 22818
rect 52110 22754 52162 22766
rect 1822 22706 1874 22718
rect 22318 22706 22370 22718
rect 2370 22654 2382 22706
rect 2434 22654 2446 22706
rect 1822 22642 1874 22654
rect 22318 22642 22370 22654
rect 24782 22706 24834 22718
rect 24782 22642 24834 22654
rect 25566 22706 25618 22718
rect 25566 22642 25618 22654
rect 25790 22706 25842 22718
rect 25790 22642 25842 22654
rect 35422 22706 35474 22718
rect 35422 22642 35474 22654
rect 35646 22706 35698 22718
rect 35646 22642 35698 22654
rect 35870 22706 35922 22718
rect 35870 22642 35922 22654
rect 36206 22706 36258 22718
rect 36206 22642 36258 22654
rect 37326 22706 37378 22718
rect 37326 22642 37378 22654
rect 37550 22706 37602 22718
rect 38446 22706 38498 22718
rect 38098 22654 38110 22706
rect 38162 22654 38174 22706
rect 37550 22642 37602 22654
rect 38446 22642 38498 22654
rect 41582 22706 41634 22718
rect 41582 22642 41634 22654
rect 42142 22706 42194 22718
rect 42142 22642 42194 22654
rect 53006 22706 53058 22718
rect 53006 22642 53058 22654
rect 53678 22706 53730 22718
rect 53678 22642 53730 22654
rect 54238 22706 54290 22718
rect 54238 22642 54290 22654
rect 57598 22706 57650 22718
rect 57598 22642 57650 22654
rect 15710 22594 15762 22606
rect 15710 22530 15762 22542
rect 16270 22594 16322 22606
rect 16270 22530 16322 22542
rect 16382 22594 16434 22606
rect 16382 22530 16434 22542
rect 16942 22594 16994 22606
rect 16942 22530 16994 22542
rect 21310 22594 21362 22606
rect 21310 22530 21362 22542
rect 21646 22594 21698 22606
rect 21646 22530 21698 22542
rect 21982 22594 22034 22606
rect 23438 22594 23490 22606
rect 22754 22542 22766 22594
rect 22818 22542 22830 22594
rect 21982 22530 22034 22542
rect 23438 22530 23490 22542
rect 25230 22594 25282 22606
rect 25230 22530 25282 22542
rect 26014 22594 26066 22606
rect 26014 22530 26066 22542
rect 27694 22594 27746 22606
rect 27694 22530 27746 22542
rect 33294 22594 33346 22606
rect 33294 22530 33346 22542
rect 35086 22594 35138 22606
rect 35086 22530 35138 22542
rect 36094 22594 36146 22606
rect 36094 22530 36146 22542
rect 36318 22594 36370 22606
rect 36318 22530 36370 22542
rect 52670 22594 52722 22606
rect 52670 22530 52722 22542
rect 53342 22594 53394 22606
rect 53342 22530 53394 22542
rect 54798 22594 54850 22606
rect 54798 22530 54850 22542
rect 20302 22482 20354 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 20302 22418 20354 22430
rect 24110 22482 24162 22494
rect 24110 22418 24162 22430
rect 24894 22482 24946 22494
rect 24894 22418 24946 22430
rect 32510 22482 32562 22494
rect 32510 22418 32562 22430
rect 33630 22482 33682 22494
rect 33630 22418 33682 22430
rect 34526 22482 34578 22494
rect 34526 22418 34578 22430
rect 44942 22482 44994 22494
rect 44942 22418 44994 22430
rect 50430 22482 50482 22494
rect 50430 22418 50482 22430
rect 51214 22482 51266 22494
rect 51214 22418 51266 22430
rect 55470 22482 55522 22494
rect 56466 22430 56478 22482
rect 56530 22430 56542 22482
rect 55470 22418 55522 22430
rect 15250 22318 15262 22370
rect 15314 22318 15326 22370
rect 1344 22202 58576 22236
rect 1344 22150 19838 22202
rect 19890 22150 19942 22202
rect 19994 22150 20046 22202
rect 20098 22150 50558 22202
rect 50610 22150 50662 22202
rect 50714 22150 50766 22202
rect 50818 22150 58576 22202
rect 1344 22116 58576 22150
rect 22642 21982 22654 22034
rect 22706 22031 22718 22034
rect 23426 22031 23438 22034
rect 22706 21985 23438 22031
rect 22706 21982 22718 21985
rect 23426 21982 23438 21985
rect 23490 21982 23502 22034
rect 39442 21982 39454 22034
rect 39506 22031 39518 22034
rect 39890 22031 39902 22034
rect 39506 21985 39902 22031
rect 39506 21982 39518 21985
rect 39890 21982 39902 21985
rect 39954 21982 39966 22034
rect 18286 21922 18338 21934
rect 15810 21870 15822 21922
rect 15874 21870 15886 21922
rect 18286 21858 18338 21870
rect 20526 21922 20578 21934
rect 20526 21858 20578 21870
rect 22094 21922 22146 21934
rect 22094 21858 22146 21870
rect 33630 21922 33682 21934
rect 38670 21922 38722 21934
rect 36642 21870 36654 21922
rect 36706 21870 36718 21922
rect 33630 21858 33682 21870
rect 38670 21858 38722 21870
rect 39454 21922 39506 21934
rect 39454 21858 39506 21870
rect 41022 21922 41074 21934
rect 41022 21858 41074 21870
rect 49758 21922 49810 21934
rect 49758 21858 49810 21870
rect 50206 21922 50258 21934
rect 50206 21858 50258 21870
rect 52894 21922 52946 21934
rect 52894 21858 52946 21870
rect 1822 21810 1874 21822
rect 1822 21746 1874 21758
rect 2270 21810 2322 21822
rect 2270 21746 2322 21758
rect 17838 21810 17890 21822
rect 17838 21746 17890 21758
rect 18622 21810 18674 21822
rect 18622 21746 18674 21758
rect 22766 21810 22818 21822
rect 22766 21746 22818 21758
rect 23214 21810 23266 21822
rect 23214 21746 23266 21758
rect 23886 21810 23938 21822
rect 23886 21746 23938 21758
rect 25118 21810 25170 21822
rect 25118 21746 25170 21758
rect 26014 21810 26066 21822
rect 26014 21746 26066 21758
rect 29150 21810 29202 21822
rect 29150 21746 29202 21758
rect 30046 21810 30098 21822
rect 30046 21746 30098 21758
rect 34750 21810 34802 21822
rect 37886 21810 37938 21822
rect 35970 21758 35982 21810
rect 36034 21758 36046 21810
rect 34750 21746 34802 21758
rect 37886 21746 37938 21758
rect 39902 21810 39954 21822
rect 39902 21746 39954 21758
rect 40350 21810 40402 21822
rect 40350 21746 40402 21758
rect 45838 21810 45890 21822
rect 45838 21746 45890 21758
rect 48862 21810 48914 21822
rect 48862 21746 48914 21758
rect 50654 21810 50706 21822
rect 50654 21746 50706 21758
rect 50766 21810 50818 21822
rect 50766 21746 50818 21758
rect 53566 21810 53618 21822
rect 53566 21746 53618 21758
rect 54014 21810 54066 21822
rect 54014 21746 54066 21758
rect 56702 21810 56754 21822
rect 56702 21746 56754 21758
rect 16830 21698 16882 21710
rect 25566 21698 25618 21710
rect 16370 21646 16382 21698
rect 16434 21646 16446 21698
rect 21186 21646 21198 21698
rect 21250 21646 21262 21698
rect 16830 21634 16882 21646
rect 25566 21634 25618 21646
rect 29598 21698 29650 21710
rect 41806 21698 41858 21710
rect 35186 21646 35198 21698
rect 35250 21646 35262 21698
rect 38770 21646 38782 21698
rect 38834 21646 38846 21698
rect 29598 21634 29650 21646
rect 24222 21586 24274 21598
rect 24222 21522 24274 21534
rect 24670 21586 24722 21598
rect 24670 21522 24722 21534
rect 26238 21586 26290 21598
rect 26238 21522 26290 21534
rect 26798 21586 26850 21598
rect 26798 21522 26850 21534
rect 28926 21586 28978 21598
rect 28926 21522 28978 21534
rect 30382 21586 30434 21598
rect 30382 21522 30434 21534
rect 32062 21586 32114 21598
rect 32062 21522 32114 21534
rect 32510 21586 32562 21598
rect 32510 21522 32562 21534
rect 33182 21586 33234 21598
rect 36194 21590 36206 21642
rect 36258 21590 36270 21642
rect 41806 21634 41858 21646
rect 43038 21698 43090 21710
rect 43038 21634 43090 21646
rect 43374 21698 43426 21710
rect 43374 21634 43426 21646
rect 43710 21698 43762 21710
rect 43710 21634 43762 21646
rect 44046 21698 44098 21710
rect 44046 21634 44098 21646
rect 44606 21698 44658 21710
rect 44606 21634 44658 21646
rect 45166 21698 45218 21710
rect 45166 21634 45218 21646
rect 47742 21698 47794 21710
rect 47742 21634 47794 21646
rect 50990 21698 51042 21710
rect 50990 21634 51042 21646
rect 54574 21698 54626 21710
rect 54574 21634 54626 21646
rect 55470 21698 55522 21710
rect 55682 21646 55694 21698
rect 55746 21646 55758 21698
rect 55470 21634 55522 21646
rect 33182 21522 33234 21534
rect 38334 21586 38386 21598
rect 38334 21522 38386 21534
rect 41582 21586 41634 21598
rect 41582 21522 41634 21534
rect 42254 21586 42306 21598
rect 42254 21522 42306 21534
rect 42702 21586 42754 21598
rect 42702 21522 42754 21534
rect 48190 21586 48242 21598
rect 48190 21522 48242 21534
rect 49310 21586 49362 21598
rect 57150 21586 57202 21598
rect 54338 21534 54350 21586
rect 54402 21534 54414 21586
rect 49310 21522 49362 21534
rect 57150 21522 57202 21534
rect 41470 21474 41522 21486
rect 41470 21410 41522 21422
rect 37762 21310 37774 21362
rect 37826 21359 37838 21362
rect 38322 21359 38334 21362
rect 37826 21313 38334 21359
rect 37826 21310 37838 21313
rect 38322 21310 38334 21313
rect 38386 21310 38398 21362
rect 55122 21310 55134 21362
rect 55186 21310 55198 21362
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 25442 20974 25454 21026
rect 25506 20974 25518 21026
rect 29698 20974 29710 21026
rect 29762 20974 29774 21026
rect 39106 20974 39118 21026
rect 39170 21023 39182 21026
rect 39442 21023 39454 21026
rect 39170 20977 39454 21023
rect 39170 20974 39182 20977
rect 39442 20974 39454 20977
rect 39506 20974 39518 21026
rect 43026 20974 43038 21026
rect 43090 20974 43102 21026
rect 50082 20974 50094 21026
rect 50146 20974 50158 21026
rect 56466 20974 56478 21026
rect 56530 20974 56542 21026
rect 24558 20914 24610 20926
rect 40686 20914 40738 20926
rect 24770 20862 24782 20914
rect 24834 20911 24846 20914
rect 24994 20911 25006 20914
rect 24834 20865 25006 20911
rect 24834 20862 24846 20865
rect 24994 20862 25006 20865
rect 25058 20862 25070 20914
rect 45490 20862 45502 20914
rect 45554 20911 45566 20914
rect 45554 20865 46111 20911
rect 45554 20862 45566 20865
rect 24558 20850 24610 20862
rect 40686 20850 40738 20862
rect 19182 20802 19234 20814
rect 16930 20750 16942 20802
rect 16994 20750 17006 20802
rect 19182 20738 19234 20750
rect 19854 20802 19906 20814
rect 19854 20738 19906 20750
rect 20302 20802 20354 20814
rect 20302 20738 20354 20750
rect 20750 20802 20802 20814
rect 20750 20738 20802 20750
rect 25006 20802 25058 20814
rect 25006 20738 25058 20750
rect 26350 20802 26402 20814
rect 26350 20738 26402 20750
rect 28590 20802 28642 20814
rect 28590 20738 28642 20750
rect 34638 20802 34690 20814
rect 34638 20738 34690 20750
rect 35086 20802 35138 20814
rect 35086 20738 35138 20750
rect 35534 20802 35586 20814
rect 35534 20738 35586 20750
rect 35982 20802 36034 20814
rect 35982 20738 36034 20750
rect 41134 20802 41186 20814
rect 41134 20738 41186 20750
rect 45502 20802 45554 20814
rect 45502 20738 45554 20750
rect 45950 20802 46002 20814
rect 46065 20799 46111 20865
rect 47630 20802 47682 20814
rect 46722 20799 46734 20802
rect 46065 20753 46734 20799
rect 46722 20750 46734 20753
rect 46786 20750 46798 20802
rect 45950 20738 46002 20750
rect 47630 20738 47682 20750
rect 51438 20802 51490 20814
rect 51438 20738 51490 20750
rect 51886 20802 51938 20814
rect 51886 20738 51938 20750
rect 56814 20802 56866 20814
rect 56814 20738 56866 20750
rect 57262 20802 57314 20814
rect 57262 20738 57314 20750
rect 21422 20690 21474 20702
rect 14690 20638 14702 20690
rect 14754 20638 14766 20690
rect 21422 20626 21474 20638
rect 23662 20690 23714 20702
rect 36430 20690 36482 20702
rect 29138 20638 29150 20690
rect 29202 20638 29214 20690
rect 23662 20626 23714 20638
rect 36430 20626 36482 20638
rect 37774 20690 37826 20702
rect 25342 20578 25394 20590
rect 21634 20526 21646 20578
rect 21698 20526 21710 20578
rect 25342 20514 25394 20526
rect 33406 20578 33458 20590
rect 37650 20582 37662 20634
rect 37714 20582 37726 20634
rect 37774 20626 37826 20638
rect 38222 20690 38274 20702
rect 38222 20626 38274 20638
rect 38558 20690 38610 20702
rect 38558 20626 38610 20638
rect 39118 20690 39170 20702
rect 39118 20626 39170 20638
rect 40350 20690 40402 20702
rect 45054 20690 45106 20702
rect 46734 20690 46786 20702
rect 43698 20638 43710 20690
rect 43762 20638 43774 20690
rect 46498 20638 46510 20690
rect 46562 20638 46574 20690
rect 40350 20626 40402 20638
rect 45054 20626 45106 20638
rect 46734 20626 46786 20638
rect 48302 20690 48354 20702
rect 55358 20690 55410 20702
rect 52882 20638 52894 20690
rect 52946 20638 52958 20690
rect 54338 20638 54350 20690
rect 54402 20638 54414 20690
rect 55906 20638 55918 20690
rect 55970 20638 55982 20690
rect 48302 20626 48354 20638
rect 55358 20626 55410 20638
rect 33406 20514 33458 20526
rect 39230 20578 39282 20590
rect 39230 20514 39282 20526
rect 40014 20578 40066 20590
rect 40014 20514 40066 20526
rect 41582 20578 41634 20590
rect 41582 20514 41634 20526
rect 43486 20578 43538 20590
rect 43486 20514 43538 20526
rect 44046 20578 44098 20590
rect 44046 20514 44098 20526
rect 46174 20578 46226 20590
rect 50094 20578 50146 20590
rect 48402 20526 48414 20578
rect 48466 20526 48478 20578
rect 53554 20526 53566 20578
rect 53618 20526 53630 20578
rect 46174 20514 46226 20526
rect 50094 20514 50146 20526
rect 25902 20466 25954 20478
rect 25902 20402 25954 20414
rect 33070 20466 33122 20478
rect 33070 20402 33122 20414
rect 34190 20466 34242 20478
rect 42814 20466 42866 20478
rect 37314 20414 37326 20466
rect 37378 20414 37390 20466
rect 34190 20402 34242 20414
rect 42814 20402 42866 20414
rect 54126 20466 54178 20478
rect 54126 20402 54178 20414
rect 54798 20466 54850 20478
rect 54798 20402 54850 20414
rect 47170 20302 47182 20354
rect 47234 20302 47246 20354
rect 1344 20186 58576 20220
rect 1344 20134 19838 20186
rect 19890 20134 19942 20186
rect 19994 20134 20046 20186
rect 20098 20134 50558 20186
rect 50610 20134 50662 20186
rect 50714 20134 50766 20186
rect 50818 20134 58576 20186
rect 1344 20100 58576 20134
rect 25778 19966 25790 20018
rect 25842 19966 25854 20018
rect 31378 19966 31390 20018
rect 31442 19966 31454 20018
rect 16718 19906 16770 19918
rect 16718 19842 16770 19854
rect 23998 19906 24050 19918
rect 23998 19842 24050 19854
rect 25566 19906 25618 19918
rect 25566 19842 25618 19854
rect 27470 19906 27522 19918
rect 27470 19842 27522 19854
rect 34526 19906 34578 19918
rect 45502 19906 45554 19918
rect 38210 19854 38222 19906
rect 38274 19854 38286 19906
rect 34526 19842 34578 19854
rect 45502 19842 45554 19854
rect 49758 19906 49810 19918
rect 49758 19842 49810 19854
rect 55470 19906 55522 19918
rect 55470 19842 55522 19854
rect 17726 19794 17778 19806
rect 17726 19730 17778 19742
rect 18174 19794 18226 19806
rect 18174 19730 18226 19742
rect 19630 19794 19682 19806
rect 19630 19730 19682 19742
rect 26798 19794 26850 19806
rect 26798 19730 26850 19742
rect 33854 19794 33906 19806
rect 33854 19730 33906 19742
rect 34190 19794 34242 19806
rect 34190 19730 34242 19742
rect 36206 19794 36258 19806
rect 36206 19730 36258 19742
rect 38782 19794 38834 19806
rect 38782 19730 38834 19742
rect 40350 19794 40402 19806
rect 40350 19730 40402 19742
rect 49086 19794 49138 19806
rect 51550 19794 51602 19806
rect 50194 19742 50206 19794
rect 50258 19742 50270 19794
rect 49086 19730 49138 19742
rect 51550 19730 51602 19742
rect 53342 19794 53394 19806
rect 54798 19794 54850 19806
rect 54114 19742 54126 19794
rect 54178 19742 54190 19794
rect 53342 19730 53394 19742
rect 54798 19730 54850 19742
rect 18958 19682 19010 19694
rect 16818 19630 16830 19682
rect 16882 19630 16894 19682
rect 17938 19630 17950 19682
rect 18002 19630 18014 19682
rect 18958 19618 19010 19630
rect 19294 19682 19346 19694
rect 19294 19618 19346 19630
rect 23214 19682 23266 19694
rect 23214 19618 23266 19630
rect 26238 19682 26290 19694
rect 31726 19682 31778 19694
rect 28354 19630 28366 19682
rect 28418 19630 28430 19682
rect 26238 19618 26290 19630
rect 31726 19618 31778 19630
rect 36094 19682 36146 19694
rect 36094 19618 36146 19630
rect 36654 19682 36706 19694
rect 36654 19618 36706 19630
rect 37774 19682 37826 19694
rect 37774 19618 37826 19630
rect 40910 19682 40962 19694
rect 40910 19618 40962 19630
rect 41022 19682 41074 19694
rect 41022 19618 41074 19630
rect 41470 19682 41522 19694
rect 41470 19618 41522 19630
rect 42030 19682 42082 19694
rect 42030 19618 42082 19630
rect 44494 19682 44546 19694
rect 44494 19618 44546 19630
rect 46174 19682 46226 19694
rect 46174 19618 46226 19630
rect 46398 19682 46450 19694
rect 46398 19618 46450 19630
rect 48750 19682 48802 19694
rect 48750 19618 48802 19630
rect 49422 19682 49474 19694
rect 49422 19618 49474 19630
rect 50878 19682 50930 19694
rect 50878 19618 50930 19630
rect 52670 19682 52722 19694
rect 52670 19618 52722 19630
rect 53006 19682 53058 19694
rect 53006 19618 53058 19630
rect 53678 19682 53730 19694
rect 53678 19618 53730 19630
rect 20190 19570 20242 19582
rect 26910 19570 26962 19582
rect 32174 19570 32226 19582
rect 22754 19518 22766 19570
rect 22818 19518 22830 19570
rect 29474 19518 29486 19570
rect 29538 19518 29550 19570
rect 20190 19506 20242 19518
rect 26910 19506 26962 19518
rect 32174 19506 32226 19518
rect 33182 19570 33234 19582
rect 33182 19506 33234 19518
rect 47518 19570 47570 19582
rect 47518 19506 47570 19518
rect 52334 19570 52386 19582
rect 52334 19506 52386 19518
rect 56702 19570 56754 19582
rect 56702 19506 56754 19518
rect 33518 19458 33570 19470
rect 33518 19394 33570 19406
rect 40014 19458 40066 19470
rect 40014 19394 40066 19406
rect 18610 19294 18622 19346
rect 18674 19294 18686 19346
rect 27010 19294 27022 19346
rect 27074 19343 27086 19346
rect 27346 19343 27358 19346
rect 27074 19297 27358 19343
rect 27074 19294 27086 19297
rect 27346 19294 27358 19297
rect 27410 19294 27422 19346
rect 45714 19294 45726 19346
rect 45778 19343 45790 19346
rect 46162 19343 46174 19346
rect 45778 19297 46174 19343
rect 45778 19294 45790 19297
rect 46162 19294 46174 19297
rect 46226 19294 46238 19346
rect 1344 19178 58576 19212
rect 1344 19126 4478 19178
rect 4530 19126 4582 19178
rect 4634 19126 4686 19178
rect 4738 19126 35198 19178
rect 35250 19126 35302 19178
rect 35354 19126 35406 19178
rect 35458 19126 58576 19178
rect 1344 19092 58576 19126
rect 31602 18958 31614 19010
rect 31666 19007 31678 19010
rect 32050 19007 32062 19010
rect 31666 18961 32062 19007
rect 31666 18958 31678 18961
rect 32050 18958 32062 18961
rect 32114 18958 32126 19010
rect 41010 18958 41022 19010
rect 41074 18958 41086 19010
rect 51426 18958 51438 19010
rect 51490 19007 51502 19010
rect 52210 19007 52222 19010
rect 51490 18961 52222 19007
rect 51490 18958 51502 18961
rect 52210 18958 52222 18961
rect 52274 18958 52286 19010
rect 35410 18846 35422 18898
rect 35474 18895 35486 18898
rect 35970 18895 35982 18898
rect 35474 18849 35982 18895
rect 35474 18846 35486 18849
rect 35970 18846 35982 18849
rect 36034 18846 36046 18898
rect 50978 18846 50990 18898
rect 51042 18895 51054 18898
rect 51874 18895 51886 18898
rect 51042 18849 51886 18895
rect 51042 18846 51054 18849
rect 51874 18846 51886 18849
rect 51938 18846 51950 18898
rect 54786 18846 54798 18898
rect 54850 18846 54862 18898
rect 20750 18786 20802 18798
rect 17826 18734 17838 18786
rect 17890 18734 17902 18786
rect 20750 18722 20802 18734
rect 25566 18786 25618 18798
rect 25566 18722 25618 18734
rect 26462 18786 26514 18798
rect 26462 18722 26514 18734
rect 27358 18786 27410 18798
rect 27358 18722 27410 18734
rect 30158 18786 30210 18798
rect 30158 18722 30210 18734
rect 30942 18786 30994 18798
rect 30942 18722 30994 18734
rect 31726 18786 31778 18798
rect 34526 18786 34578 18798
rect 33170 18734 33182 18786
rect 33234 18734 33246 18786
rect 31726 18722 31778 18734
rect 34526 18722 34578 18734
rect 35422 18786 35474 18798
rect 35422 18722 35474 18734
rect 35870 18786 35922 18798
rect 35870 18722 35922 18734
rect 37102 18786 37154 18798
rect 37102 18722 37154 18734
rect 38670 18786 38722 18798
rect 38670 18722 38722 18734
rect 39118 18786 39170 18798
rect 46062 18786 46114 18798
rect 43586 18734 43598 18786
rect 43650 18734 43662 18786
rect 39118 18722 39170 18734
rect 46062 18722 46114 18734
rect 51438 18786 51490 18798
rect 54674 18734 54686 18786
rect 54738 18734 54750 18786
rect 51438 18722 51490 18734
rect 24222 18674 24274 18686
rect 15138 18622 15150 18674
rect 15202 18622 15214 18674
rect 24222 18610 24274 18622
rect 25006 18674 25058 18686
rect 25006 18610 25058 18622
rect 30494 18674 30546 18686
rect 30494 18610 30546 18622
rect 32062 18674 32114 18686
rect 32062 18610 32114 18622
rect 34974 18674 35026 18686
rect 34974 18610 35026 18622
rect 46958 18674 47010 18686
rect 46958 18610 47010 18622
rect 47630 18674 47682 18686
rect 47630 18610 47682 18622
rect 47966 18674 48018 18686
rect 52882 18678 52894 18730
rect 52946 18678 52958 18730
rect 47966 18610 48018 18622
rect 57150 18674 57202 18686
rect 57150 18610 57202 18622
rect 26014 18562 26066 18574
rect 26014 18498 26066 18510
rect 28590 18562 28642 18574
rect 28590 18498 28642 18510
rect 34078 18562 34130 18574
rect 34078 18498 34130 18510
rect 36318 18562 36370 18574
rect 36318 18498 36370 18510
rect 39454 18562 39506 18574
rect 39454 18498 39506 18510
rect 40126 18562 40178 18574
rect 40126 18498 40178 18510
rect 45614 18562 45666 18574
rect 45614 18498 45666 18510
rect 47294 18562 47346 18574
rect 47294 18498 47346 18510
rect 48526 18562 48578 18574
rect 48526 18498 48578 18510
rect 49086 18562 49138 18574
rect 49086 18498 49138 18510
rect 49758 18562 49810 18574
rect 49758 18498 49810 18510
rect 50542 18562 50594 18574
rect 50542 18498 50594 18510
rect 53230 18562 53282 18574
rect 53230 18498 53282 18510
rect 55134 18562 55186 18574
rect 57698 18510 57710 18562
rect 57762 18510 57774 18562
rect 55134 18498 55186 18510
rect 39790 18450 39842 18462
rect 22642 18398 22654 18450
rect 22706 18398 22718 18450
rect 39790 18386 39842 18398
rect 41358 18450 41410 18462
rect 41358 18386 41410 18398
rect 50990 18450 51042 18462
rect 50990 18386 51042 18398
rect 51886 18450 51938 18462
rect 51886 18386 51938 18398
rect 51202 18286 51214 18338
rect 51266 18335 51278 18338
rect 51874 18335 51886 18338
rect 51266 18289 51886 18335
rect 51266 18286 51278 18289
rect 51874 18286 51886 18289
rect 51938 18286 51950 18338
rect 1344 18170 58576 18204
rect 1344 18118 19838 18170
rect 19890 18118 19942 18170
rect 19994 18118 20046 18170
rect 20098 18118 50558 18170
rect 50610 18118 50662 18170
rect 50714 18118 50766 18170
rect 50818 18118 58576 18170
rect 1344 18084 58576 18118
rect 23874 17950 23886 18002
rect 23938 17999 23950 18002
rect 24210 17999 24222 18002
rect 23938 17953 24222 17999
rect 23938 17950 23950 17953
rect 24210 17950 24222 17953
rect 24274 17999 24286 18002
rect 24658 17999 24670 18002
rect 24274 17953 24670 17999
rect 24274 17950 24286 17953
rect 24658 17950 24670 17953
rect 24722 17950 24734 18002
rect 30594 17950 30606 18002
rect 30658 17999 30670 18002
rect 31602 17999 31614 18002
rect 30658 17953 31614 17999
rect 30658 17950 30670 17953
rect 31602 17950 31614 17953
rect 31666 17950 31678 18002
rect 49074 17950 49086 18002
rect 49138 17950 49150 18002
rect 16830 17890 16882 17902
rect 24222 17890 24274 17902
rect 22642 17838 22654 17890
rect 22706 17838 22718 17890
rect 16830 17826 16882 17838
rect 24222 17826 24274 17838
rect 24670 17890 24722 17902
rect 24670 17826 24722 17838
rect 27806 17890 27858 17902
rect 27806 17826 27858 17838
rect 30606 17890 30658 17902
rect 30606 17826 30658 17838
rect 31054 17890 31106 17902
rect 31054 17826 31106 17838
rect 31502 17890 31554 17902
rect 31502 17826 31554 17838
rect 39454 17890 39506 17902
rect 39454 17826 39506 17838
rect 39902 17890 39954 17902
rect 39902 17826 39954 17838
rect 41022 17890 41074 17902
rect 41022 17826 41074 17838
rect 41470 17890 41522 17902
rect 41470 17826 41522 17838
rect 46062 17890 46114 17902
rect 46062 17826 46114 17838
rect 48302 17890 48354 17902
rect 48302 17826 48354 17838
rect 51662 17890 51714 17902
rect 51662 17826 51714 17838
rect 53678 17890 53730 17902
rect 53678 17826 53730 17838
rect 25342 17778 25394 17790
rect 25342 17714 25394 17726
rect 27134 17778 27186 17790
rect 27134 17714 27186 17726
rect 28366 17778 28418 17790
rect 28366 17714 28418 17726
rect 29598 17778 29650 17790
rect 29598 17714 29650 17726
rect 33182 17778 33234 17790
rect 33182 17714 33234 17726
rect 35982 17778 36034 17790
rect 35982 17714 36034 17726
rect 42254 17778 42306 17790
rect 42254 17714 42306 17726
rect 43374 17778 43426 17790
rect 43374 17714 43426 17726
rect 52670 17778 52722 17790
rect 52670 17714 52722 17726
rect 53342 17778 53394 17790
rect 53342 17714 53394 17726
rect 54798 17778 54850 17790
rect 54798 17714 54850 17726
rect 55470 17778 55522 17790
rect 55470 17714 55522 17726
rect 17726 17666 17778 17678
rect 17726 17602 17778 17614
rect 26798 17666 26850 17678
rect 26798 17602 26850 17614
rect 27470 17666 27522 17678
rect 27470 17602 27522 17614
rect 28926 17666 28978 17678
rect 28926 17602 28978 17614
rect 33518 17666 33570 17678
rect 33518 17602 33570 17614
rect 33854 17666 33906 17678
rect 33854 17602 33906 17614
rect 34190 17666 34242 17678
rect 34190 17602 34242 17614
rect 34750 17666 34802 17678
rect 34750 17602 34802 17614
rect 35310 17666 35362 17678
rect 35310 17602 35362 17614
rect 41918 17666 41970 17678
rect 41918 17602 41970 17614
rect 42702 17666 42754 17678
rect 42702 17602 42754 17614
rect 48974 17666 49026 17678
rect 48974 17602 49026 17614
rect 49310 17666 49362 17678
rect 49310 17602 49362 17614
rect 53006 17666 53058 17678
rect 53006 17602 53058 17614
rect 54238 17666 54290 17678
rect 54238 17602 54290 17614
rect 18734 17554 18786 17566
rect 18734 17490 18786 17502
rect 23662 17554 23714 17566
rect 32286 17554 32338 17566
rect 26450 17502 26462 17554
rect 26514 17502 26526 17554
rect 23662 17490 23714 17502
rect 32286 17490 32338 17502
rect 36766 17554 36818 17566
rect 36766 17490 36818 17502
rect 40350 17554 40402 17566
rect 40350 17490 40402 17502
rect 47294 17554 47346 17566
rect 47294 17490 47346 17502
rect 47742 17554 47794 17566
rect 47742 17490 47794 17502
rect 49870 17554 49922 17566
rect 49870 17490 49922 17502
rect 50766 17554 50818 17566
rect 50766 17490 50818 17502
rect 51214 17554 51266 17566
rect 51214 17490 51266 17502
rect 52334 17554 52386 17566
rect 52334 17490 52386 17502
rect 51090 17278 51102 17330
rect 51154 17327 51166 17330
rect 51650 17327 51662 17330
rect 51154 17281 51662 17327
rect 51154 17278 51166 17281
rect 51650 17278 51662 17281
rect 51714 17278 51726 17330
rect 1344 17162 58576 17196
rect 1344 17110 4478 17162
rect 4530 17110 4582 17162
rect 4634 17110 4686 17162
rect 4738 17110 35198 17162
rect 35250 17110 35302 17162
rect 35354 17110 35406 17162
rect 35458 17110 58576 17162
rect 1344 17076 58576 17110
rect 55682 16942 55694 16994
rect 55746 16942 55758 16994
rect 35522 16830 35534 16882
rect 35586 16830 35598 16882
rect 20302 16770 20354 16782
rect 20302 16706 20354 16718
rect 22094 16770 22146 16782
rect 22094 16706 22146 16718
rect 22542 16770 22594 16782
rect 22542 16706 22594 16718
rect 22990 16770 23042 16782
rect 22990 16706 23042 16718
rect 23886 16770 23938 16782
rect 23886 16706 23938 16718
rect 28478 16770 28530 16782
rect 28478 16706 28530 16718
rect 45726 16770 45778 16782
rect 45726 16706 45778 16718
rect 50990 16770 51042 16782
rect 50990 16706 51042 16718
rect 24222 16658 24274 16670
rect 24782 16658 24834 16670
rect 24434 16606 24446 16658
rect 24498 16606 24510 16658
rect 24222 16594 24274 16606
rect 24782 16594 24834 16606
rect 25342 16658 25394 16670
rect 30046 16658 30098 16670
rect 45054 16658 45106 16670
rect 29250 16606 29262 16658
rect 29314 16606 29326 16658
rect 32050 16606 32062 16658
rect 32114 16606 32126 16658
rect 25342 16594 25394 16606
rect 30046 16594 30098 16606
rect 45054 16594 45106 16606
rect 45390 16658 45442 16670
rect 53678 16658 53730 16670
rect 53218 16606 53230 16658
rect 53282 16606 53294 16658
rect 45390 16594 45442 16606
rect 53678 16594 53730 16606
rect 54126 16658 54178 16670
rect 54126 16594 54178 16606
rect 54574 16658 54626 16670
rect 54574 16594 54626 16606
rect 54910 16658 54962 16670
rect 54910 16594 54962 16606
rect 55134 16658 55186 16670
rect 55134 16594 55186 16606
rect 55358 16658 55410 16670
rect 55358 16594 55410 16606
rect 55582 16658 55634 16670
rect 55582 16594 55634 16606
rect 56142 16658 56194 16670
rect 56142 16594 56194 16606
rect 23438 16546 23490 16558
rect 23438 16482 23490 16494
rect 27806 16546 27858 16558
rect 27806 16482 27858 16494
rect 30830 16546 30882 16558
rect 30830 16482 30882 16494
rect 31054 16546 31106 16558
rect 31054 16482 31106 16494
rect 31502 16546 31554 16558
rect 31502 16482 31554 16494
rect 34414 16546 34466 16558
rect 34414 16482 34466 16494
rect 39678 16546 39730 16558
rect 39678 16482 39730 16494
rect 40014 16546 40066 16558
rect 40014 16482 40066 16494
rect 40350 16546 40402 16558
rect 41806 16546 41858 16558
rect 41122 16494 41134 16546
rect 41186 16494 41198 16546
rect 40350 16482 40402 16494
rect 41806 16482 41858 16494
rect 46958 16546 47010 16558
rect 46958 16482 47010 16494
rect 56590 16546 56642 16558
rect 56590 16482 56642 16494
rect 40686 16434 40738 16446
rect 40686 16370 40738 16382
rect 42478 16434 42530 16446
rect 42478 16370 42530 16382
rect 47294 16434 47346 16446
rect 47294 16370 47346 16382
rect 48414 16434 48466 16446
rect 48414 16370 48466 16382
rect 48862 16434 48914 16446
rect 48862 16370 48914 16382
rect 49646 16434 49698 16446
rect 49646 16370 49698 16382
rect 50094 16434 50146 16446
rect 50094 16370 50146 16382
rect 50542 16434 50594 16446
rect 50542 16370 50594 16382
rect 51438 16434 51490 16446
rect 51438 16370 51490 16382
rect 52110 16434 52162 16446
rect 57038 16434 57090 16446
rect 53442 16382 53454 16434
rect 53506 16382 53518 16434
rect 52110 16370 52162 16382
rect 57038 16370 57090 16382
rect 57486 16434 57538 16446
rect 57486 16370 57538 16382
rect 30370 16270 30382 16322
rect 30434 16270 30446 16322
rect 1344 16154 58576 16188
rect 1344 16102 19838 16154
rect 19890 16102 19942 16154
rect 19994 16102 20046 16154
rect 20098 16102 50558 16154
rect 50610 16102 50662 16154
rect 50714 16102 50766 16154
rect 50818 16102 58576 16154
rect 1344 16068 58576 16102
rect 28018 15934 28030 15986
rect 28082 15934 28094 15986
rect 31266 15934 31278 15986
rect 31330 15934 31342 15986
rect 51090 15934 51102 15986
rect 51154 15983 51166 15986
rect 51426 15983 51438 15986
rect 51154 15937 51438 15983
rect 51154 15934 51166 15937
rect 51426 15934 51438 15937
rect 51490 15983 51502 15986
rect 51762 15983 51774 15986
rect 51490 15937 51774 15983
rect 51490 15934 51502 15937
rect 51762 15934 51774 15937
rect 51826 15934 51838 15986
rect 23214 15874 23266 15886
rect 23214 15810 23266 15822
rect 23662 15874 23714 15886
rect 23662 15810 23714 15822
rect 24110 15874 24162 15886
rect 24110 15810 24162 15822
rect 37102 15874 37154 15886
rect 37102 15810 37154 15822
rect 39230 15874 39282 15886
rect 39230 15810 39282 15822
rect 40238 15874 40290 15886
rect 40238 15810 40290 15822
rect 41246 15874 41298 15886
rect 41246 15810 41298 15822
rect 42142 15874 42194 15886
rect 42142 15810 42194 15822
rect 49198 15874 49250 15886
rect 49198 15810 49250 15822
rect 49534 15874 49586 15886
rect 49534 15810 49586 15822
rect 50094 15874 50146 15886
rect 50094 15810 50146 15822
rect 50990 15874 51042 15886
rect 50990 15810 51042 15822
rect 51438 15874 51490 15886
rect 51438 15810 51490 15822
rect 52334 15874 52386 15886
rect 52334 15810 52386 15822
rect 53678 15874 53730 15886
rect 53678 15810 53730 15822
rect 19742 15762 19794 15774
rect 19742 15698 19794 15710
rect 24670 15762 24722 15774
rect 24670 15698 24722 15710
rect 25230 15762 25282 15774
rect 25230 15698 25282 15710
rect 29710 15762 29762 15774
rect 29710 15698 29762 15710
rect 32174 15762 32226 15774
rect 32174 15698 32226 15710
rect 37550 15762 37602 15774
rect 37550 15698 37602 15710
rect 38558 15762 38610 15774
rect 38558 15698 38610 15710
rect 48190 15762 48242 15774
rect 48190 15698 48242 15710
rect 53006 15762 53058 15774
rect 53006 15698 53058 15710
rect 53342 15762 53394 15774
rect 53342 15698 53394 15710
rect 54238 15762 54290 15774
rect 54238 15698 54290 15710
rect 55470 15762 55522 15774
rect 55470 15698 55522 15710
rect 17726 15650 17778 15662
rect 17726 15586 17778 15598
rect 30494 15650 30546 15662
rect 30494 15586 30546 15598
rect 31726 15650 31778 15662
rect 31726 15586 31778 15598
rect 32958 15650 33010 15662
rect 32958 15586 33010 15598
rect 33182 15650 33234 15662
rect 33182 15586 33234 15598
rect 33742 15650 33794 15662
rect 33742 15586 33794 15598
rect 34190 15650 34242 15662
rect 34190 15586 34242 15598
rect 36654 15650 36706 15662
rect 36654 15586 36706 15598
rect 37998 15650 38050 15662
rect 49646 15650 49698 15662
rect 48962 15598 48974 15650
rect 49026 15598 49038 15650
rect 37998 15586 38050 15598
rect 49646 15586 49698 15598
rect 52670 15650 52722 15662
rect 52670 15586 52722 15598
rect 54798 15650 54850 15662
rect 54798 15586 54850 15598
rect 32398 15538 32450 15550
rect 28914 15486 28926 15538
rect 28978 15486 28990 15538
rect 32398 15474 32450 15486
rect 38670 15538 38722 15550
rect 38670 15474 38722 15486
rect 41694 15538 41746 15550
rect 41694 15474 41746 15486
rect 47294 15538 47346 15550
rect 47294 15474 47346 15486
rect 47742 15538 47794 15550
rect 47742 15474 47794 15486
rect 50542 15538 50594 15550
rect 50542 15474 50594 15486
rect 51886 15538 51938 15550
rect 51886 15474 51938 15486
rect 48638 15426 48690 15438
rect 20178 15374 20190 15426
rect 20242 15374 20254 15426
rect 48638 15362 48690 15374
rect 1344 15146 58576 15180
rect 1344 15094 4478 15146
rect 4530 15094 4582 15146
rect 4634 15094 4686 15146
rect 4738 15094 35198 15146
rect 35250 15094 35302 15146
rect 35354 15094 35406 15146
rect 35458 15094 58576 15146
rect 1344 15060 58576 15094
rect 33842 14926 33854 14978
rect 33906 14926 33918 14978
rect 42254 14866 42306 14878
rect 19282 14814 19294 14866
rect 19346 14863 19358 14866
rect 20178 14863 20190 14866
rect 19346 14817 20190 14863
rect 19346 14814 19358 14817
rect 20178 14814 20190 14817
rect 20242 14814 20254 14866
rect 29250 14814 29262 14866
rect 29314 14863 29326 14866
rect 29810 14863 29822 14866
rect 29314 14817 29822 14863
rect 29314 14814 29326 14817
rect 29810 14814 29822 14817
rect 29874 14863 29886 14866
rect 30146 14863 30158 14866
rect 29874 14817 30158 14863
rect 29874 14814 29886 14817
rect 30146 14814 30158 14817
rect 30210 14814 30222 14866
rect 42254 14802 42306 14814
rect 19182 14754 19234 14766
rect 19182 14690 19234 14702
rect 27134 14754 27186 14766
rect 27134 14690 27186 14702
rect 29262 14754 29314 14766
rect 29262 14690 29314 14702
rect 30158 14754 30210 14766
rect 30158 14690 30210 14702
rect 35982 14754 36034 14766
rect 35982 14690 36034 14702
rect 36430 14754 36482 14766
rect 36430 14690 36482 14702
rect 37326 14754 37378 14766
rect 37326 14690 37378 14702
rect 51774 14754 51826 14766
rect 56242 14702 56254 14754
rect 56306 14702 56318 14754
rect 51774 14690 51826 14702
rect 19630 14642 19682 14654
rect 19630 14578 19682 14590
rect 23886 14642 23938 14654
rect 23886 14578 23938 14590
rect 25006 14642 25058 14654
rect 35086 14642 35138 14654
rect 27570 14590 27582 14642
rect 27634 14590 27646 14642
rect 25006 14578 25058 14590
rect 35086 14578 35138 14590
rect 37774 14642 37826 14654
rect 37774 14578 37826 14590
rect 37886 14642 37938 14654
rect 37886 14578 37938 14590
rect 38222 14642 38274 14654
rect 38222 14578 38274 14590
rect 39006 14642 39058 14654
rect 39006 14578 39058 14590
rect 43822 14642 43874 14654
rect 48638 14642 48690 14654
rect 44930 14590 44942 14642
rect 44994 14590 45006 14642
rect 43822 14578 43874 14590
rect 48638 14578 48690 14590
rect 48974 14642 49026 14654
rect 48974 14578 49026 14590
rect 49310 14642 49362 14654
rect 49310 14578 49362 14590
rect 49870 14642 49922 14654
rect 49870 14578 49922 14590
rect 52894 14642 52946 14654
rect 57026 14590 57038 14642
rect 57090 14590 57102 14642
rect 52894 14578 52946 14590
rect 20078 14530 20130 14542
rect 20078 14466 20130 14478
rect 21422 14530 21474 14542
rect 21422 14466 21474 14478
rect 22206 14530 22258 14542
rect 22206 14466 22258 14478
rect 22878 14530 22930 14542
rect 22878 14466 22930 14478
rect 23214 14530 23266 14542
rect 23214 14466 23266 14478
rect 23550 14530 23602 14542
rect 23550 14466 23602 14478
rect 24446 14530 24498 14542
rect 24446 14466 24498 14478
rect 26686 14530 26738 14542
rect 26686 14466 26738 14478
rect 28254 14530 28306 14542
rect 28254 14466 28306 14478
rect 31278 14530 31330 14542
rect 31278 14466 31330 14478
rect 41246 14530 41298 14542
rect 41246 14466 41298 14478
rect 44270 14530 44322 14542
rect 44270 14466 44322 14478
rect 45502 14530 45554 14542
rect 45502 14466 45554 14478
rect 47854 14530 47906 14542
rect 47854 14466 47906 14478
rect 48302 14530 48354 14542
rect 48302 14466 48354 14478
rect 50430 14530 50482 14542
rect 50430 14466 50482 14478
rect 51102 14530 51154 14542
rect 51102 14466 51154 14478
rect 52670 14530 52722 14542
rect 52670 14466 52722 14478
rect 54462 14530 54514 14542
rect 54898 14478 54910 14530
rect 54962 14478 54974 14530
rect 56130 14478 56142 14530
rect 56194 14478 56206 14530
rect 54462 14466 54514 14478
rect 21870 14418 21922 14430
rect 21870 14354 21922 14366
rect 22542 14418 22594 14430
rect 22542 14354 22594 14366
rect 25678 14418 25730 14430
rect 25678 14354 25730 14366
rect 28702 14418 28754 14430
rect 28702 14354 28754 14366
rect 29710 14418 29762 14430
rect 29710 14354 29762 14366
rect 30942 14418 30994 14430
rect 30942 14354 30994 14366
rect 35534 14418 35586 14430
rect 35534 14354 35586 14366
rect 19842 14254 19854 14306
rect 19906 14303 19918 14306
rect 20066 14303 20078 14306
rect 19906 14257 20078 14303
rect 19906 14254 19918 14257
rect 20066 14254 20078 14257
rect 20130 14254 20142 14306
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 54786 13918 54798 13970
rect 54850 13918 54862 13970
rect 19182 13858 19234 13870
rect 19182 13794 19234 13806
rect 24446 13858 24498 13870
rect 24446 13794 24498 13806
rect 25342 13858 25394 13870
rect 25342 13794 25394 13806
rect 25790 13858 25842 13870
rect 25790 13794 25842 13806
rect 26686 13858 26738 13870
rect 26686 13794 26738 13806
rect 29150 13858 29202 13870
rect 29150 13794 29202 13806
rect 30942 13858 30994 13870
rect 30942 13794 30994 13806
rect 32062 13858 32114 13870
rect 32062 13794 32114 13806
rect 32510 13858 32562 13870
rect 32510 13794 32562 13806
rect 33294 13858 33346 13870
rect 33294 13794 33346 13806
rect 33630 13858 33682 13870
rect 33630 13794 33682 13806
rect 36318 13858 36370 13870
rect 36318 13794 36370 13806
rect 38110 13858 38162 13870
rect 38110 13794 38162 13806
rect 46062 13858 46114 13870
rect 56030 13858 56082 13870
rect 54562 13806 54574 13858
rect 54626 13806 54638 13858
rect 46062 13794 46114 13806
rect 56030 13794 56082 13806
rect 16830 13746 16882 13758
rect 20078 13746 20130 13758
rect 18395 13694 18407 13746
rect 18459 13694 18471 13746
rect 16830 13682 16882 13694
rect 20078 13682 20130 13694
rect 23326 13746 23378 13758
rect 23326 13682 23378 13694
rect 28590 13746 28642 13758
rect 28590 13682 28642 13694
rect 35646 13746 35698 13758
rect 41134 13746 41186 13758
rect 36754 13694 36766 13746
rect 36818 13694 36830 13746
rect 35646 13682 35698 13694
rect 41134 13682 41186 13694
rect 45390 13746 45442 13758
rect 45390 13682 45442 13694
rect 46622 13746 46674 13758
rect 46622 13682 46674 13694
rect 47182 13746 47234 13758
rect 47182 13682 47234 13694
rect 47854 13746 47906 13758
rect 54238 13746 54290 13758
rect 50530 13694 50542 13746
rect 50594 13694 50606 13746
rect 47854 13682 47906 13694
rect 54238 13682 54290 13694
rect 54910 13746 54962 13758
rect 54910 13682 54962 13694
rect 55022 13746 55074 13758
rect 55022 13682 55074 13694
rect 19742 13634 19794 13646
rect 20974 13634 21026 13646
rect 17490 13582 17502 13634
rect 17554 13582 17566 13634
rect 20402 13582 20414 13634
rect 20466 13582 20478 13634
rect 19742 13570 19794 13582
rect 20974 13570 21026 13582
rect 35310 13634 35362 13646
rect 35310 13570 35362 13582
rect 35982 13634 36034 13646
rect 35982 13570 36034 13582
rect 37438 13634 37490 13646
rect 37438 13570 37490 13582
rect 38894 13634 38946 13646
rect 43710 13634 43762 13646
rect 41682 13582 41694 13634
rect 41746 13582 41758 13634
rect 38894 13570 38946 13582
rect 43710 13570 43762 13582
rect 45054 13634 45106 13646
rect 45054 13570 45106 13582
rect 45726 13634 45778 13646
rect 52658 13582 52670 13634
rect 52722 13582 52734 13634
rect 45726 13570 45778 13582
rect 26238 13522 26290 13534
rect 44494 13522 44546 13534
rect 39778 13470 39790 13522
rect 39842 13470 39854 13522
rect 26238 13458 26290 13470
rect 44494 13458 44546 13470
rect 55582 13522 55634 13534
rect 55582 13458 55634 13470
rect 1344 13130 58576 13164
rect 1344 13078 4478 13130
rect 4530 13078 4582 13130
rect 4634 13078 4686 13130
rect 4738 13078 35198 13130
rect 35250 13078 35302 13130
rect 35354 13078 35406 13130
rect 35458 13078 58576 13130
rect 1344 13044 58576 13078
rect 42590 12850 42642 12862
rect 19282 12798 19294 12850
rect 19346 12798 19358 12850
rect 42590 12786 42642 12798
rect 55918 12850 55970 12862
rect 55918 12786 55970 12798
rect 22430 12738 22482 12750
rect 22430 12674 22482 12686
rect 27022 12738 27074 12750
rect 27022 12674 27074 12686
rect 33742 12738 33794 12750
rect 33742 12674 33794 12686
rect 48302 12738 48354 12750
rect 48302 12674 48354 12686
rect 50990 12738 51042 12750
rect 50990 12674 51042 12686
rect 51550 12738 51602 12750
rect 51550 12674 51602 12686
rect 51886 12738 51938 12750
rect 51886 12674 51938 12686
rect 52782 12738 52834 12750
rect 53890 12686 53902 12738
rect 53954 12686 53966 12738
rect 52782 12674 52834 12686
rect 17502 12626 17554 12638
rect 17502 12562 17554 12574
rect 23662 12626 23714 12638
rect 23662 12562 23714 12574
rect 24334 12626 24386 12638
rect 24334 12562 24386 12574
rect 24894 12626 24946 12638
rect 24894 12562 24946 12574
rect 30382 12626 30434 12638
rect 30382 12562 30434 12574
rect 31614 12626 31666 12638
rect 31614 12562 31666 12574
rect 39454 12626 39506 12638
rect 46722 12574 46734 12626
rect 46786 12574 46798 12626
rect 55346 12574 55358 12626
rect 55410 12574 55422 12626
rect 39454 12562 39506 12574
rect 18958 12514 19010 12526
rect 18958 12450 19010 12462
rect 21310 12514 21362 12526
rect 21310 12450 21362 12462
rect 23326 12514 23378 12526
rect 23326 12450 23378 12462
rect 23998 12514 24050 12526
rect 23998 12450 24050 12462
rect 25454 12514 25506 12526
rect 25454 12450 25506 12462
rect 30046 12514 30098 12526
rect 30046 12450 30098 12462
rect 30718 12514 30770 12526
rect 30718 12450 30770 12462
rect 32174 12514 32226 12526
rect 32174 12450 32226 12462
rect 38446 12514 38498 12526
rect 38446 12450 38498 12462
rect 38558 12514 38610 12526
rect 38558 12450 38610 12462
rect 39230 12514 39282 12526
rect 39230 12450 39282 12462
rect 53678 12514 53730 12526
rect 53678 12450 53730 12462
rect 26126 12402 26178 12414
rect 26126 12338 26178 12350
rect 31054 12402 31106 12414
rect 31054 12338 31106 12350
rect 32846 12402 32898 12414
rect 32846 12338 32898 12350
rect 35534 12402 35586 12414
rect 35534 12338 35586 12350
rect 35982 12402 36034 12414
rect 35982 12338 36034 12350
rect 36430 12402 36482 12414
rect 36430 12338 36482 12350
rect 37326 12402 37378 12414
rect 37326 12338 37378 12350
rect 37774 12402 37826 12414
rect 37774 12338 37826 12350
rect 38222 12402 38274 12414
rect 38222 12338 38274 12350
rect 46398 12402 46450 12414
rect 46398 12338 46450 12350
rect 1344 12122 58576 12156
rect 1344 12070 19838 12122
rect 19890 12070 19942 12122
rect 19994 12070 20046 12122
rect 20098 12070 50558 12122
rect 50610 12070 50662 12122
rect 50714 12070 50766 12122
rect 50818 12070 58576 12122
rect 1344 12036 58576 12070
rect 22754 11902 22766 11954
rect 22818 11951 22830 11954
rect 23314 11951 23326 11954
rect 22818 11905 23326 11951
rect 22818 11902 22830 11905
rect 23314 11902 23326 11905
rect 23378 11902 23390 11954
rect 31042 11902 31054 11954
rect 31106 11951 31118 11954
rect 31714 11951 31726 11954
rect 31106 11905 31726 11951
rect 31106 11902 31118 11905
rect 31714 11902 31726 11905
rect 31778 11902 31790 11954
rect 30606 11842 30658 11854
rect 30606 11778 30658 11790
rect 52782 11842 52834 11854
rect 52782 11778 52834 11790
rect 53790 11842 53842 11854
rect 53790 11778 53842 11790
rect 20526 11730 20578 11742
rect 20526 11666 20578 11678
rect 25902 11730 25954 11742
rect 31166 11730 31218 11742
rect 29474 11678 29486 11730
rect 29538 11678 29550 11730
rect 25902 11666 25954 11678
rect 31166 11666 31218 11678
rect 36766 11730 36818 11742
rect 36766 11666 36818 11678
rect 37662 11730 37714 11742
rect 37662 11666 37714 11678
rect 40462 11730 40514 11742
rect 48862 11730 48914 11742
rect 42354 11678 42366 11730
rect 42418 11678 42430 11730
rect 44370 11678 44382 11730
rect 44434 11678 44446 11730
rect 40462 11666 40514 11678
rect 48862 11666 48914 11678
rect 53342 11730 53394 11742
rect 53342 11666 53394 11678
rect 19742 11618 19794 11630
rect 19742 11554 19794 11566
rect 22542 11618 22594 11630
rect 22542 11554 22594 11566
rect 25454 11618 25506 11630
rect 25454 11554 25506 11566
rect 26350 11618 26402 11630
rect 26350 11554 26402 11566
rect 26798 11618 26850 11630
rect 26798 11554 26850 11566
rect 27134 11618 27186 11630
rect 33630 11618 33682 11630
rect 29810 11566 29822 11618
rect 29874 11566 29886 11618
rect 27134 11554 27186 11566
rect 33630 11554 33682 11566
rect 36318 11618 36370 11630
rect 36318 11554 36370 11566
rect 41470 11618 41522 11630
rect 41470 11554 41522 11566
rect 42030 11618 42082 11630
rect 42030 11554 42082 11566
rect 52334 11618 52386 11630
rect 52334 11554 52386 11566
rect 19406 11506 19458 11518
rect 19406 11442 19458 11454
rect 22990 11506 23042 11518
rect 22990 11442 23042 11454
rect 23438 11506 23490 11518
rect 23438 11442 23490 11454
rect 24670 11506 24722 11518
rect 24670 11442 24722 11454
rect 31614 11506 31666 11518
rect 31614 11442 31666 11454
rect 32062 11506 32114 11518
rect 32062 11442 32114 11454
rect 32510 11506 32562 11518
rect 32510 11442 32562 11454
rect 33070 11506 33122 11518
rect 33070 11442 33122 11454
rect 35870 11506 35922 11518
rect 35870 11442 35922 11454
rect 37326 11506 37378 11518
rect 37326 11442 37378 11454
rect 41022 11506 41074 11518
rect 45602 11454 45614 11506
rect 45666 11454 45678 11506
rect 41022 11442 41074 11454
rect 31602 11230 31614 11282
rect 31666 11279 31678 11282
rect 32386 11279 32398 11282
rect 31666 11233 32398 11279
rect 31666 11230 31678 11233
rect 32386 11230 32398 11233
rect 32450 11230 32462 11282
rect 1344 11114 58576 11148
rect 1344 11062 4478 11114
rect 4530 11062 4582 11114
rect 4634 11062 4686 11114
rect 4738 11062 35198 11114
rect 35250 11062 35302 11114
rect 35354 11062 35406 11114
rect 35458 11062 58576 11114
rect 1344 11028 58576 11062
rect 20290 10894 20302 10946
rect 20354 10943 20366 10946
rect 20738 10943 20750 10946
rect 20354 10897 20750 10943
rect 20354 10894 20366 10897
rect 20738 10894 20750 10897
rect 20802 10894 20814 10946
rect 36978 10894 36990 10946
rect 37042 10894 37054 10946
rect 25118 10834 25170 10846
rect 47854 10834 47906 10846
rect 35298 10782 35310 10834
rect 35362 10782 35374 10834
rect 25118 10770 25170 10782
rect 47854 10770 47906 10782
rect 20302 10722 20354 10734
rect 20302 10658 20354 10670
rect 21422 10722 21474 10734
rect 21422 10658 21474 10670
rect 30382 10722 30434 10734
rect 30382 10658 30434 10670
rect 30830 10722 30882 10734
rect 30830 10658 30882 10670
rect 31278 10722 31330 10734
rect 31278 10658 31330 10670
rect 35982 10722 36034 10734
rect 35982 10658 36034 10670
rect 36430 10722 36482 10734
rect 36430 10658 36482 10670
rect 41582 10722 41634 10734
rect 41582 10658 41634 10670
rect 42030 10722 42082 10734
rect 42030 10658 42082 10670
rect 43598 10722 43650 10734
rect 43598 10658 43650 10670
rect 53118 10722 53170 10734
rect 53118 10658 53170 10670
rect 31614 10610 31666 10622
rect 31614 10546 31666 10558
rect 34190 10610 34242 10622
rect 34190 10546 34242 10558
rect 37774 10610 37826 10622
rect 37774 10546 37826 10558
rect 38894 10610 38946 10622
rect 38894 10546 38946 10558
rect 39118 10610 39170 10622
rect 39118 10546 39170 10558
rect 41134 10610 41186 10622
rect 41134 10546 41186 10558
rect 44046 10610 44098 10622
rect 44046 10546 44098 10558
rect 45166 10610 45218 10622
rect 45166 10546 45218 10558
rect 45390 10610 45442 10622
rect 45390 10546 45442 10558
rect 45502 10610 45554 10622
rect 45502 10546 45554 10558
rect 20750 10498 20802 10510
rect 20750 10434 20802 10446
rect 21870 10498 21922 10510
rect 24446 10498 24498 10510
rect 22306 10446 22318 10498
rect 22370 10446 22382 10498
rect 21870 10434 21922 10446
rect 24446 10434 24498 10446
rect 32398 10498 32450 10510
rect 38658 10446 38670 10498
rect 38722 10446 38734 10498
rect 32398 10434 32450 10446
rect 25790 10386 25842 10398
rect 25790 10322 25842 10334
rect 1344 10106 58576 10140
rect 1344 10054 19838 10106
rect 19890 10054 19942 10106
rect 19994 10054 20046 10106
rect 20098 10054 50558 10106
rect 50610 10054 50662 10106
rect 50714 10054 50766 10106
rect 50818 10054 58576 10106
rect 1344 10020 58576 10054
rect 23650 9886 23662 9938
rect 23714 9935 23726 9938
rect 24658 9935 24670 9938
rect 23714 9889 24670 9935
rect 23714 9886 23726 9889
rect 24658 9886 24670 9889
rect 24722 9886 24734 9938
rect 30146 9886 30158 9938
rect 30210 9886 30222 9938
rect 33506 9886 33518 9938
rect 33570 9935 33582 9938
rect 34514 9935 34526 9938
rect 33570 9889 34526 9935
rect 33570 9886 33582 9889
rect 34514 9886 34526 9889
rect 34578 9886 34590 9938
rect 18174 9826 18226 9838
rect 23662 9826 23714 9838
rect 22866 9774 22878 9826
rect 22930 9774 22942 9826
rect 18174 9762 18226 9774
rect 23662 9762 23714 9774
rect 24222 9826 24274 9838
rect 24222 9762 24274 9774
rect 25678 9826 25730 9838
rect 25678 9762 25730 9774
rect 33518 9826 33570 9838
rect 33518 9762 33570 9774
rect 33966 9826 34018 9838
rect 33966 9762 34018 9774
rect 44494 9826 44546 9838
rect 44494 9762 44546 9774
rect 24670 9714 24722 9726
rect 21298 9662 21310 9714
rect 21362 9662 21374 9714
rect 24670 9650 24722 9662
rect 18622 9602 18674 9614
rect 18622 9538 18674 9550
rect 19070 9602 19122 9614
rect 26014 9602 26066 9614
rect 21634 9550 21646 9602
rect 21698 9550 21710 9602
rect 19070 9538 19122 9550
rect 26014 9538 26066 9550
rect 26574 9602 26626 9614
rect 26574 9538 26626 9550
rect 28814 9602 28866 9614
rect 28814 9538 28866 9550
rect 34526 9602 34578 9614
rect 34526 9538 34578 9550
rect 35198 9602 35250 9614
rect 35198 9538 35250 9550
rect 37538 9438 37550 9490
rect 37602 9438 37614 9490
rect 1344 9098 58576 9132
rect 1344 9046 4478 9098
rect 4530 9046 4582 9098
rect 4634 9046 4686 9098
rect 4738 9046 35198 9098
rect 35250 9046 35302 9098
rect 35354 9046 35406 9098
rect 35458 9046 58576 9098
rect 1344 9012 58576 9046
rect 26226 8878 26238 8930
rect 26290 8878 26302 8930
rect 32174 8818 32226 8830
rect 21634 8766 21646 8818
rect 21698 8815 21710 8818
rect 22978 8815 22990 8818
rect 21698 8769 22990 8815
rect 21698 8766 21710 8769
rect 22978 8766 22990 8769
rect 23042 8766 23054 8818
rect 32174 8754 32226 8766
rect 21646 8706 21698 8718
rect 21646 8642 21698 8654
rect 22094 8706 22146 8718
rect 22094 8642 22146 8654
rect 22542 8706 22594 8718
rect 22542 8642 22594 8654
rect 22990 8706 23042 8718
rect 22990 8642 23042 8654
rect 28142 8706 28194 8718
rect 28142 8642 28194 8654
rect 36430 8706 36482 8718
rect 36430 8642 36482 8654
rect 37102 8706 37154 8718
rect 37102 8642 37154 8654
rect 23662 8594 23714 8606
rect 23662 8530 23714 8542
rect 23774 8594 23826 8606
rect 23774 8530 23826 8542
rect 24894 8594 24946 8606
rect 24894 8530 24946 8542
rect 28590 8594 28642 8606
rect 28590 8530 28642 8542
rect 29262 8594 29314 8606
rect 29262 8530 29314 8542
rect 29598 8594 29650 8606
rect 29598 8530 29650 8542
rect 27694 8482 27746 8494
rect 23986 8430 23998 8482
rect 24050 8430 24062 8482
rect 27694 8418 27746 8430
rect 31726 8370 31778 8382
rect 31726 8306 31778 8318
rect 1344 8090 58576 8124
rect 1344 8038 19838 8090
rect 19890 8038 19942 8090
rect 19994 8038 20046 8090
rect 20098 8038 50558 8090
rect 50610 8038 50662 8090
rect 50714 8038 50766 8090
rect 50818 8038 58576 8090
rect 1344 8004 58576 8038
rect 3838 7810 3890 7822
rect 3838 7746 3890 7758
rect 4286 7810 4338 7822
rect 4286 7746 4338 7758
rect 22318 7810 22370 7822
rect 22318 7746 22370 7758
rect 22766 7810 22818 7822
rect 22766 7746 22818 7758
rect 28254 7810 28306 7822
rect 28254 7746 28306 7758
rect 28702 7810 28754 7822
rect 28702 7746 28754 7758
rect 29598 7810 29650 7822
rect 29598 7746 29650 7758
rect 32286 7810 32338 7822
rect 32286 7746 32338 7758
rect 29150 7698 29202 7710
rect 29150 7634 29202 7646
rect 30606 7698 30658 7710
rect 30606 7634 30658 7646
rect 31614 7698 31666 7710
rect 31614 7634 31666 7646
rect 30270 7586 30322 7598
rect 30270 7522 30322 7534
rect 30382 7586 30434 7598
rect 30382 7522 30434 7534
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 1344 6074 58576 6108
rect 1344 6022 19838 6074
rect 19890 6022 19942 6074
rect 19994 6022 20046 6074
rect 20098 6022 50558 6074
rect 50610 6022 50662 6074
rect 50714 6022 50766 6074
rect 50818 6022 58576 6074
rect 1344 5988 58576 6022
rect 1344 5066 58576 5100
rect 1344 5014 4478 5066
rect 4530 5014 4582 5066
rect 4634 5014 4686 5066
rect 4738 5014 35198 5066
rect 35250 5014 35302 5066
rect 35354 5014 35406 5066
rect 35458 5014 58576 5066
rect 1344 4980 58576 5014
rect 1344 4058 58576 4092
rect 1344 4006 19838 4058
rect 19890 4006 19942 4058
rect 19994 4006 20046 4058
rect 20098 4006 50558 4058
rect 50610 4006 50662 4058
rect 50714 4006 50766 4058
rect 50818 4006 58576 4058
rect 1344 3972 58576 4006
<< via1 >>
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4478 55414 4530 55466
rect 4582 55414 4634 55466
rect 4686 55414 4738 55466
rect 35198 55414 35250 55466
rect 35302 55414 35354 55466
rect 35406 55414 35458 55466
rect 19838 54406 19890 54458
rect 19942 54406 19994 54458
rect 20046 54406 20098 54458
rect 50558 54406 50610 54458
rect 50662 54406 50714 54458
rect 50766 54406 50818 54458
rect 3838 54126 3890 54178
rect 56030 54126 56082 54178
rect 4478 53398 4530 53450
rect 4582 53398 4634 53450
rect 4686 53398 4738 53450
rect 35198 53398 35250 53450
rect 35302 53398 35354 53450
rect 35406 53398 35458 53450
rect 19838 52390 19890 52442
rect 19942 52390 19994 52442
rect 20046 52390 20098 52442
rect 50558 52390 50610 52442
rect 50662 52390 50714 52442
rect 50766 52390 50818 52442
rect 4478 51382 4530 51434
rect 4582 51382 4634 51434
rect 4686 51382 4738 51434
rect 35198 51382 35250 51434
rect 35302 51382 35354 51434
rect 35406 51382 35458 51434
rect 19838 50374 19890 50426
rect 19942 50374 19994 50426
rect 20046 50374 20098 50426
rect 50558 50374 50610 50426
rect 50662 50374 50714 50426
rect 50766 50374 50818 50426
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 32062 49086 32114 49138
rect 33518 49086 33570 49138
rect 32062 48974 32114 49026
rect 39230 48862 39282 48914
rect 39566 48862 39618 48914
rect 21422 48750 21474 48802
rect 23662 48750 23714 48802
rect 23998 48750 24050 48802
rect 24334 48750 24386 48802
rect 25230 48750 25282 48802
rect 25790 48750 25842 48802
rect 32510 48750 32562 48802
rect 33070 48750 33122 48802
rect 33518 48750 33570 48802
rect 38782 48750 38834 48802
rect 40686 48750 40738 48802
rect 41358 48750 41410 48802
rect 42590 48750 42642 48802
rect 43150 48750 43202 48802
rect 21870 48638 21922 48690
rect 22318 48638 22370 48690
rect 24670 48638 24722 48690
rect 26462 48638 26514 48690
rect 35534 48638 35586 48690
rect 38334 48638 38386 48690
rect 41246 48638 41298 48690
rect 19838 48358 19890 48410
rect 19942 48358 19994 48410
rect 20046 48358 20098 48410
rect 50558 48358 50610 48410
rect 50662 48358 50714 48410
rect 50766 48358 50818 48410
rect 26462 48190 26514 48242
rect 27246 48190 27298 48242
rect 27694 48190 27746 48242
rect 23102 48078 23154 48130
rect 26462 48078 26514 48130
rect 35534 48078 35586 48130
rect 41470 48078 41522 48130
rect 19854 47966 19906 48018
rect 22094 47966 22146 48018
rect 26014 47966 26066 48018
rect 28478 47966 28530 48018
rect 19518 47854 19570 47906
rect 27694 47854 27746 47906
rect 36990 47854 37042 47906
rect 39006 47854 39058 47906
rect 19070 47742 19122 47794
rect 23550 47742 23602 47794
rect 23998 47742 24050 47794
rect 26910 47742 26962 47794
rect 27358 47742 27410 47794
rect 32062 47742 32114 47794
rect 32622 47742 32674 47794
rect 40350 47742 40402 47794
rect 41022 47742 41074 47794
rect 41918 47742 41970 47794
rect 42366 47742 42418 47794
rect 42814 47742 42866 47794
rect 43262 47742 43314 47794
rect 43822 47742 43874 47794
rect 44158 47742 44210 47794
rect 45166 47742 45218 47794
rect 50206 47742 50258 47794
rect 50654 47742 50706 47794
rect 52110 47742 52162 47794
rect 52670 47742 52722 47794
rect 53006 47742 53058 47794
rect 53454 47742 53506 47794
rect 31054 47630 31106 47682
rect 41022 47630 41074 47682
rect 41582 47630 41634 47682
rect 42366 47630 42418 47682
rect 43150 47630 43202 47682
rect 52110 47630 52162 47682
rect 53006 47630 53058 47682
rect 27022 47518 27074 47570
rect 27358 47518 27410 47570
rect 40798 47518 40850 47570
rect 41358 47518 41410 47570
rect 41918 47518 41970 47570
rect 42814 47518 42866 47570
rect 4478 47350 4530 47402
rect 4582 47350 4634 47402
rect 4686 47350 4738 47402
rect 35198 47350 35250 47402
rect 35302 47350 35354 47402
rect 35406 47350 35458 47402
rect 27246 47070 27298 47122
rect 27806 47070 27858 47122
rect 28478 47070 28530 47122
rect 21646 46958 21698 47010
rect 25902 46958 25954 47010
rect 27246 46958 27298 47010
rect 28142 46958 28194 47010
rect 28590 46958 28642 47010
rect 43150 46958 43202 47010
rect 43598 46958 43650 47010
rect 22430 46846 22482 46898
rect 22878 46846 22930 46898
rect 29374 46846 29426 46898
rect 29822 46846 29874 46898
rect 32174 46846 32226 46898
rect 32622 46846 32674 46898
rect 34078 46846 34130 46898
rect 34862 46846 34914 46898
rect 37550 46846 37602 46898
rect 41246 46846 41298 46898
rect 45502 46846 45554 46898
rect 52782 46846 52834 46898
rect 53678 46846 53730 46898
rect 17838 46734 17890 46786
rect 39118 46734 39170 46786
rect 39454 46734 39506 46786
rect 39790 46734 39842 46786
rect 40686 46734 40738 46786
rect 17390 46622 17442 46674
rect 18510 46622 18562 46674
rect 20526 46622 20578 46674
rect 22094 46622 22146 46674
rect 25118 46622 25170 46674
rect 27694 46622 27746 46674
rect 33182 46622 33234 46674
rect 33854 46622 33906 46674
rect 37102 46622 37154 46674
rect 37998 46622 38050 46674
rect 40126 46622 40178 46674
rect 41918 46622 41970 46674
rect 42702 46622 42754 46674
rect 44046 46622 44098 46674
rect 44942 46622 44994 46674
rect 53230 46622 53282 46674
rect 54126 46622 54178 46674
rect 21646 46510 21698 46562
rect 22094 46510 22146 46562
rect 22430 46510 22482 46562
rect 35646 46510 35698 46562
rect 43150 46510 43202 46562
rect 43934 46510 43986 46562
rect 50990 46510 51042 46562
rect 53230 46510 53282 46562
rect 53790 46510 53842 46562
rect 19838 46342 19890 46394
rect 19942 46342 19994 46394
rect 20046 46342 20098 46394
rect 50558 46342 50610 46394
rect 50662 46342 50714 46394
rect 50766 46342 50818 46394
rect 32286 46174 32338 46226
rect 41918 46174 41970 46226
rect 22654 46062 22706 46114
rect 23326 46062 23378 46114
rect 24222 46062 24274 46114
rect 25454 46062 25506 46114
rect 26462 46062 26514 46114
rect 27246 46062 27298 46114
rect 30606 46062 30658 46114
rect 35870 46062 35922 46114
rect 39566 46062 39618 46114
rect 46174 46062 46226 46114
rect 25230 45950 25282 46002
rect 28254 45950 28306 46002
rect 31950 45950 32002 46002
rect 33070 45950 33122 46002
rect 34526 45950 34578 46002
rect 35198 45950 35250 46002
rect 40126 45950 40178 46002
rect 41134 45950 41186 46002
rect 44046 45950 44098 46002
rect 50878 45950 50930 46002
rect 51550 45950 51602 46002
rect 53006 45950 53058 46002
rect 53790 45950 53842 46002
rect 54910 45950 54962 46002
rect 55358 45950 55410 46002
rect 17950 45838 18002 45890
rect 18286 45838 18338 45890
rect 20526 45838 20578 45890
rect 27806 45838 27858 45890
rect 31502 45838 31554 45890
rect 33406 45838 33458 45890
rect 33742 45838 33794 45890
rect 34078 45838 34130 45890
rect 37886 45838 37938 45890
rect 39118 45838 39170 45890
rect 41358 45838 41410 45890
rect 41582 45838 41634 45890
rect 41806 45838 41858 45890
rect 42814 45838 42866 45890
rect 43934 45838 43986 45890
rect 45278 45865 45330 45917
rect 48750 45838 48802 45890
rect 49086 45838 49138 45890
rect 49422 45838 49474 45890
rect 49758 45838 49810 45890
rect 50318 45838 50370 45890
rect 53454 45838 53506 45890
rect 54014 45838 54066 45890
rect 17502 45726 17554 45778
rect 21758 45726 21810 45778
rect 23774 45726 23826 45778
rect 24670 45726 24722 45778
rect 36990 45726 37042 45778
rect 37550 45726 37602 45778
rect 46622 45726 46674 45778
rect 47070 45726 47122 45778
rect 48190 45726 48242 45778
rect 52334 45726 52386 45778
rect 53678 45726 53730 45778
rect 23774 45614 23826 45666
rect 24670 45614 24722 45666
rect 43822 45614 43874 45666
rect 4478 45334 4530 45386
rect 4582 45334 4634 45386
rect 4686 45334 4738 45386
rect 35198 45334 35250 45386
rect 35302 45334 35354 45386
rect 35406 45334 35458 45386
rect 38670 45166 38722 45218
rect 48526 45166 48578 45218
rect 35310 45054 35362 45106
rect 34078 44942 34130 44994
rect 37550 44942 37602 44994
rect 17166 44830 17218 44882
rect 17502 44830 17554 44882
rect 18062 44830 18114 44882
rect 24558 44830 24610 44882
rect 27358 44830 27410 44882
rect 32062 44830 32114 44882
rect 32622 44830 32674 44882
rect 34526 44830 34578 44882
rect 36094 44830 36146 44882
rect 37102 44830 37154 44882
rect 37886 44830 37938 44882
rect 38110 44830 38162 44882
rect 38334 44830 38386 44882
rect 39566 44830 39618 44882
rect 43710 44830 43762 44882
rect 44832 44830 44884 44882
rect 45278 44830 45330 44882
rect 46622 44830 46674 44882
rect 50990 44830 51042 44882
rect 53006 44830 53058 44882
rect 54798 44830 54850 44882
rect 21310 44718 21362 44770
rect 21870 44718 21922 44770
rect 28142 44718 28194 44770
rect 30494 44718 30546 44770
rect 30830 44718 30882 44770
rect 31166 44718 31218 44770
rect 39230 44718 39282 44770
rect 39902 44718 39954 44770
rect 40798 44718 40850 44770
rect 41358 44718 41410 44770
rect 43262 44718 43314 44770
rect 43486 44718 43538 44770
rect 43934 44718 43986 44770
rect 45054 44718 45106 44770
rect 50654 44718 50706 44770
rect 51214 44718 51266 44770
rect 51886 44718 51938 44770
rect 52670 44718 52722 44770
rect 53342 44718 53394 44770
rect 54126 44718 54178 44770
rect 20302 44606 20354 44658
rect 20638 44606 20690 44658
rect 24222 44606 24274 44658
rect 25342 44606 25394 44658
rect 26014 44606 26066 44658
rect 28254 44606 28306 44658
rect 31502 44606 31554 44658
rect 33294 44606 33346 44658
rect 40238 44606 40290 44658
rect 42030 44606 42082 44658
rect 43598 44606 43650 44658
rect 44942 44606 44994 44658
rect 51438 44606 51490 44658
rect 53678 44606 53730 44658
rect 55470 44606 55522 44658
rect 19838 44326 19890 44378
rect 19942 44326 19994 44378
rect 20046 44326 20098 44378
rect 50558 44326 50610 44378
rect 50662 44326 50714 44378
rect 50766 44326 50818 44378
rect 20302 44158 20354 44210
rect 21198 44158 21250 44210
rect 24222 44158 24274 44210
rect 24558 44158 24610 44210
rect 31278 44158 31330 44210
rect 38110 44158 38162 44210
rect 39006 44158 39058 44210
rect 40798 44158 40850 44210
rect 41358 44158 41410 44210
rect 20302 44046 20354 44098
rect 21198 44046 21250 44098
rect 21646 44046 21698 44098
rect 24222 44046 24274 44098
rect 24670 44046 24722 44098
rect 25678 44046 25730 44098
rect 27246 44046 27298 44098
rect 28702 44046 28754 44098
rect 30494 44046 30546 44098
rect 34190 44046 34242 44098
rect 39006 44046 39058 44098
rect 43486 44046 43538 44098
rect 45950 44046 46002 44098
rect 48078 44046 48130 44098
rect 55470 44046 55522 44098
rect 29038 43934 29090 43986
rect 32174 43934 32226 43986
rect 42142 43934 42194 43986
rect 42590 43934 42642 43986
rect 49646 43934 49698 43986
rect 51886 43934 51938 43986
rect 53118 43934 53170 43986
rect 54686 43934 54738 43986
rect 56702 43934 56754 43986
rect 57150 43934 57202 43986
rect 31726 43822 31778 43874
rect 38558 43822 38610 43874
rect 39454 43822 39506 43874
rect 44046 43822 44098 43874
rect 45166 43822 45218 43874
rect 46958 43822 47010 43874
rect 47294 43822 47346 43874
rect 47406 43822 47458 43874
rect 47630 43822 47682 43874
rect 50878 43822 50930 43874
rect 52894 43822 52946 43874
rect 55022 43822 55074 43874
rect 19854 43710 19906 43762
rect 20750 43710 20802 43762
rect 26126 43710 26178 43762
rect 28030 43710 28082 43762
rect 37326 43710 37378 43762
rect 37774 43710 37826 43762
rect 38110 43710 38162 43762
rect 39902 43710 39954 43762
rect 40350 43710 40402 43762
rect 41022 43710 41074 43762
rect 41470 43710 41522 43762
rect 42814 43710 42866 43762
rect 49534 43710 49586 43762
rect 38670 43598 38722 43650
rect 39118 43598 39170 43650
rect 39902 43598 39954 43650
rect 40350 43598 40402 43650
rect 20750 43486 20802 43538
rect 21646 43486 21698 43538
rect 41694 43486 41746 43538
rect 4478 43318 4530 43370
rect 4582 43318 4634 43370
rect 4686 43318 4738 43370
rect 35198 43318 35250 43370
rect 35302 43318 35354 43370
rect 35406 43318 35458 43370
rect 47294 43150 47346 43202
rect 48638 43150 48690 43202
rect 50654 43150 50706 43202
rect 51550 43150 51602 43202
rect 33966 43038 34018 43090
rect 37102 43038 37154 43090
rect 37550 43038 37602 43090
rect 38334 43038 38386 43090
rect 47742 43038 47794 43090
rect 49086 43038 49138 43090
rect 21646 42926 21698 42978
rect 27246 42926 27298 42978
rect 27694 42926 27746 42978
rect 37550 42926 37602 42978
rect 39790 42926 39842 42978
rect 42478 42926 42530 42978
rect 47294 42926 47346 42978
rect 47742 42926 47794 42978
rect 48638 42926 48690 42978
rect 49086 42926 49138 42978
rect 55134 42926 55186 42978
rect 7534 42814 7586 42866
rect 8094 42814 8146 42866
rect 23102 42814 23154 42866
rect 23438 42814 23490 42866
rect 23774 42814 23826 42866
rect 24670 42814 24722 42866
rect 25230 42814 25282 42866
rect 29038 42814 29090 42866
rect 30270 42814 30322 42866
rect 32958 42814 33010 42866
rect 33294 42814 33346 42866
rect 38670 42814 38722 42866
rect 39454 42814 39506 42866
rect 42590 42814 42642 42866
rect 42702 42814 42754 42866
rect 43598 42814 43650 42866
rect 43934 42814 43986 42866
rect 45390 42814 45442 42866
rect 46398 42814 46450 42866
rect 50206 42814 50258 42866
rect 53230 42814 53282 42866
rect 53454 42814 53506 42866
rect 53790 42814 53842 42866
rect 54348 42814 54400 42866
rect 55358 42814 55410 42866
rect 56142 42814 56194 42866
rect 56478 42814 56530 42866
rect 25902 42702 25954 42754
rect 28142 42702 28194 42754
rect 29374 42702 29426 42754
rect 29598 42702 29650 42754
rect 39230 42702 39282 42754
rect 40462 42702 40514 42754
rect 41246 42702 41298 42754
rect 45166 42702 45218 42754
rect 45614 42702 45666 42754
rect 54238 42702 54290 42754
rect 55694 42702 55746 42754
rect 56926 42702 56978 42754
rect 7198 42590 7250 42642
rect 10222 42590 10274 42642
rect 10670 42590 10722 42642
rect 20414 42590 20466 42642
rect 22094 42590 22146 42642
rect 24110 42590 24162 42642
rect 26798 42590 26850 42642
rect 28590 42590 28642 42642
rect 36430 42590 36482 42642
rect 37102 42590 37154 42642
rect 37998 42590 38050 42642
rect 41918 42590 41970 42642
rect 46846 42590 46898 42642
rect 48190 42590 48242 42642
rect 49758 42590 49810 42642
rect 50654 42590 50706 42642
rect 51102 42590 51154 42642
rect 51550 42590 51602 42642
rect 51998 42590 52050 42642
rect 53342 42590 53394 42642
rect 55806 42590 55858 42642
rect 57374 42590 57426 42642
rect 57822 42590 57874 42642
rect 37102 42478 37154 42530
rect 37998 42478 38050 42530
rect 44718 42478 44770 42530
rect 55022 42478 55074 42530
rect 56702 42478 56754 42530
rect 57822 42478 57874 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 6862 42030 6914 42082
rect 35086 42030 35138 42082
rect 44046 42030 44098 42082
rect 48974 42030 49026 42082
rect 50878 42030 50930 42082
rect 52670 42030 52722 42082
rect 56702 42030 56754 42082
rect 9662 41918 9714 41970
rect 9774 41918 9826 41970
rect 19294 41918 19346 41970
rect 19518 41918 19570 41970
rect 21646 41918 21698 41970
rect 22766 41918 22818 41970
rect 25342 41918 25394 41970
rect 27470 41918 27522 41970
rect 27918 41918 27970 41970
rect 30270 41918 30322 41970
rect 30830 41918 30882 41970
rect 34414 41918 34466 41970
rect 36878 41918 36930 41970
rect 39566 41918 39618 41970
rect 41918 41918 41970 41970
rect 42366 41918 42418 41970
rect 43038 41918 43090 41970
rect 43710 41918 43762 41970
rect 45166 41918 45218 41970
rect 45838 41918 45890 41970
rect 52222 41918 52274 41970
rect 53790 41918 53842 41970
rect 54798 41918 54850 41970
rect 55694 41918 55746 41970
rect 4062 41806 4114 41858
rect 4622 41806 4674 41858
rect 11006 41806 11058 41858
rect 25566 41806 25618 41858
rect 26798 41806 26850 41858
rect 33966 41806 34018 41858
rect 36318 41806 36370 41858
rect 36430 41806 36482 41858
rect 37774 41806 37826 41858
rect 39902 41806 39954 41858
rect 42142 41806 42194 41858
rect 43374 41806 43426 41858
rect 44606 41806 44658 41858
rect 46622 41806 46674 41858
rect 52334 41806 52386 41858
rect 56030 41806 56082 41858
rect 1822 41694 1874 41746
rect 3726 41694 3778 41746
rect 24670 41694 24722 41746
rect 28142 41694 28194 41746
rect 28814 41694 28866 41746
rect 30942 41694 30994 41746
rect 31502 41694 31554 41746
rect 33406 41694 33458 41746
rect 40350 41694 40402 41746
rect 41358 41694 41410 41746
rect 49422 41694 49474 41746
rect 49870 41694 49922 41746
rect 50430 41694 50482 41746
rect 51326 41694 51378 41746
rect 57150 41694 57202 41746
rect 57598 41694 57650 41746
rect 7198 41582 7250 41634
rect 23886 41582 23938 41634
rect 37214 41582 37266 41634
rect 49422 41582 49474 41634
rect 50430 41582 50482 41634
rect 55470 41582 55522 41634
rect 10894 41470 10946 41522
rect 21534 41470 21586 41522
rect 27022 41470 27074 41522
rect 29822 41470 29874 41522
rect 41470 41470 41522 41522
rect 49870 41470 49922 41522
rect 50878 41470 50930 41522
rect 51102 41470 51154 41522
rect 51326 41470 51378 41522
rect 4478 41302 4530 41354
rect 4582 41302 4634 41354
rect 4686 41302 4738 41354
rect 35198 41302 35250 41354
rect 35302 41302 35354 41354
rect 35406 41302 35458 41354
rect 6190 41134 6242 41186
rect 42702 41134 42754 41186
rect 43374 41134 43426 41186
rect 55918 41134 55970 41186
rect 56254 41134 56306 41186
rect 12126 41022 12178 41074
rect 19854 40910 19906 40962
rect 20302 40910 20354 40962
rect 27134 40910 27186 40962
rect 34638 40910 34690 40962
rect 35534 40910 35586 40962
rect 41918 40910 41970 40962
rect 43150 40910 43202 40962
rect 43598 40910 43650 40962
rect 51214 40910 51266 40962
rect 51998 40910 52050 40962
rect 56254 40910 56306 40962
rect 1822 40798 1874 40850
rect 2382 40798 2434 40850
rect 6302 40798 6354 40850
rect 8990 40798 9042 40850
rect 9550 40798 9602 40850
rect 16606 40798 16658 40850
rect 19294 40798 19346 40850
rect 22766 40798 22818 40850
rect 25454 40798 25506 40850
rect 25790 40798 25842 40850
rect 31838 40798 31890 40850
rect 36430 40798 36482 40850
rect 38446 40798 38498 40850
rect 38894 40798 38946 40850
rect 47966 40798 48018 40850
rect 52670 40798 52722 40850
rect 53006 40798 53058 40850
rect 53342 40798 53394 40850
rect 54798 40798 54850 40850
rect 20750 40686 20802 40738
rect 21534 40686 21586 40738
rect 21870 40686 21922 40738
rect 22318 40686 22370 40738
rect 35982 40686 36034 40738
rect 37886 40686 37938 40738
rect 39678 40686 39730 40738
rect 47070 40686 47122 40738
rect 47742 40686 47794 40738
rect 48302 40686 48354 40738
rect 49534 40686 49586 40738
rect 49982 40686 50034 40738
rect 50542 40686 50594 40738
rect 50654 40686 50706 40738
rect 54238 40686 54290 40738
rect 55470 40686 55522 40738
rect 4622 40574 4674 40626
rect 4958 40574 5010 40626
rect 5742 40574 5794 40626
rect 7982 40574 8034 40626
rect 8654 40574 8706 40626
rect 11678 40574 11730 40626
rect 16158 40574 16210 40626
rect 17278 40574 17330 40626
rect 31278 40574 31330 40626
rect 33182 40574 33234 40626
rect 35086 40574 35138 40626
rect 39566 40574 39618 40626
rect 42702 40574 42754 40626
rect 45390 40574 45442 40626
rect 49198 40574 49250 40626
rect 53678 40574 53730 40626
rect 5630 40462 5682 40514
rect 7870 40462 7922 40514
rect 26574 40462 26626 40514
rect 47294 40462 47346 40514
rect 19838 40294 19890 40346
rect 19942 40294 19994 40346
rect 20046 40294 20098 40346
rect 50558 40294 50610 40346
rect 50662 40294 50714 40346
rect 50766 40294 50818 40346
rect 30382 40126 30434 40178
rect 48638 40126 48690 40178
rect 1822 40014 1874 40066
rect 4846 40014 4898 40066
rect 5294 40014 5346 40066
rect 8542 40014 8594 40066
rect 8878 40014 8930 40066
rect 12574 40014 12626 40066
rect 21310 40014 21362 40066
rect 23662 40014 23714 40066
rect 24670 40014 24722 40066
rect 35086 40014 35138 40066
rect 41022 40014 41074 40066
rect 44494 40014 44546 40066
rect 44942 40014 44994 40066
rect 45390 40014 45442 40066
rect 46398 40014 46450 40066
rect 53902 40014 53954 40066
rect 18174 39902 18226 39954
rect 20862 39902 20914 39954
rect 22542 39902 22594 39954
rect 26350 39902 26402 39954
rect 33406 39902 33458 39954
rect 33854 39902 33906 39954
rect 36542 39902 36594 39954
rect 37550 39902 37602 39954
rect 38446 39902 38498 39954
rect 45726 39902 45778 39954
rect 49086 39902 49138 39954
rect 49646 39902 49698 39954
rect 50206 39902 50258 39954
rect 51102 39902 51154 39954
rect 54350 39902 54402 39954
rect 55694 39902 55746 39954
rect 2158 39790 2210 39842
rect 2718 39790 2770 39842
rect 5742 39790 5794 39842
rect 6302 39790 6354 39842
rect 9774 39790 9826 39842
rect 10334 39790 10386 39842
rect 12910 39790 12962 39842
rect 13470 39790 13522 39842
rect 17502 39790 17554 39842
rect 20190 39790 20242 39842
rect 21646 39790 21698 39842
rect 30718 39790 30770 39842
rect 32062 39790 32114 39842
rect 35758 39790 35810 39842
rect 37998 39790 38050 39842
rect 38782 39790 38834 39842
rect 41470 39790 41522 39842
rect 41918 39790 41970 39842
rect 48190 39790 48242 39842
rect 49422 39790 49474 39842
rect 50430 39790 50482 39842
rect 50654 39796 50706 39848
rect 50878 39790 50930 39842
rect 51774 39790 51826 39842
rect 52110 39790 52162 39842
rect 52446 39790 52498 39842
rect 52894 39790 52946 39842
rect 53230 39790 53282 39842
rect 53566 39790 53618 39842
rect 55022 39790 55074 39842
rect 57262 39790 57314 39842
rect 16830 39678 16882 39730
rect 25454 39678 25506 39730
rect 31166 39678 31218 39730
rect 31726 39678 31778 39730
rect 34078 39678 34130 39730
rect 39790 39678 39842 39730
rect 40238 39678 40290 39730
rect 44046 39678 44098 39730
rect 13358 39566 13410 39618
rect 32398 39566 32450 39618
rect 41022 39566 41074 39618
rect 41806 39566 41858 39618
rect 47518 39566 47570 39618
rect 32958 39454 33010 39506
rect 51214 39454 51266 39506
rect 56814 39454 56866 39506
rect 4478 39286 4530 39338
rect 4582 39286 4634 39338
rect 4686 39286 4738 39338
rect 35198 39286 35250 39338
rect 35302 39286 35354 39338
rect 35406 39286 35458 39338
rect 6078 39118 6130 39170
rect 52558 39118 52610 39170
rect 53230 39118 53282 39170
rect 55806 39118 55858 39170
rect 56814 39118 56866 39170
rect 17166 39006 17218 39058
rect 34638 39006 34690 39058
rect 35086 39006 35138 39058
rect 53454 39006 53506 39058
rect 55358 39006 55410 39058
rect 5630 38894 5682 38946
rect 13470 38894 13522 38946
rect 34862 38894 34914 38946
rect 35310 38894 35362 38946
rect 44270 38894 44322 38946
rect 52782 38894 52834 38946
rect 53230 38894 53282 38946
rect 53566 38894 53618 38946
rect 53790 38894 53842 38946
rect 54126 38894 54178 38946
rect 56478 38894 56530 38946
rect 56926 38894 56978 38946
rect 1822 38782 1874 38834
rect 2382 38782 2434 38834
rect 6190 38782 6242 38834
rect 9662 38782 9714 38834
rect 10222 38782 10274 38834
rect 19854 38782 19906 38834
rect 23774 38782 23826 38834
rect 24110 38782 24162 38834
rect 24446 38782 24498 38834
rect 24782 38782 24834 38834
rect 25902 38782 25954 38834
rect 36990 38782 37042 38834
rect 37326 38782 37378 38834
rect 37662 38782 37714 38834
rect 38558 38782 38610 38834
rect 39118 38782 39170 38834
rect 42030 38782 42082 38834
rect 45390 38782 45442 38834
rect 47630 38782 47682 38834
rect 48974 38782 49026 38834
rect 49310 38782 49362 38834
rect 49646 38782 49698 38834
rect 54238 38782 54290 38834
rect 55582 38782 55634 38834
rect 4958 38670 5010 38722
rect 5742 38670 5794 38722
rect 12798 38670 12850 38722
rect 13582 38670 13634 38722
rect 20638 38670 20690 38722
rect 25342 38670 25394 38722
rect 26574 38670 26626 38722
rect 27358 38670 27410 38722
rect 30158 38670 30210 38722
rect 30606 38670 30658 38722
rect 36430 38670 36482 38722
rect 39790 38670 39842 38722
rect 40462 38670 40514 38722
rect 40798 38670 40850 38722
rect 41134 38670 41186 38722
rect 42590 38670 42642 38722
rect 43262 38670 43314 38722
rect 44942 38670 44994 38722
rect 46734 38670 46786 38722
rect 48190 38670 48242 38722
rect 48638 38670 48690 38722
rect 50094 38670 50146 38722
rect 50766 38670 50818 38722
rect 51438 38670 51490 38722
rect 53790 38670 53842 38722
rect 54686 38670 54738 38722
rect 56030 38670 56082 38722
rect 4622 38558 4674 38610
rect 6638 38558 6690 38610
rect 8878 38558 8930 38610
rect 9326 38558 9378 38610
rect 12462 38558 12514 38610
rect 16830 38558 16882 38610
rect 19182 38558 19234 38610
rect 33854 38558 33906 38610
rect 37998 38558 38050 38610
rect 41470 38558 41522 38610
rect 19838 38278 19890 38330
rect 19942 38278 19994 38330
rect 20046 38278 20098 38330
rect 50558 38278 50610 38330
rect 50662 38278 50714 38330
rect 50766 38278 50818 38330
rect 40238 38110 40290 38162
rect 47630 38110 47682 38162
rect 48190 38110 48242 38162
rect 1822 37998 1874 38050
rect 2270 37998 2322 38050
rect 5742 37998 5794 38050
rect 13022 37998 13074 38050
rect 20862 37998 20914 38050
rect 23102 37998 23154 38050
rect 23774 37998 23826 38050
rect 33182 37998 33234 38050
rect 47742 37998 47794 38050
rect 48190 37998 48242 38050
rect 49758 37998 49810 38050
rect 55806 37998 55858 38050
rect 18398 37886 18450 37938
rect 25230 37886 25282 37938
rect 27358 37886 27410 37938
rect 31726 37886 31778 37938
rect 32174 37886 32226 37938
rect 38894 37886 38946 37938
rect 42030 37886 42082 37938
rect 43262 37886 43314 37938
rect 44606 37886 44658 37938
rect 46510 37886 46562 37938
rect 49086 37886 49138 37938
rect 53790 37886 53842 37938
rect 55022 37886 55074 37938
rect 2606 37774 2658 37826
rect 3054 37774 3106 37826
rect 3614 37774 3666 37826
rect 10222 37774 10274 37826
rect 10782 37774 10834 37826
rect 13358 37774 13410 37826
rect 13918 37774 13970 37826
rect 17614 37774 17666 37826
rect 25566 37774 25618 37826
rect 31838 37774 31890 37826
rect 33518 37774 33570 37826
rect 38222 37774 38274 37826
rect 41358 37774 41410 37826
rect 41582 37774 41634 37826
rect 41806 37774 41858 37826
rect 42366 37774 42418 37826
rect 42590 37774 42642 37826
rect 46286 37774 46338 37826
rect 51550 37774 51602 37826
rect 52222 37774 52274 37826
rect 52558 37774 52610 37826
rect 52894 37774 52946 37826
rect 53230 37774 53282 37826
rect 54350 37774 54402 37826
rect 1934 37550 1986 37602
rect 2606 37662 2658 37714
rect 9886 37662 9938 37714
rect 16830 37662 16882 37714
rect 21422 37662 21474 37714
rect 21870 37662 21922 37714
rect 24222 37662 24274 37714
rect 24670 37662 24722 37714
rect 31054 37662 31106 37714
rect 36654 37662 36706 37714
rect 37102 37662 37154 37714
rect 37662 37662 37714 37714
rect 6190 37550 6242 37602
rect 13806 37550 13858 37602
rect 20414 37550 20466 37602
rect 41918 37550 41970 37602
rect 2718 37438 2770 37490
rect 28366 37438 28418 37490
rect 32622 37438 32674 37490
rect 4478 37270 4530 37322
rect 4582 37270 4634 37322
rect 4686 37270 4738 37322
rect 35198 37270 35250 37322
rect 35302 37270 35354 37322
rect 35406 37270 35458 37322
rect 52222 37102 52274 37154
rect 1934 36990 1986 37042
rect 43934 36990 43986 37042
rect 50318 36990 50370 37042
rect 55134 36990 55186 37042
rect 6078 36878 6130 36930
rect 9326 36878 9378 36930
rect 16718 36878 16770 36930
rect 20190 36878 20242 36930
rect 23102 36878 23154 36930
rect 24222 36878 24274 36930
rect 32062 36878 32114 36930
rect 36430 36878 36482 36930
rect 43150 36878 43202 36930
rect 49534 36878 49586 36930
rect 53118 36878 53170 36930
rect 54126 36878 54178 36930
rect 4510 36766 4562 36818
rect 5070 36766 5122 36818
rect 6190 36766 6242 36818
rect 9662 36766 9714 36818
rect 10222 36766 10274 36818
rect 19518 36766 19570 36818
rect 21646 36766 21698 36818
rect 21870 36766 21922 36818
rect 23886 36766 23938 36818
rect 28366 36766 28418 36818
rect 34078 36766 34130 36818
rect 38334 36766 38386 36818
rect 39454 36766 39506 36818
rect 42702 36766 42754 36818
rect 45950 36766 46002 36818
rect 48190 36766 48242 36818
rect 51774 36766 51826 36818
rect 56030 36766 56082 36818
rect 57486 36766 57538 36818
rect 5630 36654 5682 36706
rect 22094 36654 22146 36706
rect 26014 36654 26066 36706
rect 37550 36654 37602 36706
rect 37774 36654 37826 36706
rect 38670 36654 38722 36706
rect 39118 36654 39170 36706
rect 39790 36654 39842 36706
rect 40574 36654 40626 36706
rect 41246 36654 41298 36706
rect 41918 36654 41970 36706
rect 44270 36654 44322 36706
rect 45166 36654 45218 36706
rect 47854 36654 47906 36706
rect 49870 36654 49922 36706
rect 50654 36654 50706 36706
rect 51102 36654 51154 36706
rect 51326 36654 51378 36706
rect 52782 36654 52834 36706
rect 54574 36654 54626 36706
rect 57598 36654 57650 36706
rect 2270 36542 2322 36594
rect 5742 36542 5794 36594
rect 12462 36542 12514 36594
rect 12798 36542 12850 36594
rect 13582 36542 13634 36594
rect 16382 36542 16434 36594
rect 18734 36542 18786 36594
rect 20638 36542 20690 36594
rect 21198 36542 21250 36594
rect 23550 36542 23602 36594
rect 27358 36542 27410 36594
rect 29262 36542 29314 36594
rect 31502 36542 31554 36594
rect 37102 36542 37154 36594
rect 40126 36542 40178 36594
rect 43598 36542 43650 36594
rect 49086 36542 49138 36594
rect 13470 36430 13522 36482
rect 27918 36430 27970 36482
rect 42702 36430 42754 36482
rect 43598 36430 43650 36482
rect 19838 36262 19890 36314
rect 19942 36262 19994 36314
rect 20046 36262 20098 36314
rect 50558 36262 50610 36314
rect 50662 36262 50714 36314
rect 50766 36262 50818 36314
rect 17726 36094 17778 36146
rect 19182 36094 19234 36146
rect 20750 36094 20802 36146
rect 36654 36094 36706 36146
rect 37102 36094 37154 36146
rect 1822 35982 1874 36034
rect 3054 35982 3106 36034
rect 6190 35982 6242 36034
rect 14142 35982 14194 36034
rect 36206 35982 36258 36034
rect 36654 35982 36706 36034
rect 39678 35982 39730 36034
rect 55694 35982 55746 36034
rect 56702 35982 56754 36034
rect 11006 35870 11058 35922
rect 18174 35870 18226 35922
rect 18622 35870 18674 35922
rect 18846 35870 18898 35922
rect 20190 35870 20242 35922
rect 23886 35870 23938 35922
rect 25902 35870 25954 35922
rect 26462 35870 26514 35922
rect 27806 35870 27858 35922
rect 37102 35870 37154 35922
rect 43038 35870 43090 35922
rect 49422 35870 49474 35922
rect 50206 35870 50258 35922
rect 54350 35870 54402 35922
rect 3390 35758 3442 35810
rect 3950 35758 4002 35810
rect 6526 35758 6578 35810
rect 11342 35758 11394 35810
rect 11902 35758 11954 35810
rect 19630 35758 19682 35810
rect 20302 35758 20354 35810
rect 21086 35758 21138 35810
rect 21870 35758 21922 35810
rect 24558 35758 24610 35810
rect 27022 35758 27074 35810
rect 29822 35758 29874 35810
rect 31838 35758 31890 35810
rect 33518 35758 33570 35810
rect 37662 35758 37714 35810
rect 37886 35758 37938 35810
rect 38334 35758 38386 35810
rect 40350 35758 40402 35810
rect 41246 35758 41298 35810
rect 42814 35758 42866 35810
rect 44046 35758 44098 35810
rect 44382 35758 44434 35810
rect 50654 35758 50706 35810
rect 51102 35758 51154 35810
rect 52110 35758 52162 35810
rect 52334 35758 52386 35810
rect 16382 35646 16434 35698
rect 16830 35646 16882 35698
rect 17614 35646 17666 35698
rect 21534 35646 21586 35698
rect 26574 35646 26626 35698
rect 33182 35646 33234 35698
rect 34078 35646 34130 35698
rect 41694 35646 41746 35698
rect 44494 35646 44546 35698
rect 44942 35646 44994 35698
rect 45390 35646 45442 35698
rect 48974 35646 49026 35698
rect 50094 35646 50146 35698
rect 52894 35758 52946 35810
rect 53230 35758 53282 35810
rect 53566 35758 53618 35810
rect 53902 35758 53954 35810
rect 55022 35758 55074 35810
rect 57150 35758 57202 35810
rect 52894 35646 52946 35698
rect 56814 35646 56866 35698
rect 14478 35534 14530 35586
rect 31502 35534 31554 35586
rect 40014 35534 40066 35586
rect 40910 35534 40962 35586
rect 43374 35534 43426 35586
rect 25454 35422 25506 35474
rect 33630 35422 33682 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 5630 35086 5682 35138
rect 13470 35086 13522 35138
rect 17278 35086 17330 35138
rect 17726 35086 17778 35138
rect 18174 35086 18226 35138
rect 18734 35086 18786 35138
rect 27134 35086 27186 35138
rect 35310 35086 35362 35138
rect 50766 35086 50818 35138
rect 51102 35086 51154 35138
rect 20750 34974 20802 35026
rect 39678 34974 39730 35026
rect 51886 34974 51938 35026
rect 56142 34974 56194 35026
rect 56702 34974 56754 35026
rect 18398 34862 18450 34914
rect 19854 34862 19906 34914
rect 21422 34862 21474 34914
rect 30606 34862 30658 34914
rect 44046 34862 44098 34914
rect 44942 34862 44994 34914
rect 49422 34862 49474 34914
rect 50766 34862 50818 34914
rect 51214 34862 51266 34914
rect 54686 34862 54738 34914
rect 56142 34862 56194 34914
rect 20414 34750 20466 34802
rect 21310 34750 21362 34802
rect 21534 34750 21586 34802
rect 22878 34750 22930 34802
rect 23326 34750 23378 34802
rect 24894 34750 24946 34802
rect 25678 34750 25730 34802
rect 26686 34750 26738 34802
rect 27806 34750 27858 34802
rect 28030 34750 28082 34802
rect 29486 34750 29538 34802
rect 30942 34750 30994 34802
rect 33742 34750 33794 34802
rect 35198 34750 35250 34802
rect 36990 34750 37042 34802
rect 37214 34750 37266 34802
rect 38110 34750 38162 34802
rect 38334 34750 38386 34802
rect 38670 34750 38722 34802
rect 38894 34750 38946 34802
rect 49870 34750 49922 34802
rect 52782 34750 52834 34802
rect 53006 34750 53058 34802
rect 54910 34750 54962 34802
rect 16606 34638 16658 34690
rect 17726 34638 17778 34690
rect 18174 34638 18226 34690
rect 19182 34638 19234 34690
rect 19630 34638 19682 34690
rect 21758 34638 21810 34690
rect 21982 34638 22034 34690
rect 22430 34638 22482 34690
rect 23774 34638 23826 34690
rect 25118 34638 25170 34690
rect 26014 34638 26066 34690
rect 26126 34638 26178 34690
rect 28366 34638 28418 34690
rect 33966 34638 34018 34690
rect 34862 34638 34914 34690
rect 40014 34638 40066 34690
rect 42814 34638 42866 34690
rect 51550 34638 51602 34690
rect 55694 34638 55746 34690
rect 56590 34638 56642 34690
rect 5742 34526 5794 34578
rect 13582 34526 13634 34578
rect 16270 34526 16322 34578
rect 17054 34526 17106 34578
rect 22318 34526 22370 34578
rect 22766 34526 22818 34578
rect 24670 34526 24722 34578
rect 25230 34526 25282 34578
rect 25454 34526 25506 34578
rect 29374 34526 29426 34578
rect 31726 34526 31778 34578
rect 38670 34526 38722 34578
rect 40686 34526 40738 34578
rect 41358 34526 41410 34578
rect 41806 34526 41858 34578
rect 42254 34526 42306 34578
rect 43150 34526 43202 34578
rect 45390 34526 45442 34578
rect 45838 34526 45890 34578
rect 46286 34526 46338 34578
rect 50318 34526 50370 34578
rect 54014 34526 54066 34578
rect 55246 34526 55298 34578
rect 27358 34414 27410 34466
rect 37326 34414 37378 34466
rect 37998 34414 38050 34466
rect 19838 34246 19890 34298
rect 19942 34246 19994 34298
rect 20046 34246 20098 34298
rect 50558 34246 50610 34298
rect 50662 34246 50714 34298
rect 50766 34246 50818 34298
rect 23438 34078 23490 34130
rect 32286 34078 32338 34130
rect 50206 34078 50258 34130
rect 51102 34078 51154 34130
rect 3278 33966 3330 34018
rect 3726 33966 3778 34018
rect 4062 33966 4114 34018
rect 16830 33966 16882 34018
rect 19854 33966 19906 34018
rect 20862 33966 20914 34018
rect 25342 33966 25394 34018
rect 26462 33966 26514 34018
rect 27022 33966 27074 34018
rect 28814 33966 28866 34018
rect 30270 33966 30322 34018
rect 36542 33966 36594 34018
rect 37214 33966 37266 34018
rect 40350 33966 40402 34018
rect 42142 33966 42194 34018
rect 44718 33966 44770 34018
rect 47182 33966 47234 34018
rect 48190 33966 48242 34018
rect 50206 33966 50258 34018
rect 50654 33966 50706 34018
rect 51102 33966 51154 34018
rect 51550 33966 51602 34018
rect 51998 33966 52050 34018
rect 55022 33966 55074 34018
rect 11902 33854 11954 33906
rect 16382 33854 16434 33906
rect 18846 33854 18898 33906
rect 20974 33854 21026 33906
rect 21310 33854 21362 33906
rect 21982 33854 22034 33906
rect 22430 33854 22482 33906
rect 22654 33854 22706 33906
rect 23886 33854 23938 33906
rect 24334 33854 24386 33906
rect 25790 33854 25842 33906
rect 27358 33854 27410 33906
rect 31278 33854 31330 33906
rect 31838 33854 31890 33906
rect 33630 33854 33682 33906
rect 34190 33854 34242 33906
rect 35534 33854 35586 33906
rect 36206 33854 36258 33906
rect 36878 33854 36930 33906
rect 42366 33854 42418 33906
rect 53118 33854 53170 33906
rect 54350 33854 54402 33906
rect 6302 33742 6354 33794
rect 6862 33742 6914 33794
rect 18286 33742 18338 33794
rect 20190 33742 20242 33794
rect 22206 33742 22258 33794
rect 24110 33742 24162 33794
rect 25118 33742 25170 33794
rect 26014 33742 26066 33794
rect 26686 33742 26738 33794
rect 27582 33742 27634 33794
rect 30718 33742 30770 33794
rect 35086 33742 35138 33794
rect 35310 33742 35362 33794
rect 42254 33742 42306 33794
rect 44270 33742 44322 33794
rect 45726 33742 45778 33794
rect 52670 33742 52722 33794
rect 52894 33742 52946 33794
rect 12126 33630 12178 33682
rect 17726 33630 17778 33682
rect 18958 33630 19010 33682
rect 23214 33630 23266 33682
rect 25566 33630 25618 33682
rect 27246 33630 27298 33682
rect 31166 33630 31218 33682
rect 34302 33630 34354 33682
rect 37998 33630 38050 33682
rect 41022 33630 41074 33682
rect 43822 33630 43874 33682
rect 45390 33630 45442 33682
rect 46062 33630 46114 33682
rect 46734 33630 46786 33682
rect 53902 33630 53954 33682
rect 55806 33630 55858 33682
rect 12238 33518 12290 33570
rect 17838 33518 17890 33570
rect 21646 33518 21698 33570
rect 22206 33518 22258 33570
rect 46062 33518 46114 33570
rect 33182 33406 33234 33458
rect 34638 33406 34690 33458
rect 46846 33406 46898 33458
rect 50654 33406 50706 33458
rect 51550 33406 51602 33458
rect 52222 33406 52274 33458
rect 4478 33238 4530 33290
rect 4582 33238 4634 33290
rect 4686 33238 4738 33290
rect 35198 33238 35250 33290
rect 35302 33238 35354 33290
rect 35406 33238 35458 33290
rect 5742 33070 5794 33122
rect 12910 32958 12962 33010
rect 34414 32958 34466 33010
rect 34750 32958 34802 33010
rect 19742 32846 19794 32898
rect 21758 32846 21810 32898
rect 28590 32846 28642 32898
rect 43486 32846 43538 32898
rect 43934 32846 43986 32898
rect 45054 32846 45106 32898
rect 50654 32846 50706 32898
rect 9774 32734 9826 32786
rect 10110 32734 10162 32786
rect 14030 32734 14082 32786
rect 15262 32734 15314 32786
rect 15710 32734 15762 32786
rect 18398 32734 18450 32786
rect 20190 32734 20242 32786
rect 20638 32734 20690 32786
rect 22094 32734 22146 32786
rect 23550 32734 23602 32786
rect 24334 32734 24386 32786
rect 24446 32734 24498 32786
rect 25342 32734 25394 32786
rect 29822 32734 29874 32786
rect 30830 32734 30882 32786
rect 33518 32734 33570 32786
rect 34078 32734 34130 32786
rect 38222 32734 38274 32786
rect 38334 32734 38386 32786
rect 39790 32734 39842 32786
rect 44270 32734 44322 32786
rect 45390 32734 45442 32786
rect 45726 32734 45778 32786
rect 45838 32734 45890 32786
rect 46062 32734 46114 32786
rect 46846 32734 46898 32786
rect 47070 32734 47122 32786
rect 47294 32734 47346 32786
rect 51886 32734 51938 32786
rect 52894 32734 52946 32786
rect 53230 32734 53282 32786
rect 54014 32734 54066 32786
rect 54126 32734 54178 32786
rect 56590 32734 56642 32786
rect 16382 32622 16434 32674
rect 19070 32622 19122 32674
rect 19518 32622 19570 32674
rect 20302 32622 20354 32674
rect 20414 32622 20466 32674
rect 23662 32622 23714 32674
rect 25902 32622 25954 32674
rect 29486 32622 29538 32674
rect 30046 32622 30098 32674
rect 30494 32622 30546 32674
rect 31502 32622 31554 32674
rect 35086 32622 35138 32674
rect 35534 32622 35586 32674
rect 37102 32622 37154 32674
rect 39118 32622 39170 32674
rect 39454 32622 39506 32674
rect 40126 32622 40178 32674
rect 41022 32622 41074 32674
rect 41582 32622 41634 32674
rect 42254 32622 42306 32674
rect 46622 32622 46674 32674
rect 47966 32622 48018 32674
rect 48414 32622 48466 32674
rect 48974 32622 49026 32674
rect 49758 32622 49810 32674
rect 51326 32622 51378 32674
rect 51774 32622 51826 32674
rect 55022 32622 55074 32674
rect 5630 32510 5682 32562
rect 6078 32510 6130 32562
rect 10894 32510 10946 32562
rect 13470 32510 13522 32562
rect 13582 32510 13634 32562
rect 23214 32510 23266 32562
rect 23886 32510 23938 32562
rect 24110 32510 24162 32562
rect 24670 32510 24722 32562
rect 24894 32510 24946 32562
rect 25118 32510 25170 32562
rect 25566 32510 25618 32562
rect 37550 32510 37602 32562
rect 40462 32510 40514 32562
rect 43038 32510 43090 32562
rect 46846 32510 46898 32562
rect 47630 32510 47682 32562
rect 50206 32510 50258 32562
rect 52894 32510 52946 32562
rect 57038 32510 57090 32562
rect 6190 32398 6242 32450
rect 13918 32398 13970 32450
rect 18622 32398 18674 32450
rect 49310 32398 49362 32450
rect 50878 32398 50930 32450
rect 54686 32398 54738 32450
rect 55582 32398 55634 32450
rect 19838 32230 19890 32282
rect 19942 32230 19994 32282
rect 20046 32230 20098 32282
rect 50558 32230 50610 32282
rect 50662 32230 50714 32282
rect 50766 32230 50818 32282
rect 41694 32062 41746 32114
rect 4174 31950 4226 32002
rect 8878 31950 8930 32002
rect 9886 31950 9938 32002
rect 14142 31950 14194 32002
rect 16942 31950 16994 32002
rect 18174 31950 18226 32002
rect 26014 31950 26066 32002
rect 30494 31950 30546 32002
rect 44382 31950 44434 32002
rect 52558 31950 52610 32002
rect 56814 31950 56866 32002
rect 57150 31950 57202 32002
rect 3838 31838 3890 31890
rect 10334 31838 10386 31890
rect 10446 31838 10498 31890
rect 12238 31838 12290 31890
rect 13806 31838 13858 31890
rect 14814 31838 14866 31890
rect 15374 31838 15426 31890
rect 21310 31838 21362 31890
rect 24222 31838 24274 31890
rect 29374 31838 29426 31890
rect 34078 31838 34130 31890
rect 37326 31838 37378 31890
rect 40126 31838 40178 31890
rect 42814 31838 42866 31890
rect 45054 31838 45106 31890
rect 45726 31838 45778 31890
rect 47854 31838 47906 31890
rect 48862 31838 48914 31890
rect 49870 31838 49922 31890
rect 50430 31838 50482 31890
rect 51998 31838 52050 31890
rect 52894 31838 52946 31890
rect 53230 31838 53282 31890
rect 54350 31838 54402 31890
rect 55694 31838 55746 31890
rect 58158 31838 58210 31890
rect 3390 31726 3442 31778
rect 6414 31726 6466 31778
rect 6974 31726 7026 31778
rect 7422 31726 7474 31778
rect 15150 31726 15202 31778
rect 16382 31726 16434 31778
rect 17390 31726 17442 31778
rect 20862 31726 20914 31778
rect 21422 31726 21474 31778
rect 24670 31726 24722 31778
rect 25230 31726 25282 31778
rect 29710 31726 29762 31778
rect 33854 31726 33906 31778
rect 34302 31726 34354 31778
rect 36654 31726 36706 31778
rect 37102 31726 37154 31778
rect 39006 31726 39058 31778
rect 41134 31726 41186 31778
rect 41358 31726 41410 31778
rect 43038 31726 43090 31778
rect 45390 31726 45442 31778
rect 46062 31726 46114 31778
rect 46622 31726 46674 31778
rect 47182 31726 47234 31778
rect 49086 31726 49138 31778
rect 50094 31726 50146 31778
rect 51326 31726 51378 31778
rect 51550 31726 51602 31778
rect 51774 31726 51826 31778
rect 52446 31726 52498 31778
rect 53566 31726 53618 31778
rect 53902 31726 53954 31778
rect 55022 31726 55074 31778
rect 56478 31726 56530 31778
rect 57374 31726 57426 31778
rect 8542 31614 8594 31666
rect 14366 31614 14418 31666
rect 20190 31614 20242 31666
rect 22206 31614 22258 31666
rect 34750 31614 34802 31666
rect 35982 31614 36034 31666
rect 37326 31614 37378 31666
rect 12910 31502 12962 31554
rect 28030 31502 28082 31554
rect 32510 31502 32562 31554
rect 36990 31502 37042 31554
rect 37774 31614 37826 31666
rect 38558 31614 38610 31666
rect 42926 31614 42978 31666
rect 48750 31614 48802 31666
rect 52222 31614 52274 31666
rect 56814 31614 56866 31666
rect 57710 31614 57762 31666
rect 7310 31390 7362 31442
rect 8990 31390 9042 31442
rect 20414 31390 20466 31442
rect 24558 31390 24610 31442
rect 33966 31390 34018 31442
rect 37662 31390 37714 31442
rect 38110 31390 38162 31442
rect 49422 31390 49474 31442
rect 4478 31222 4530 31274
rect 4582 31222 4634 31274
rect 4686 31222 4738 31274
rect 35198 31222 35250 31274
rect 35302 31222 35354 31274
rect 35406 31222 35458 31274
rect 28478 31054 28530 31106
rect 8766 30942 8818 30994
rect 26014 30942 26066 30994
rect 38782 30942 38834 30994
rect 14926 30830 14978 30882
rect 22878 30830 22930 30882
rect 31166 30830 31218 30882
rect 32062 30830 32114 30882
rect 33742 30830 33794 30882
rect 36990 30830 37042 30882
rect 37662 30830 37714 30882
rect 38222 30830 38274 30882
rect 50206 30830 50258 30882
rect 51214 30830 51266 30882
rect 51550 30830 51602 30882
rect 1822 30718 1874 30770
rect 2382 30718 2434 30770
rect 5630 30718 5682 30770
rect 6190 30718 6242 30770
rect 9886 30718 9938 30770
rect 12462 30718 12514 30770
rect 17950 30718 18002 30770
rect 18622 30718 18674 30770
rect 23214 30718 23266 30770
rect 27470 30718 27522 30770
rect 28590 30718 28642 30770
rect 30158 30712 30210 30764
rect 30828 30718 30880 30770
rect 31502 30718 31554 30770
rect 32622 30718 32674 30770
rect 33070 30718 33122 30770
rect 33406 30718 33458 30770
rect 33854 30718 33906 30770
rect 34974 30718 35026 30770
rect 35198 30718 35250 30770
rect 35422 30718 35474 30770
rect 35646 30718 35698 30770
rect 37326 30718 37378 30770
rect 38446 30718 38498 30770
rect 42142 30718 42194 30770
rect 42366 30718 42418 30770
rect 43374 30718 43426 30770
rect 45950 30718 46002 30770
rect 46510 30718 46562 30770
rect 50990 30718 51042 30770
rect 52670 30718 52722 30770
rect 54014 30718 54066 30770
rect 56142 30718 56194 30770
rect 57598 30718 57650 30770
rect 14030 30606 14082 30658
rect 14702 30606 14754 30658
rect 17614 30606 17666 30658
rect 18286 30606 18338 30658
rect 19070 30606 19122 30658
rect 19742 30606 19794 30658
rect 23998 30606 24050 30658
rect 26686 30606 26738 30658
rect 27022 30606 27074 30658
rect 28142 30606 28194 30658
rect 29150 30606 29202 30658
rect 29934 30606 29986 30658
rect 30606 30606 30658 30658
rect 31278 30606 31330 30658
rect 32846 30606 32898 30658
rect 33630 30606 33682 30658
rect 34638 30606 34690 30658
rect 36430 30606 36482 30658
rect 37886 30606 37938 30658
rect 39118 30606 39170 30658
rect 39454 30606 39506 30658
rect 40798 30606 40850 30658
rect 45166 30606 45218 30658
rect 48750 30606 48802 30658
rect 49758 30606 49810 30658
rect 51326 30606 51378 30658
rect 54462 30606 54514 30658
rect 57262 30606 57314 30658
rect 4622 30494 4674 30546
rect 4958 30494 5010 30546
rect 8318 30494 8370 30546
rect 10558 30494 10610 30546
rect 12126 30494 12178 30546
rect 14366 30494 14418 30546
rect 20414 30494 20466 30546
rect 27246 30494 27298 30546
rect 27806 30494 27858 30546
rect 29486 30494 29538 30546
rect 32958 30494 33010 30546
rect 34302 30494 34354 30546
rect 35086 30494 35138 30546
rect 36094 30494 36146 30546
rect 37550 30494 37602 30546
rect 39790 30494 39842 30546
rect 40462 30494 40514 30546
rect 41134 30494 41186 30546
rect 44382 30494 44434 30546
rect 45502 30494 45554 30546
rect 52110 30494 52162 30546
rect 55022 30494 55074 30546
rect 11678 30382 11730 30434
rect 15038 30382 15090 30434
rect 27022 30382 27074 30434
rect 30046 30382 30098 30434
rect 30718 30382 30770 30434
rect 38110 30382 38162 30434
rect 47630 30382 47682 30434
rect 50654 30382 50706 30434
rect 53006 30382 53058 30434
rect 19838 30214 19890 30266
rect 19942 30214 19994 30266
rect 20046 30214 20098 30266
rect 50558 30214 50610 30266
rect 50662 30214 50714 30266
rect 50766 30214 50818 30266
rect 11790 30046 11842 30098
rect 12126 30046 12178 30098
rect 21422 30046 21474 30098
rect 27134 30046 27186 30098
rect 39902 30046 39954 30098
rect 40462 30046 40514 30098
rect 41694 30046 41746 30098
rect 42142 30046 42194 30098
rect 42590 30046 42642 30098
rect 1822 29934 1874 29986
rect 2830 29934 2882 29986
rect 3726 29934 3778 29986
rect 4062 29934 4114 29986
rect 7310 29934 7362 29986
rect 11678 29934 11730 29986
rect 16270 29934 16322 29986
rect 20414 29934 20466 29986
rect 25678 29934 25730 29986
rect 28478 29934 28530 29986
rect 28814 29934 28866 29986
rect 30494 29934 30546 29986
rect 31838 29934 31890 29986
rect 34750 29934 34802 29986
rect 35086 29934 35138 29986
rect 38222 29934 38274 29986
rect 39230 29934 39282 29986
rect 41246 29934 41298 29986
rect 41694 29934 41746 29986
rect 42590 29934 42642 29986
rect 45726 29934 45778 29986
rect 50318 29934 50370 29986
rect 51662 29934 51714 29986
rect 53902 29934 53954 29986
rect 55694 29934 55746 29986
rect 12574 29822 12626 29874
rect 13134 29822 13186 29874
rect 13246 29822 13298 29874
rect 14926 29822 14978 29874
rect 16158 29822 16210 29874
rect 21870 29822 21922 29874
rect 22318 29822 22370 29874
rect 25902 29822 25954 29874
rect 26574 29822 26626 29874
rect 27022 29822 27074 29874
rect 27134 29822 27186 29874
rect 27470 29822 27522 29874
rect 28142 29822 28194 29874
rect 29150 29822 29202 29874
rect 33518 29822 33570 29874
rect 33854 29822 33906 29874
rect 38334 29822 38386 29874
rect 40910 29822 40962 29874
rect 44718 29822 44770 29874
rect 45390 29822 45442 29874
rect 46286 29822 46338 29874
rect 46846 29822 46898 29874
rect 47518 29822 47570 29874
rect 52894 29822 52946 29874
rect 53230 29822 53282 29874
rect 3278 29710 3330 29762
rect 6302 29710 6354 29762
rect 6862 29710 6914 29762
rect 11118 29710 11170 29762
rect 11230 29710 11282 29762
rect 14366 29710 14418 29762
rect 15934 29710 15986 29762
rect 16382 29710 16434 29762
rect 21086 29710 21138 29762
rect 22094 29710 22146 29762
rect 22990 29710 23042 29762
rect 23102 29710 23154 29762
rect 24222 29710 24274 29762
rect 24446 29710 24498 29762
rect 24670 29710 24722 29762
rect 26126 29710 26178 29762
rect 26350 29710 26402 29762
rect 34190 29710 34242 29762
rect 35422 29710 35474 29762
rect 35646 29710 35698 29762
rect 35870 29716 35922 29768
rect 36094 29710 36146 29762
rect 36654 29710 36706 29762
rect 36878 29710 36930 29762
rect 37102 29710 37154 29762
rect 37326 29710 37378 29762
rect 37886 29710 37938 29762
rect 45054 29710 45106 29762
rect 53566 29710 53618 29762
rect 54462 29710 54514 29762
rect 55022 29710 55074 29762
rect 10446 29598 10498 29650
rect 15038 29598 15090 29650
rect 18062 29598 18114 29650
rect 25678 29598 25730 29650
rect 26686 29598 26738 29650
rect 33182 29598 33234 29650
rect 33854 29598 33906 29650
rect 36766 29598 36818 29650
rect 39902 29598 39954 29650
rect 40350 29598 40402 29650
rect 42142 29598 42194 29650
rect 44382 29598 44434 29650
rect 48862 29598 48914 29650
rect 49870 29598 49922 29650
rect 50766 29598 50818 29650
rect 51214 29598 51266 29650
rect 52334 29598 52386 29650
rect 18398 29486 18450 29538
rect 49870 29486 49922 29538
rect 50878 29486 50930 29538
rect 51326 29486 51378 29538
rect 3166 29374 3218 29426
rect 13918 29374 13970 29426
rect 24110 29374 24162 29426
rect 25230 29374 25282 29426
rect 34974 29374 35026 29426
rect 36206 29374 36258 29426
rect 50990 29374 51042 29426
rect 51214 29374 51266 29426
rect 4478 29206 4530 29258
rect 4582 29206 4634 29258
rect 4686 29206 4738 29258
rect 35198 29206 35250 29258
rect 35302 29206 35354 29258
rect 35406 29206 35458 29258
rect 5630 29038 5682 29090
rect 15486 29038 15538 29090
rect 18734 29038 18786 29090
rect 21646 29038 21698 29090
rect 26350 29038 26402 29090
rect 41246 29038 41298 29090
rect 43038 29038 43090 29090
rect 53790 29038 53842 29090
rect 55582 29038 55634 29090
rect 16942 28926 16994 28978
rect 20638 28926 20690 28978
rect 35086 28926 35138 28978
rect 38446 28926 38498 28978
rect 15150 28814 15202 28866
rect 16606 28814 16658 28866
rect 19854 28814 19906 28866
rect 29150 28814 29202 28866
rect 31166 28814 31218 28866
rect 31614 28814 31666 28866
rect 36430 28814 36482 28866
rect 37102 28814 37154 28866
rect 38446 28814 38498 28866
rect 1822 28702 1874 28754
rect 2382 28702 2434 28754
rect 5742 28702 5794 28754
rect 12350 28702 12402 28754
rect 12910 28702 12962 28754
rect 14030 28702 14082 28754
rect 17390 28702 17442 28754
rect 17726 28702 17778 28754
rect 20302 28702 20354 28754
rect 21310 28702 21362 28754
rect 21758 28702 21810 28754
rect 24446 28702 24498 28754
rect 24670 28702 24722 28754
rect 24894 28702 24946 28754
rect 26462 28702 26514 28754
rect 26686 28702 26738 28754
rect 26910 28702 26962 28754
rect 27134 28702 27186 28754
rect 29486 28702 29538 28754
rect 29934 28702 29986 28754
rect 33294 28702 33346 28754
rect 33742 28702 33794 28754
rect 34302 28702 34354 28754
rect 34526 28702 34578 28754
rect 34750 28702 34802 28754
rect 34974 28702 35026 28754
rect 35310 28702 35362 28754
rect 35646 28702 35698 28754
rect 36878 28702 36930 28754
rect 37214 28702 37266 28754
rect 4958 28590 5010 28642
rect 6078 28590 6130 28642
rect 6190 28590 6242 28642
rect 12238 28590 12290 28642
rect 13470 28590 13522 28642
rect 14478 28590 14530 28642
rect 15038 28590 15090 28642
rect 15934 28590 15986 28642
rect 16494 28590 16546 28642
rect 17950 28590 18002 28642
rect 19182 28590 19234 28642
rect 19630 28590 19682 28642
rect 21534 28590 21586 28642
rect 25118 28590 25170 28642
rect 25790 28590 25842 28642
rect 26014 28590 26066 28642
rect 27358 28590 27410 28642
rect 28030 28590 28082 28642
rect 28254 28590 28306 28642
rect 30718 28590 30770 28642
rect 32398 28590 32450 28642
rect 35534 28590 35586 28642
rect 35982 28590 36034 28642
rect 37438 28590 37490 28642
rect 4510 28478 4562 28530
rect 13582 28478 13634 28530
rect 24334 28478 24386 28530
rect 25566 28478 25618 28530
rect 27806 28478 27858 28530
rect 30382 28478 30434 28530
rect 32062 28478 32114 28530
rect 32734 28478 32786 28530
rect 33070 28478 33122 28530
rect 37998 28478 38050 28530
rect 45950 28926 46002 28978
rect 46510 28926 46562 28978
rect 46846 28926 46898 28978
rect 42142 28814 42194 28866
rect 43038 28814 43090 28866
rect 45950 28814 46002 28866
rect 46398 28814 46450 28866
rect 50542 28814 50594 28866
rect 52782 28814 52834 28866
rect 53230 28814 53282 28866
rect 54126 28814 54178 28866
rect 39342 28702 39394 28754
rect 40238 28702 40290 28754
rect 41246 28702 41298 28754
rect 47070 28702 47122 28754
rect 47630 28702 47682 28754
rect 48078 28702 48130 28754
rect 48302 28702 48354 28754
rect 55694 28702 55746 28754
rect 42590 28590 42642 28642
rect 54574 28590 54626 28642
rect 12798 28366 12850 28418
rect 25342 28366 25394 28418
rect 27582 28366 27634 28418
rect 38894 28478 38946 28530
rect 41694 28478 41746 28530
rect 45054 28478 45106 28530
rect 45502 28478 45554 28530
rect 48974 28478 49026 28530
rect 50094 28478 50146 28530
rect 50990 28478 51042 28530
rect 51662 28478 51714 28530
rect 52110 28478 52162 28530
rect 56702 28478 56754 28530
rect 39230 28366 39282 28418
rect 39902 28366 39954 28418
rect 40910 28366 40962 28418
rect 47518 28366 47570 28418
rect 50094 28366 50146 28418
rect 50990 28366 51042 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 1822 28030 1874 28082
rect 2382 28030 2434 28082
rect 2606 28030 2658 28082
rect 18510 28030 18562 28082
rect 25342 28030 25394 28082
rect 27022 28030 27074 28082
rect 31166 28030 31218 28082
rect 33518 28030 33570 28082
rect 36206 28030 36258 28082
rect 48862 28030 48914 28082
rect 50206 28030 50258 28082
rect 3166 27918 3218 27970
rect 3614 27918 3666 27970
rect 14254 27918 14306 27970
rect 14702 27918 14754 27970
rect 26910 27918 26962 27970
rect 27806 27918 27858 27970
rect 28478 27918 28530 27970
rect 29710 27918 29762 27970
rect 30718 27918 30770 27970
rect 34414 27918 34466 27970
rect 37886 27918 37938 27970
rect 39230 27918 39282 27970
rect 42142 27918 42194 27970
rect 42814 27918 42866 27970
rect 43262 27918 43314 27970
rect 44718 27918 44770 27970
rect 45166 27918 45218 27970
rect 45614 27918 45666 27970
rect 46062 27918 46114 27970
rect 46846 27918 46898 27970
rect 48862 27918 48914 27970
rect 49310 27918 49362 27970
rect 50206 27918 50258 27970
rect 50654 27918 50706 27970
rect 53118 27918 53170 27970
rect 54798 27918 54850 27970
rect 55358 27918 55410 27970
rect 1822 27806 1874 27858
rect 2270 27806 2322 27858
rect 16046 27806 16098 27858
rect 18958 27806 19010 27858
rect 19406 27806 19458 27858
rect 25902 27806 25954 27858
rect 26126 27806 26178 27858
rect 27134 27806 27186 27858
rect 27358 27806 27410 27858
rect 28142 27806 28194 27858
rect 28814 27806 28866 27858
rect 30046 27806 30098 27858
rect 30382 27806 30434 27858
rect 31502 27806 31554 27858
rect 32062 27806 32114 27858
rect 33070 27806 33122 27858
rect 33406 27806 33458 27858
rect 33518 27806 33570 27858
rect 33854 27806 33906 27858
rect 35534 27806 35586 27858
rect 35982 27806 36034 27858
rect 36318 27806 36370 27858
rect 36542 27806 36594 27858
rect 36766 27806 36818 27858
rect 39678 27806 39730 27858
rect 40014 27806 40066 27858
rect 41358 27806 41410 27858
rect 46510 27806 46562 27858
rect 47182 27806 47234 27858
rect 48190 27806 48242 27858
rect 51102 27806 51154 27858
rect 51662 27806 51714 27858
rect 52110 27806 52162 27858
rect 52334 27806 52386 27858
rect 53454 27806 53506 27858
rect 54350 27806 54402 27858
rect 54910 27806 54962 27858
rect 55806 27806 55858 27858
rect 2718 27694 2770 27746
rect 5742 27694 5794 27746
rect 6302 27694 6354 27746
rect 11566 27694 11618 27746
rect 12126 27694 12178 27746
rect 15486 27694 15538 27746
rect 15710 27694 15762 27746
rect 19518 27694 19570 27746
rect 25678 27694 25730 27746
rect 26350 27694 26402 27746
rect 26574 27694 26626 27746
rect 34190 27694 34242 27746
rect 37326 27694 37378 27746
rect 37550 27694 37602 27746
rect 37774 27694 37826 27746
rect 37998 27694 38050 27746
rect 39118 27694 39170 27746
rect 39790 27694 39842 27746
rect 40910 27694 40962 27746
rect 42254 27694 42306 27746
rect 51886 27694 51938 27746
rect 53342 27694 53394 27746
rect 11230 27582 11282 27634
rect 25454 27582 25506 27634
rect 29262 27582 29314 27634
rect 31838 27582 31890 27634
rect 32510 27582 32562 27634
rect 38446 27582 38498 27634
rect 40238 27582 40290 27634
rect 40350 27582 40402 27634
rect 43710 27582 43762 27634
rect 46286 27582 46338 27634
rect 49758 27582 49810 27634
rect 31726 27470 31778 27522
rect 41022 27470 41074 27522
rect 47854 27470 47906 27522
rect 48974 27470 49026 27522
rect 49870 27470 49922 27522
rect 50094 27470 50146 27522
rect 51886 27582 51938 27634
rect 56702 27582 56754 27634
rect 51998 27470 52050 27522
rect 15038 27358 15090 27410
rect 4478 27190 4530 27242
rect 4582 27190 4634 27242
rect 4686 27190 4738 27242
rect 35198 27190 35250 27242
rect 35302 27190 35354 27242
rect 35406 27190 35458 27242
rect 37438 27022 37490 27074
rect 35310 26910 35362 26962
rect 4958 26798 5010 26850
rect 9326 26798 9378 26850
rect 23438 26798 23490 26850
rect 24558 26798 24610 26850
rect 26126 26798 26178 26850
rect 28142 26798 28194 26850
rect 33518 26798 33570 26850
rect 36318 26798 36370 26850
rect 39006 26798 39058 26850
rect 43374 26798 43426 26850
rect 44270 26798 44322 26850
rect 44718 26798 44770 26850
rect 46398 26798 46450 26850
rect 50654 26798 50706 26850
rect 1822 26686 1874 26738
rect 2382 26686 2434 26738
rect 12350 26686 12402 26738
rect 12910 26686 12962 26738
rect 13470 26686 13522 26738
rect 14030 26686 14082 26738
rect 28478 26686 28530 26738
rect 30830 26686 30882 26738
rect 33070 26686 33122 26738
rect 33742 26686 33794 26738
rect 34190 26686 34242 26738
rect 34750 26686 34802 26738
rect 35086 26686 35138 26738
rect 35646 26686 35698 26738
rect 37102 26686 37154 26738
rect 37326 26686 37378 26738
rect 37550 26686 37602 26738
rect 37774 26686 37826 26738
rect 38894 26686 38946 26738
rect 39342 26686 39394 26738
rect 39790 26686 39842 26738
rect 40238 26686 40290 26738
rect 40574 26686 40626 26738
rect 42142 26686 42194 26738
rect 45502 26686 45554 26738
rect 46846 26686 46898 26738
rect 49758 26686 49810 26738
rect 51326 26686 51378 26738
rect 51550 26686 51602 26738
rect 52670 26686 52722 26738
rect 53006 26686 53058 26738
rect 53678 26686 53730 26738
rect 54238 26686 54290 26738
rect 54798 26686 54850 26738
rect 9774 26574 9826 26626
rect 23550 26574 23602 26626
rect 24110 26574 24162 26626
rect 26686 26574 26738 26626
rect 27022 26574 27074 26626
rect 27358 26574 27410 26626
rect 27918 26574 27970 26626
rect 28254 26574 28306 26626
rect 31278 26574 31330 26626
rect 31614 26574 31666 26626
rect 35982 26574 36034 26626
rect 39118 26574 39170 26626
rect 40798 26574 40850 26626
rect 41694 26574 41746 26626
rect 42254 26574 42306 26626
rect 42926 26574 42978 26626
rect 45166 26574 45218 26626
rect 45614 26574 45666 26626
rect 50878 26574 50930 26626
rect 51886 26574 51938 26626
rect 53342 26574 53394 26626
rect 4510 26462 4562 26514
rect 10110 26462 10162 26514
rect 16158 26462 16210 26514
rect 16606 26462 16658 26514
rect 20750 26462 20802 26514
rect 21422 26462 21474 26514
rect 21870 26462 21922 26514
rect 24894 26462 24946 26514
rect 26350 26462 26402 26514
rect 27470 26462 27522 26514
rect 29598 26462 29650 26514
rect 30046 26462 30098 26514
rect 30494 26462 30546 26514
rect 30942 26462 30994 26514
rect 38334 26462 38386 26514
rect 43934 26462 43986 26514
rect 46286 26462 46338 26514
rect 50206 26462 50258 26514
rect 27358 26350 27410 26402
rect 41246 26350 41298 26402
rect 55470 26462 55522 26514
rect 46510 26350 46562 26402
rect 47294 26350 47346 26402
rect 49646 26350 49698 26402
rect 50654 26350 50706 26402
rect 19838 26182 19890 26234
rect 19942 26182 19994 26234
rect 20046 26182 20098 26234
rect 50558 26182 50610 26234
rect 50662 26182 50714 26234
rect 50766 26182 50818 26234
rect 30270 26014 30322 26066
rect 30830 26014 30882 26066
rect 35758 26014 35810 26066
rect 44830 26014 44882 26066
rect 1822 25902 1874 25954
rect 2718 25902 2770 25954
rect 4958 25902 5010 25954
rect 10558 25902 10610 25954
rect 11006 25902 11058 25954
rect 11454 25902 11506 25954
rect 14590 25902 14642 25954
rect 14926 25902 14978 25954
rect 22206 25902 22258 25954
rect 25566 25902 25618 25954
rect 25902 25902 25954 25954
rect 30270 25902 30322 25954
rect 37886 25902 37938 25954
rect 38782 25902 38834 25954
rect 41470 25902 41522 25954
rect 42142 25902 42194 25954
rect 53342 25902 53394 25954
rect 55358 25902 55410 25954
rect 55806 25902 55858 25954
rect 56702 25902 56754 25954
rect 23998 25790 24050 25842
rect 29710 25790 29762 25842
rect 31390 25790 31442 25842
rect 32510 25790 32562 25842
rect 33294 25790 33346 25842
rect 35534 25790 35586 25842
rect 35758 25790 35810 25842
rect 35982 25790 36034 25842
rect 36766 25790 36818 25842
rect 37550 25790 37602 25842
rect 38670 25790 38722 25842
rect 40126 25790 40178 25842
rect 42366 25790 42418 25842
rect 43822 25790 43874 25842
rect 45390 25790 45442 25842
rect 45726 25790 45778 25842
rect 46510 25790 46562 25842
rect 47182 25790 47234 25842
rect 47854 25790 47906 25842
rect 49646 25790 49698 25842
rect 53902 25790 53954 25842
rect 3054 25678 3106 25730
rect 3614 25678 3666 25730
rect 4062 25678 4114 25730
rect 7198 25678 7250 25730
rect 7758 25678 7810 25730
rect 8206 25678 8258 25730
rect 8766 25678 8818 25730
rect 11790 25678 11842 25730
rect 12350 25678 12402 25730
rect 17502 25678 17554 25730
rect 17838 25678 17890 25730
rect 19966 25678 20018 25730
rect 20750 25678 20802 25730
rect 21198 25678 21250 25730
rect 21534 25678 21586 25730
rect 21870 25678 21922 25730
rect 22766 25678 22818 25730
rect 23326 25678 23378 25730
rect 26238 25678 26290 25730
rect 26462 25678 26514 25730
rect 27022 25678 27074 25730
rect 28366 25689 28418 25741
rect 28590 25678 28642 25730
rect 28814 25678 28866 25730
rect 29038 25678 29090 25730
rect 29486 25678 29538 25730
rect 29598 25678 29650 25730
rect 30718 25678 30770 25730
rect 31166 25678 31218 25730
rect 31726 25678 31778 25730
rect 32174 25678 32226 25730
rect 32286 25678 32338 25730
rect 34078 25678 34130 25730
rect 34190 25678 34242 25730
rect 34526 25678 34578 25730
rect 34862 25678 34914 25730
rect 35198 25678 35250 25730
rect 36542 25678 36594 25730
rect 36654 25678 36706 25730
rect 36990 25678 37042 25730
rect 37214 25678 37266 25730
rect 38446 25678 38498 25730
rect 38894 25678 38946 25730
rect 39566 25678 39618 25730
rect 41246 25678 41298 25730
rect 42030 25678 42082 25730
rect 44382 25678 44434 25730
rect 45054 25678 45106 25730
rect 46062 25678 46114 25730
rect 49086 25678 49138 25730
rect 50990 25678 51042 25730
rect 52222 25678 52274 25730
rect 53230 25678 53282 25730
rect 54910 25678 54962 25730
rect 3950 25566 4002 25618
rect 16830 25566 16882 25618
rect 28030 25566 28082 25618
rect 31390 25566 31442 25618
rect 40238 25566 40290 25618
rect 41694 25566 41746 25618
rect 43710 25566 43762 25618
rect 57150 25566 57202 25618
rect 4622 25454 4674 25506
rect 26910 25454 26962 25506
rect 33630 25454 33682 25506
rect 3166 25342 3218 25394
rect 3502 25342 3554 25394
rect 8094 25342 8146 25394
rect 8878 25342 8930 25394
rect 10894 25342 10946 25394
rect 11342 25342 11394 25394
rect 28702 25342 28754 25394
rect 39118 25342 39170 25394
rect 4478 25174 4530 25226
rect 4582 25174 4634 25226
rect 4686 25174 4738 25226
rect 35198 25174 35250 25226
rect 35302 25174 35354 25226
rect 35406 25174 35458 25226
rect 5742 25006 5794 25058
rect 13470 25006 13522 25058
rect 32510 25006 32562 25058
rect 53230 25006 53282 25058
rect 53790 25006 53842 25058
rect 4958 24894 5010 24946
rect 6190 24894 6242 24946
rect 12798 24894 12850 24946
rect 20526 24894 20578 24946
rect 19406 24782 19458 24834
rect 24110 24782 24162 24834
rect 27022 24782 27074 24834
rect 28142 24782 28194 24834
rect 29486 24782 29538 24834
rect 31614 24782 31666 24834
rect 34190 24782 34242 24834
rect 45278 24782 45330 24834
rect 1822 24670 1874 24722
rect 2382 24670 2434 24722
rect 5630 24670 5682 24722
rect 8766 24670 8818 24722
rect 9326 24670 9378 24722
rect 9662 24670 9714 24722
rect 10222 24670 10274 24722
rect 13582 24670 13634 24722
rect 16270 24670 16322 24722
rect 16718 24670 16770 24722
rect 19070 24670 19122 24722
rect 21422 24670 21474 24722
rect 21982 24670 22034 24722
rect 25566 24670 25618 24722
rect 27694 24670 27746 24722
rect 29150 24670 29202 24722
rect 29822 24670 29874 24722
rect 32398 24670 32450 24722
rect 32622 24670 32674 24722
rect 35198 24670 35250 24722
rect 35646 24670 35698 24722
rect 35870 24670 35922 24722
rect 36878 24670 36930 24722
rect 39118 24670 39170 24722
rect 39230 24670 39282 24722
rect 39566 24670 39618 24722
rect 42366 24726 42418 24778
rect 45726 24782 45778 24834
rect 47854 24782 47906 24834
rect 52782 24782 52834 24834
rect 53230 24782 53282 24834
rect 53678 24782 53730 24834
rect 55358 24782 55410 24834
rect 41694 24670 41746 24722
rect 49534 24670 49586 24722
rect 54462 24670 54514 24722
rect 55806 24670 55858 24722
rect 56702 24670 56754 24722
rect 24894 24558 24946 24610
rect 25006 24558 25058 24610
rect 26238 24558 26290 24610
rect 27470 24558 27522 24610
rect 34862 24558 34914 24610
rect 37550 24558 37602 24610
rect 37774 24558 37826 24610
rect 38446 24558 38498 24610
rect 39342 24558 39394 24610
rect 41246 24558 41298 24610
rect 50654 24614 50706 24666
rect 57822 24670 57874 24722
rect 58046 24658 58098 24710
rect 42814 24558 42866 24610
rect 57598 24558 57650 24610
rect 4622 24446 4674 24498
rect 6526 24446 6578 24498
rect 12350 24446 12402 24498
rect 14030 24446 14082 24498
rect 26574 24446 26626 24498
rect 29262 24446 29314 24498
rect 29710 24446 29762 24498
rect 32062 24446 32114 24498
rect 32846 24446 32898 24498
rect 33294 24446 33346 24498
rect 33742 24446 33794 24498
rect 34526 24446 34578 24498
rect 36206 24446 36258 24498
rect 37214 24446 37266 24498
rect 38110 24446 38162 24498
rect 40126 24446 40178 24498
rect 40574 24446 40626 24498
rect 51214 24446 51266 24498
rect 51886 24446 51938 24498
rect 2494 24334 2546 24386
rect 3054 24334 3106 24386
rect 26014 24334 26066 24386
rect 27582 24334 27634 24386
rect 37438 24334 37490 24386
rect 52558 24334 52610 24386
rect 53566 24334 53618 24386
rect 54126 24334 54178 24386
rect 57486 24334 57538 24386
rect 19838 24166 19890 24218
rect 19942 24166 19994 24218
rect 20046 24166 20098 24218
rect 50558 24166 50610 24218
rect 50662 24166 50714 24218
rect 50766 24166 50818 24218
rect 22094 23998 22146 24050
rect 22990 23998 23042 24050
rect 32062 23998 32114 24050
rect 36094 23998 36146 24050
rect 36990 23998 37042 24050
rect 39230 23998 39282 24050
rect 1822 23886 1874 23938
rect 2270 23886 2322 23938
rect 2606 23886 2658 23938
rect 5854 23886 5906 23938
rect 6190 23886 6242 23938
rect 9662 23886 9714 23938
rect 21422 23886 21474 23938
rect 22094 23886 22146 23938
rect 22990 23886 23042 23938
rect 24558 23886 24610 23938
rect 25566 23886 25618 23938
rect 26574 23886 26626 23938
rect 26686 23886 26738 23938
rect 28254 23886 28306 23938
rect 33182 23886 33234 23938
rect 34190 23886 34242 23938
rect 34302 23886 34354 23938
rect 35086 23886 35138 23938
rect 35870 23886 35922 23938
rect 36766 23886 36818 23938
rect 37662 23886 37714 23938
rect 38558 23886 38610 23938
rect 39342 23886 39394 23938
rect 39790 23886 39842 23938
rect 40014 23886 40066 23938
rect 40238 23886 40290 23938
rect 43934 23886 43986 23938
rect 44382 23886 44434 23938
rect 45054 23886 45106 23938
rect 47630 23886 47682 23938
rect 48078 23886 48130 23938
rect 49982 23886 50034 23938
rect 53902 23886 53954 23938
rect 55694 23886 55746 23938
rect 57150 23886 57202 23938
rect 17614 23774 17666 23826
rect 25342 23774 25394 23826
rect 25790 23774 25842 23826
rect 26350 23774 26402 23826
rect 28702 23774 28754 23826
rect 28926 23774 28978 23826
rect 30942 23774 30994 23826
rect 35422 23774 35474 23826
rect 35758 23774 35810 23826
rect 36542 23774 36594 23826
rect 37102 23774 37154 23826
rect 37326 23774 37378 23826
rect 38894 23774 38946 23826
rect 42254 23774 42306 23826
rect 42478 23774 42530 23826
rect 46062 23774 46114 23826
rect 46398 23774 46450 23826
rect 48862 23774 48914 23826
rect 50654 23774 50706 23826
rect 52894 23774 52946 23826
rect 53230 23774 53282 23826
rect 53566 23774 53618 23826
rect 54350 23774 54402 23826
rect 4846 23662 4898 23714
rect 5406 23662 5458 23714
rect 8430 23662 8482 23714
rect 8990 23662 9042 23714
rect 17950 23662 18002 23714
rect 18510 23662 18562 23714
rect 18846 23662 18898 23714
rect 25118 23662 25170 23714
rect 26014 23662 26066 23714
rect 26126 23662 26178 23714
rect 26910 23662 26962 23714
rect 29038 23662 29090 23714
rect 33742 23662 33794 23714
rect 33966 23662 34018 23714
rect 34414 23662 34466 23714
rect 34750 23662 34802 23714
rect 36318 23662 36370 23714
rect 37886 23662 37938 23714
rect 38222 23662 38274 23714
rect 41582 23662 41634 23714
rect 42142 23662 42194 23714
rect 49534 23662 49586 23714
rect 16830 23550 16882 23602
rect 22542 23550 22594 23602
rect 23438 23550 23490 23602
rect 24110 23550 24162 23602
rect 45726 23606 45778 23658
rect 51774 23662 51826 23714
rect 55022 23662 55074 23714
rect 27806 23550 27858 23602
rect 50430 23550 50482 23602
rect 52558 23550 52610 23602
rect 56702 23550 56754 23602
rect 27694 23438 27746 23490
rect 28478 23438 28530 23490
rect 39118 23438 39170 23490
rect 39790 23438 39842 23490
rect 40238 23438 40290 23490
rect 4478 23158 4530 23210
rect 4582 23158 4634 23210
rect 4686 23158 4738 23210
rect 35198 23158 35250 23210
rect 35302 23158 35354 23210
rect 35406 23158 35458 23210
rect 33630 22990 33682 23042
rect 34414 22990 34466 23042
rect 35646 22990 35698 23042
rect 35870 22990 35922 23042
rect 40350 22990 40402 23042
rect 41246 22990 41298 23042
rect 4958 22878 5010 22930
rect 28366 22878 28418 22930
rect 36990 22878 37042 22930
rect 37886 22878 37938 22930
rect 41694 22878 41746 22930
rect 5742 22766 5794 22818
rect 6190 22766 6242 22818
rect 20750 22766 20802 22818
rect 25230 22766 25282 22818
rect 32958 22766 33010 22818
rect 34078 22766 34130 22818
rect 39118 22766 39170 22818
rect 39902 22766 39954 22818
rect 40350 22766 40402 22818
rect 40798 22766 40850 22818
rect 41246 22766 41298 22818
rect 41918 22766 41970 22818
rect 42590 22766 42642 22818
rect 43038 22766 43090 22818
rect 43486 22766 43538 22818
rect 44270 22766 44322 22818
rect 49534 22766 49586 22818
rect 49982 22766 50034 22818
rect 51662 22766 51714 22818
rect 52110 22766 52162 22818
rect 57710 22766 57762 22818
rect 1822 22654 1874 22706
rect 2382 22654 2434 22706
rect 22318 22654 22370 22706
rect 24782 22654 24834 22706
rect 25566 22654 25618 22706
rect 25790 22654 25842 22706
rect 35422 22654 35474 22706
rect 35646 22654 35698 22706
rect 35870 22654 35922 22706
rect 36206 22654 36258 22706
rect 37326 22654 37378 22706
rect 37550 22654 37602 22706
rect 38110 22654 38162 22706
rect 38446 22654 38498 22706
rect 41582 22654 41634 22706
rect 42142 22654 42194 22706
rect 53006 22654 53058 22706
rect 53678 22654 53730 22706
rect 54238 22654 54290 22706
rect 57598 22654 57650 22706
rect 15710 22542 15762 22594
rect 16270 22542 16322 22594
rect 16382 22542 16434 22594
rect 16942 22542 16994 22594
rect 21310 22542 21362 22594
rect 21646 22542 21698 22594
rect 21982 22542 22034 22594
rect 22766 22542 22818 22594
rect 23438 22542 23490 22594
rect 25230 22542 25282 22594
rect 26014 22542 26066 22594
rect 27694 22542 27746 22594
rect 33294 22542 33346 22594
rect 35086 22542 35138 22594
rect 36094 22542 36146 22594
rect 36318 22542 36370 22594
rect 52670 22542 52722 22594
rect 53342 22542 53394 22594
rect 54798 22542 54850 22594
rect 4622 22430 4674 22482
rect 20302 22430 20354 22482
rect 24110 22430 24162 22482
rect 24894 22430 24946 22482
rect 32510 22430 32562 22482
rect 33630 22430 33682 22482
rect 34526 22430 34578 22482
rect 44942 22430 44994 22482
rect 50430 22430 50482 22482
rect 51214 22430 51266 22482
rect 55470 22430 55522 22482
rect 56478 22430 56530 22482
rect 15262 22318 15314 22370
rect 19838 22150 19890 22202
rect 19942 22150 19994 22202
rect 20046 22150 20098 22202
rect 50558 22150 50610 22202
rect 50662 22150 50714 22202
rect 50766 22150 50818 22202
rect 22654 21982 22706 22034
rect 23438 21982 23490 22034
rect 39454 21982 39506 22034
rect 39902 21982 39954 22034
rect 15822 21870 15874 21922
rect 18286 21870 18338 21922
rect 20526 21870 20578 21922
rect 22094 21870 22146 21922
rect 33630 21870 33682 21922
rect 36654 21870 36706 21922
rect 38670 21870 38722 21922
rect 39454 21870 39506 21922
rect 41022 21870 41074 21922
rect 49758 21870 49810 21922
rect 50206 21870 50258 21922
rect 52894 21870 52946 21922
rect 1822 21758 1874 21810
rect 2270 21758 2322 21810
rect 17838 21758 17890 21810
rect 18622 21758 18674 21810
rect 22766 21758 22818 21810
rect 23214 21758 23266 21810
rect 23886 21758 23938 21810
rect 25118 21758 25170 21810
rect 26014 21758 26066 21810
rect 29150 21758 29202 21810
rect 30046 21758 30098 21810
rect 34750 21758 34802 21810
rect 35982 21758 36034 21810
rect 37886 21758 37938 21810
rect 39902 21758 39954 21810
rect 40350 21758 40402 21810
rect 45838 21758 45890 21810
rect 48862 21758 48914 21810
rect 50654 21758 50706 21810
rect 50766 21758 50818 21810
rect 53566 21758 53618 21810
rect 54014 21758 54066 21810
rect 56702 21758 56754 21810
rect 16382 21646 16434 21698
rect 16830 21646 16882 21698
rect 21198 21646 21250 21698
rect 25566 21646 25618 21698
rect 29598 21646 29650 21698
rect 35198 21646 35250 21698
rect 38782 21646 38834 21698
rect 41806 21646 41858 21698
rect 24222 21534 24274 21586
rect 24670 21534 24722 21586
rect 26238 21534 26290 21586
rect 26798 21534 26850 21586
rect 28926 21534 28978 21586
rect 30382 21534 30434 21586
rect 32062 21534 32114 21586
rect 32510 21534 32562 21586
rect 36206 21590 36258 21642
rect 43038 21646 43090 21698
rect 43374 21646 43426 21698
rect 43710 21646 43762 21698
rect 44046 21646 44098 21698
rect 44606 21646 44658 21698
rect 45166 21646 45218 21698
rect 47742 21646 47794 21698
rect 50990 21646 51042 21698
rect 54574 21646 54626 21698
rect 55470 21646 55522 21698
rect 55694 21646 55746 21698
rect 33182 21534 33234 21586
rect 38334 21534 38386 21586
rect 41582 21534 41634 21586
rect 42254 21534 42306 21586
rect 42702 21534 42754 21586
rect 48190 21534 48242 21586
rect 49310 21534 49362 21586
rect 54350 21534 54402 21586
rect 57150 21534 57202 21586
rect 41470 21422 41522 21474
rect 37774 21310 37826 21362
rect 38334 21310 38386 21362
rect 55134 21310 55186 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 25454 20974 25506 21026
rect 29710 20974 29762 21026
rect 39118 20974 39170 21026
rect 39454 20974 39506 21026
rect 43038 20974 43090 21026
rect 50094 20974 50146 21026
rect 56478 20974 56530 21026
rect 24558 20862 24610 20914
rect 24782 20862 24834 20914
rect 25006 20862 25058 20914
rect 40686 20862 40738 20914
rect 45502 20862 45554 20914
rect 16942 20750 16994 20802
rect 19182 20750 19234 20802
rect 19854 20750 19906 20802
rect 20302 20750 20354 20802
rect 20750 20750 20802 20802
rect 25006 20750 25058 20802
rect 26350 20750 26402 20802
rect 28590 20750 28642 20802
rect 34638 20750 34690 20802
rect 35086 20750 35138 20802
rect 35534 20750 35586 20802
rect 35982 20750 36034 20802
rect 41134 20750 41186 20802
rect 45502 20750 45554 20802
rect 45950 20750 46002 20802
rect 46734 20750 46786 20802
rect 47630 20750 47682 20802
rect 51438 20750 51490 20802
rect 51886 20750 51938 20802
rect 56814 20750 56866 20802
rect 57262 20750 57314 20802
rect 14702 20638 14754 20690
rect 21422 20638 21474 20690
rect 23662 20638 23714 20690
rect 29150 20638 29202 20690
rect 36430 20638 36482 20690
rect 37774 20638 37826 20690
rect 21646 20526 21698 20578
rect 25342 20526 25394 20578
rect 37662 20582 37714 20634
rect 38222 20638 38274 20690
rect 38558 20638 38610 20690
rect 39118 20638 39170 20690
rect 40350 20638 40402 20690
rect 43710 20638 43762 20690
rect 45054 20638 45106 20690
rect 46510 20638 46562 20690
rect 46734 20638 46786 20690
rect 48302 20638 48354 20690
rect 52894 20638 52946 20690
rect 54350 20638 54402 20690
rect 55358 20638 55410 20690
rect 55918 20638 55970 20690
rect 33406 20526 33458 20578
rect 39230 20526 39282 20578
rect 40014 20526 40066 20578
rect 41582 20526 41634 20578
rect 43486 20526 43538 20578
rect 44046 20526 44098 20578
rect 46174 20526 46226 20578
rect 48414 20526 48466 20578
rect 50094 20526 50146 20578
rect 53566 20526 53618 20578
rect 25902 20414 25954 20466
rect 33070 20414 33122 20466
rect 34190 20414 34242 20466
rect 37326 20414 37378 20466
rect 42814 20414 42866 20466
rect 54126 20414 54178 20466
rect 54798 20414 54850 20466
rect 47182 20302 47234 20354
rect 19838 20134 19890 20186
rect 19942 20134 19994 20186
rect 20046 20134 20098 20186
rect 50558 20134 50610 20186
rect 50662 20134 50714 20186
rect 50766 20134 50818 20186
rect 25790 19966 25842 20018
rect 31390 19966 31442 20018
rect 16718 19854 16770 19906
rect 23998 19854 24050 19906
rect 25566 19854 25618 19906
rect 27470 19854 27522 19906
rect 34526 19854 34578 19906
rect 38222 19854 38274 19906
rect 45502 19854 45554 19906
rect 49758 19854 49810 19906
rect 55470 19854 55522 19906
rect 17726 19742 17778 19794
rect 18174 19742 18226 19794
rect 19630 19742 19682 19794
rect 26798 19742 26850 19794
rect 33854 19742 33906 19794
rect 34190 19742 34242 19794
rect 36206 19742 36258 19794
rect 38782 19742 38834 19794
rect 40350 19742 40402 19794
rect 49086 19742 49138 19794
rect 50206 19742 50258 19794
rect 51550 19742 51602 19794
rect 53342 19742 53394 19794
rect 54126 19742 54178 19794
rect 54798 19742 54850 19794
rect 16830 19630 16882 19682
rect 17950 19630 18002 19682
rect 18958 19630 19010 19682
rect 19294 19630 19346 19682
rect 23214 19630 23266 19682
rect 26238 19630 26290 19682
rect 28366 19630 28418 19682
rect 31726 19630 31778 19682
rect 36094 19630 36146 19682
rect 36654 19630 36706 19682
rect 37774 19630 37826 19682
rect 40910 19630 40962 19682
rect 41022 19630 41074 19682
rect 41470 19630 41522 19682
rect 42030 19630 42082 19682
rect 44494 19630 44546 19682
rect 46174 19630 46226 19682
rect 46398 19630 46450 19682
rect 48750 19630 48802 19682
rect 49422 19630 49474 19682
rect 50878 19630 50930 19682
rect 52670 19630 52722 19682
rect 53006 19630 53058 19682
rect 53678 19630 53730 19682
rect 20190 19518 20242 19570
rect 22766 19518 22818 19570
rect 26910 19518 26962 19570
rect 29486 19518 29538 19570
rect 32174 19518 32226 19570
rect 33182 19518 33234 19570
rect 47518 19518 47570 19570
rect 52334 19518 52386 19570
rect 56702 19518 56754 19570
rect 33518 19406 33570 19458
rect 40014 19406 40066 19458
rect 18622 19294 18674 19346
rect 27022 19294 27074 19346
rect 27358 19294 27410 19346
rect 45726 19294 45778 19346
rect 46174 19294 46226 19346
rect 4478 19126 4530 19178
rect 4582 19126 4634 19178
rect 4686 19126 4738 19178
rect 35198 19126 35250 19178
rect 35302 19126 35354 19178
rect 35406 19126 35458 19178
rect 31614 18958 31666 19010
rect 32062 18958 32114 19010
rect 41022 18958 41074 19010
rect 51438 18958 51490 19010
rect 52222 18958 52274 19010
rect 35422 18846 35474 18898
rect 35982 18846 36034 18898
rect 50990 18846 51042 18898
rect 51886 18846 51938 18898
rect 54798 18846 54850 18898
rect 17838 18734 17890 18786
rect 20750 18734 20802 18786
rect 25566 18734 25618 18786
rect 26462 18734 26514 18786
rect 27358 18734 27410 18786
rect 30158 18734 30210 18786
rect 30942 18734 30994 18786
rect 31726 18734 31778 18786
rect 33182 18734 33234 18786
rect 34526 18734 34578 18786
rect 35422 18734 35474 18786
rect 35870 18734 35922 18786
rect 37102 18734 37154 18786
rect 38670 18734 38722 18786
rect 39118 18734 39170 18786
rect 43598 18734 43650 18786
rect 46062 18734 46114 18786
rect 51438 18734 51490 18786
rect 54686 18734 54738 18786
rect 15150 18622 15202 18674
rect 24222 18622 24274 18674
rect 25006 18622 25058 18674
rect 30494 18622 30546 18674
rect 32062 18622 32114 18674
rect 34974 18622 35026 18674
rect 46958 18622 47010 18674
rect 47630 18622 47682 18674
rect 52894 18678 52946 18730
rect 47966 18622 48018 18674
rect 57150 18622 57202 18674
rect 26014 18510 26066 18562
rect 28590 18510 28642 18562
rect 34078 18510 34130 18562
rect 36318 18510 36370 18562
rect 39454 18510 39506 18562
rect 40126 18510 40178 18562
rect 45614 18510 45666 18562
rect 47294 18510 47346 18562
rect 48526 18510 48578 18562
rect 49086 18510 49138 18562
rect 49758 18510 49810 18562
rect 50542 18510 50594 18562
rect 53230 18510 53282 18562
rect 55134 18510 55186 18562
rect 57710 18510 57762 18562
rect 22654 18398 22706 18450
rect 39790 18398 39842 18450
rect 41358 18398 41410 18450
rect 50990 18398 51042 18450
rect 51886 18398 51938 18450
rect 51214 18286 51266 18338
rect 51886 18286 51938 18338
rect 19838 18118 19890 18170
rect 19942 18118 19994 18170
rect 20046 18118 20098 18170
rect 50558 18118 50610 18170
rect 50662 18118 50714 18170
rect 50766 18118 50818 18170
rect 23886 17950 23938 18002
rect 24222 17950 24274 18002
rect 24670 17950 24722 18002
rect 30606 17950 30658 18002
rect 31614 17950 31666 18002
rect 49086 17950 49138 18002
rect 16830 17838 16882 17890
rect 22654 17838 22706 17890
rect 24222 17838 24274 17890
rect 24670 17838 24722 17890
rect 27806 17838 27858 17890
rect 30606 17838 30658 17890
rect 31054 17838 31106 17890
rect 31502 17838 31554 17890
rect 39454 17838 39506 17890
rect 39902 17838 39954 17890
rect 41022 17838 41074 17890
rect 41470 17838 41522 17890
rect 46062 17838 46114 17890
rect 48302 17838 48354 17890
rect 51662 17838 51714 17890
rect 53678 17838 53730 17890
rect 25342 17726 25394 17778
rect 27134 17726 27186 17778
rect 28366 17726 28418 17778
rect 29598 17726 29650 17778
rect 33182 17726 33234 17778
rect 35982 17726 36034 17778
rect 42254 17726 42306 17778
rect 43374 17726 43426 17778
rect 52670 17726 52722 17778
rect 53342 17726 53394 17778
rect 54798 17726 54850 17778
rect 55470 17726 55522 17778
rect 17726 17614 17778 17666
rect 26798 17614 26850 17666
rect 27470 17614 27522 17666
rect 28926 17614 28978 17666
rect 33518 17614 33570 17666
rect 33854 17614 33906 17666
rect 34190 17614 34242 17666
rect 34750 17614 34802 17666
rect 35310 17614 35362 17666
rect 41918 17614 41970 17666
rect 42702 17614 42754 17666
rect 48974 17614 49026 17666
rect 49310 17614 49362 17666
rect 53006 17614 53058 17666
rect 54238 17614 54290 17666
rect 18734 17502 18786 17554
rect 23662 17502 23714 17554
rect 26462 17502 26514 17554
rect 32286 17502 32338 17554
rect 36766 17502 36818 17554
rect 40350 17502 40402 17554
rect 47294 17502 47346 17554
rect 47742 17502 47794 17554
rect 49870 17502 49922 17554
rect 50766 17502 50818 17554
rect 51214 17502 51266 17554
rect 52334 17502 52386 17554
rect 51102 17278 51154 17330
rect 51662 17278 51714 17330
rect 4478 17110 4530 17162
rect 4582 17110 4634 17162
rect 4686 17110 4738 17162
rect 35198 17110 35250 17162
rect 35302 17110 35354 17162
rect 35406 17110 35458 17162
rect 55694 16942 55746 16994
rect 35534 16830 35586 16882
rect 20302 16718 20354 16770
rect 22094 16718 22146 16770
rect 22542 16718 22594 16770
rect 22990 16718 23042 16770
rect 23886 16718 23938 16770
rect 28478 16718 28530 16770
rect 45726 16718 45778 16770
rect 50990 16718 51042 16770
rect 24222 16606 24274 16658
rect 24446 16606 24498 16658
rect 24782 16606 24834 16658
rect 25342 16606 25394 16658
rect 29262 16606 29314 16658
rect 30046 16606 30098 16658
rect 32062 16606 32114 16658
rect 45054 16606 45106 16658
rect 45390 16606 45442 16658
rect 53230 16606 53282 16658
rect 53678 16606 53730 16658
rect 54126 16606 54178 16658
rect 54574 16606 54626 16658
rect 54910 16606 54962 16658
rect 55134 16606 55186 16658
rect 55358 16606 55410 16658
rect 55582 16606 55634 16658
rect 56142 16606 56194 16658
rect 23438 16494 23490 16546
rect 27806 16494 27858 16546
rect 30830 16494 30882 16546
rect 31054 16494 31106 16546
rect 31502 16494 31554 16546
rect 34414 16494 34466 16546
rect 39678 16494 39730 16546
rect 40014 16494 40066 16546
rect 40350 16494 40402 16546
rect 41134 16494 41186 16546
rect 41806 16494 41858 16546
rect 46958 16494 47010 16546
rect 56590 16494 56642 16546
rect 40686 16382 40738 16434
rect 42478 16382 42530 16434
rect 47294 16382 47346 16434
rect 48414 16382 48466 16434
rect 48862 16382 48914 16434
rect 49646 16382 49698 16434
rect 50094 16382 50146 16434
rect 50542 16382 50594 16434
rect 51438 16382 51490 16434
rect 52110 16382 52162 16434
rect 53454 16382 53506 16434
rect 57038 16382 57090 16434
rect 57486 16382 57538 16434
rect 30382 16270 30434 16322
rect 19838 16102 19890 16154
rect 19942 16102 19994 16154
rect 20046 16102 20098 16154
rect 50558 16102 50610 16154
rect 50662 16102 50714 16154
rect 50766 16102 50818 16154
rect 28030 15934 28082 15986
rect 31278 15934 31330 15986
rect 51102 15934 51154 15986
rect 51438 15934 51490 15986
rect 51774 15934 51826 15986
rect 23214 15822 23266 15874
rect 23662 15822 23714 15874
rect 24110 15822 24162 15874
rect 37102 15822 37154 15874
rect 39230 15822 39282 15874
rect 40238 15822 40290 15874
rect 41246 15822 41298 15874
rect 42142 15822 42194 15874
rect 49198 15822 49250 15874
rect 49534 15822 49586 15874
rect 50094 15822 50146 15874
rect 50990 15822 51042 15874
rect 51438 15822 51490 15874
rect 52334 15822 52386 15874
rect 53678 15822 53730 15874
rect 19742 15710 19794 15762
rect 24670 15710 24722 15762
rect 25230 15710 25282 15762
rect 29710 15710 29762 15762
rect 32174 15710 32226 15762
rect 37550 15710 37602 15762
rect 38558 15710 38610 15762
rect 48190 15710 48242 15762
rect 53006 15710 53058 15762
rect 53342 15710 53394 15762
rect 54238 15710 54290 15762
rect 55470 15710 55522 15762
rect 17726 15598 17778 15650
rect 30494 15598 30546 15650
rect 31726 15598 31778 15650
rect 32958 15598 33010 15650
rect 33182 15598 33234 15650
rect 33742 15598 33794 15650
rect 34190 15598 34242 15650
rect 36654 15598 36706 15650
rect 37998 15598 38050 15650
rect 48974 15598 49026 15650
rect 49646 15598 49698 15650
rect 52670 15598 52722 15650
rect 54798 15598 54850 15650
rect 28926 15486 28978 15538
rect 32398 15486 32450 15538
rect 38670 15486 38722 15538
rect 41694 15486 41746 15538
rect 47294 15486 47346 15538
rect 47742 15486 47794 15538
rect 50542 15486 50594 15538
rect 51886 15486 51938 15538
rect 20190 15374 20242 15426
rect 48638 15374 48690 15426
rect 4478 15094 4530 15146
rect 4582 15094 4634 15146
rect 4686 15094 4738 15146
rect 35198 15094 35250 15146
rect 35302 15094 35354 15146
rect 35406 15094 35458 15146
rect 33854 14926 33906 14978
rect 19294 14814 19346 14866
rect 20190 14814 20242 14866
rect 29262 14814 29314 14866
rect 29822 14814 29874 14866
rect 30158 14814 30210 14866
rect 42254 14814 42306 14866
rect 19182 14702 19234 14754
rect 27134 14702 27186 14754
rect 29262 14702 29314 14754
rect 30158 14702 30210 14754
rect 35982 14702 36034 14754
rect 36430 14702 36482 14754
rect 37326 14702 37378 14754
rect 51774 14702 51826 14754
rect 56254 14702 56306 14754
rect 19630 14590 19682 14642
rect 23886 14590 23938 14642
rect 25006 14590 25058 14642
rect 27582 14590 27634 14642
rect 35086 14590 35138 14642
rect 37774 14590 37826 14642
rect 37886 14590 37938 14642
rect 38222 14590 38274 14642
rect 39006 14590 39058 14642
rect 43822 14590 43874 14642
rect 44942 14590 44994 14642
rect 48638 14590 48690 14642
rect 48974 14590 49026 14642
rect 49310 14590 49362 14642
rect 49870 14590 49922 14642
rect 52894 14590 52946 14642
rect 57038 14590 57090 14642
rect 20078 14478 20130 14530
rect 21422 14478 21474 14530
rect 22206 14478 22258 14530
rect 22878 14478 22930 14530
rect 23214 14478 23266 14530
rect 23550 14478 23602 14530
rect 24446 14478 24498 14530
rect 26686 14478 26738 14530
rect 28254 14478 28306 14530
rect 31278 14478 31330 14530
rect 41246 14478 41298 14530
rect 44270 14478 44322 14530
rect 45502 14478 45554 14530
rect 47854 14478 47906 14530
rect 48302 14478 48354 14530
rect 50430 14478 50482 14530
rect 51102 14478 51154 14530
rect 52670 14478 52722 14530
rect 54462 14478 54514 14530
rect 54910 14478 54962 14530
rect 56142 14478 56194 14530
rect 21870 14366 21922 14418
rect 22542 14366 22594 14418
rect 25678 14366 25730 14418
rect 28702 14366 28754 14418
rect 29710 14366 29762 14418
rect 30942 14366 30994 14418
rect 35534 14366 35586 14418
rect 19854 14254 19906 14306
rect 20078 14254 20130 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 54798 13918 54850 13970
rect 19182 13806 19234 13858
rect 24446 13806 24498 13858
rect 25342 13806 25394 13858
rect 25790 13806 25842 13858
rect 26686 13806 26738 13858
rect 29150 13806 29202 13858
rect 30942 13806 30994 13858
rect 32062 13806 32114 13858
rect 32510 13806 32562 13858
rect 33294 13806 33346 13858
rect 33630 13806 33682 13858
rect 36318 13806 36370 13858
rect 38110 13806 38162 13858
rect 46062 13806 46114 13858
rect 54574 13806 54626 13858
rect 56030 13806 56082 13858
rect 16830 13694 16882 13746
rect 18407 13694 18459 13746
rect 20078 13694 20130 13746
rect 23326 13694 23378 13746
rect 28590 13694 28642 13746
rect 35646 13694 35698 13746
rect 36766 13694 36818 13746
rect 41134 13694 41186 13746
rect 45390 13694 45442 13746
rect 46622 13694 46674 13746
rect 47182 13694 47234 13746
rect 47854 13694 47906 13746
rect 50542 13694 50594 13746
rect 54238 13694 54290 13746
rect 54910 13694 54962 13746
rect 55022 13694 55074 13746
rect 17502 13582 17554 13634
rect 19742 13582 19794 13634
rect 20414 13582 20466 13634
rect 20974 13582 21026 13634
rect 35310 13582 35362 13634
rect 35982 13582 36034 13634
rect 37438 13582 37490 13634
rect 38894 13582 38946 13634
rect 41694 13582 41746 13634
rect 43710 13582 43762 13634
rect 45054 13582 45106 13634
rect 45726 13582 45778 13634
rect 52670 13582 52722 13634
rect 26238 13470 26290 13522
rect 39790 13470 39842 13522
rect 44494 13470 44546 13522
rect 55582 13470 55634 13522
rect 4478 13078 4530 13130
rect 4582 13078 4634 13130
rect 4686 13078 4738 13130
rect 35198 13078 35250 13130
rect 35302 13078 35354 13130
rect 35406 13078 35458 13130
rect 19294 12798 19346 12850
rect 42590 12798 42642 12850
rect 55918 12798 55970 12850
rect 22430 12686 22482 12738
rect 27022 12686 27074 12738
rect 33742 12686 33794 12738
rect 48302 12686 48354 12738
rect 50990 12686 51042 12738
rect 51550 12686 51602 12738
rect 51886 12686 51938 12738
rect 52782 12686 52834 12738
rect 53902 12686 53954 12738
rect 17502 12574 17554 12626
rect 23662 12574 23714 12626
rect 24334 12574 24386 12626
rect 24894 12574 24946 12626
rect 30382 12574 30434 12626
rect 31614 12574 31666 12626
rect 39454 12574 39506 12626
rect 46734 12574 46786 12626
rect 55358 12574 55410 12626
rect 18958 12462 19010 12514
rect 21310 12462 21362 12514
rect 23326 12462 23378 12514
rect 23998 12462 24050 12514
rect 25454 12462 25506 12514
rect 30046 12462 30098 12514
rect 30718 12462 30770 12514
rect 32174 12462 32226 12514
rect 38446 12462 38498 12514
rect 38558 12462 38610 12514
rect 39230 12462 39282 12514
rect 53678 12462 53730 12514
rect 26126 12350 26178 12402
rect 31054 12350 31106 12402
rect 32846 12350 32898 12402
rect 35534 12350 35586 12402
rect 35982 12350 36034 12402
rect 36430 12350 36482 12402
rect 37326 12350 37378 12402
rect 37774 12350 37826 12402
rect 38222 12350 38274 12402
rect 46398 12350 46450 12402
rect 19838 12070 19890 12122
rect 19942 12070 19994 12122
rect 20046 12070 20098 12122
rect 50558 12070 50610 12122
rect 50662 12070 50714 12122
rect 50766 12070 50818 12122
rect 22766 11902 22818 11954
rect 23326 11902 23378 11954
rect 31054 11902 31106 11954
rect 31726 11902 31778 11954
rect 30606 11790 30658 11842
rect 52782 11790 52834 11842
rect 53790 11790 53842 11842
rect 20526 11678 20578 11730
rect 25902 11678 25954 11730
rect 29486 11678 29538 11730
rect 31166 11678 31218 11730
rect 36766 11678 36818 11730
rect 37662 11678 37714 11730
rect 40462 11678 40514 11730
rect 42366 11678 42418 11730
rect 44382 11678 44434 11730
rect 48862 11678 48914 11730
rect 53342 11678 53394 11730
rect 19742 11566 19794 11618
rect 22542 11566 22594 11618
rect 25454 11566 25506 11618
rect 26350 11566 26402 11618
rect 26798 11566 26850 11618
rect 27134 11566 27186 11618
rect 29822 11566 29874 11618
rect 33630 11566 33682 11618
rect 36318 11566 36370 11618
rect 41470 11566 41522 11618
rect 42030 11566 42082 11618
rect 52334 11566 52386 11618
rect 19406 11454 19458 11506
rect 22990 11454 23042 11506
rect 23438 11454 23490 11506
rect 24670 11454 24722 11506
rect 31614 11454 31666 11506
rect 32062 11454 32114 11506
rect 32510 11454 32562 11506
rect 33070 11454 33122 11506
rect 35870 11454 35922 11506
rect 37326 11454 37378 11506
rect 41022 11454 41074 11506
rect 45614 11454 45666 11506
rect 31614 11230 31666 11282
rect 32398 11230 32450 11282
rect 4478 11062 4530 11114
rect 4582 11062 4634 11114
rect 4686 11062 4738 11114
rect 35198 11062 35250 11114
rect 35302 11062 35354 11114
rect 35406 11062 35458 11114
rect 20302 10894 20354 10946
rect 20750 10894 20802 10946
rect 36990 10894 37042 10946
rect 25118 10782 25170 10834
rect 35310 10782 35362 10834
rect 47854 10782 47906 10834
rect 20302 10670 20354 10722
rect 21422 10670 21474 10722
rect 30382 10670 30434 10722
rect 30830 10670 30882 10722
rect 31278 10670 31330 10722
rect 35982 10670 36034 10722
rect 36430 10670 36482 10722
rect 41582 10670 41634 10722
rect 42030 10670 42082 10722
rect 43598 10670 43650 10722
rect 53118 10670 53170 10722
rect 31614 10558 31666 10610
rect 34190 10558 34242 10610
rect 37774 10558 37826 10610
rect 38894 10558 38946 10610
rect 39118 10558 39170 10610
rect 41134 10558 41186 10610
rect 44046 10558 44098 10610
rect 45166 10558 45218 10610
rect 45390 10558 45442 10610
rect 45502 10558 45554 10610
rect 20750 10446 20802 10498
rect 21870 10446 21922 10498
rect 22318 10446 22370 10498
rect 24446 10446 24498 10498
rect 32398 10446 32450 10498
rect 38670 10446 38722 10498
rect 25790 10334 25842 10386
rect 19838 10054 19890 10106
rect 19942 10054 19994 10106
rect 20046 10054 20098 10106
rect 50558 10054 50610 10106
rect 50662 10054 50714 10106
rect 50766 10054 50818 10106
rect 23662 9886 23714 9938
rect 24670 9886 24722 9938
rect 30158 9886 30210 9938
rect 33518 9886 33570 9938
rect 34526 9886 34578 9938
rect 18174 9774 18226 9826
rect 22878 9774 22930 9826
rect 23662 9774 23714 9826
rect 24222 9774 24274 9826
rect 25678 9774 25730 9826
rect 33518 9774 33570 9826
rect 33966 9774 34018 9826
rect 44494 9774 44546 9826
rect 21310 9662 21362 9714
rect 24670 9662 24722 9714
rect 18622 9550 18674 9602
rect 19070 9550 19122 9602
rect 21646 9550 21698 9602
rect 26014 9550 26066 9602
rect 26574 9550 26626 9602
rect 28814 9550 28866 9602
rect 34526 9550 34578 9602
rect 35198 9550 35250 9602
rect 37550 9438 37602 9490
rect 4478 9046 4530 9098
rect 4582 9046 4634 9098
rect 4686 9046 4738 9098
rect 35198 9046 35250 9098
rect 35302 9046 35354 9098
rect 35406 9046 35458 9098
rect 26238 8878 26290 8930
rect 21646 8766 21698 8818
rect 22990 8766 23042 8818
rect 32174 8766 32226 8818
rect 21646 8654 21698 8706
rect 22094 8654 22146 8706
rect 22542 8654 22594 8706
rect 22990 8654 23042 8706
rect 28142 8654 28194 8706
rect 36430 8654 36482 8706
rect 37102 8654 37154 8706
rect 23662 8542 23714 8594
rect 23774 8542 23826 8594
rect 24894 8542 24946 8594
rect 28590 8542 28642 8594
rect 29262 8542 29314 8594
rect 29598 8542 29650 8594
rect 23998 8430 24050 8482
rect 27694 8430 27746 8482
rect 31726 8318 31778 8370
rect 19838 8038 19890 8090
rect 19942 8038 19994 8090
rect 20046 8038 20098 8090
rect 50558 8038 50610 8090
rect 50662 8038 50714 8090
rect 50766 8038 50818 8090
rect 3838 7758 3890 7810
rect 4286 7758 4338 7810
rect 22318 7758 22370 7810
rect 22766 7758 22818 7810
rect 28254 7758 28306 7810
rect 28702 7758 28754 7810
rect 29598 7758 29650 7810
rect 32286 7758 32338 7810
rect 29150 7646 29202 7698
rect 30606 7646 30658 7698
rect 31614 7646 31666 7698
rect 30270 7534 30322 7586
rect 30382 7534 30434 7586
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6022 19890 6074
rect 19942 6022 19994 6074
rect 20046 6022 20098 6074
rect 50558 6022 50610 6074
rect 50662 6022 50714 6074
rect 50766 6022 50818 6074
rect 4478 5014 4530 5066
rect 4582 5014 4634 5066
rect 4686 5014 4738 5066
rect 35198 5014 35250 5066
rect 35302 5014 35354 5066
rect 35406 5014 35458 5066
rect 19838 4006 19890 4058
rect 19942 4006 19994 4058
rect 20046 4006 20098 4058
rect 50558 4006 50610 4058
rect 50662 4006 50714 4058
rect 50766 4006 50818 4058
<< metal2 >>
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 4476 55468 4740 55478
rect 4532 55412 4580 55468
rect 4636 55412 4684 55468
rect 4476 55402 4740 55412
rect 35196 55468 35460 55478
rect 35252 55412 35300 55468
rect 35356 55412 35404 55468
rect 35196 55402 35460 55412
rect 19836 54460 20100 54470
rect 19892 54404 19940 54460
rect 19996 54404 20044 54460
rect 19836 54394 20100 54404
rect 50556 54460 50820 54470
rect 50612 54404 50660 54460
rect 50716 54404 50764 54460
rect 50556 54394 50820 54404
rect 3836 54178 3892 54190
rect 3836 54126 3838 54178
rect 3890 54126 3892 54178
rect 3836 53844 3892 54126
rect 56028 54180 56084 54190
rect 56028 54178 56196 54180
rect 56028 54126 56030 54178
rect 56082 54126 56196 54178
rect 56028 54124 56196 54126
rect 56028 54114 56084 54124
rect 3836 53778 3892 53788
rect 56140 53844 56196 54124
rect 56140 53778 56196 53788
rect 4476 53452 4740 53462
rect 4532 53396 4580 53452
rect 4636 53396 4684 53452
rect 4476 53386 4740 53396
rect 35196 53452 35460 53462
rect 35252 53396 35300 53452
rect 35356 53396 35404 53452
rect 35196 53386 35460 53396
rect 19836 52444 20100 52454
rect 19892 52388 19940 52444
rect 19996 52388 20044 52444
rect 19836 52378 20100 52388
rect 50556 52444 50820 52454
rect 50612 52388 50660 52444
rect 50716 52388 50764 52444
rect 50556 52378 50820 52388
rect 4476 51436 4740 51446
rect 4532 51380 4580 51436
rect 4636 51380 4684 51436
rect 4476 51370 4740 51380
rect 35196 51436 35460 51446
rect 35252 51380 35300 51436
rect 35356 51380 35404 51436
rect 35196 51370 35460 51380
rect 19836 50428 20100 50438
rect 19892 50372 19940 50428
rect 19996 50372 20044 50428
rect 19836 50362 20100 50372
rect 50556 50428 50820 50438
rect 50612 50372 50660 50428
rect 50716 50372 50764 50428
rect 50556 50362 50820 50372
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 32060 49138 32116 49150
rect 32060 49086 32062 49138
rect 32114 49086 32116 49138
rect 32060 49026 32116 49086
rect 32060 48974 32062 49026
rect 32114 48974 32116 49026
rect 32060 48962 32116 48974
rect 33516 49138 33572 49150
rect 33516 49086 33518 49138
rect 33570 49086 33572 49138
rect 21420 48802 21476 48814
rect 21420 48750 21422 48802
rect 21474 48750 21476 48802
rect 19836 48412 20100 48422
rect 19892 48356 19940 48412
rect 19996 48356 20044 48412
rect 19836 48346 20100 48356
rect 19852 48018 19908 48030
rect 19852 47966 19854 48018
rect 19906 47966 19908 48018
rect 19516 47908 19572 47918
rect 19516 47814 19572 47852
rect 19068 47794 19124 47806
rect 19068 47742 19070 47794
rect 19122 47742 19124 47794
rect 19068 47684 19124 47742
rect 19852 47684 19908 47966
rect 19068 47628 19908 47684
rect 20188 47908 20244 47918
rect 4476 47404 4740 47414
rect 4532 47348 4580 47404
rect 4636 47348 4684 47404
rect 4476 47338 4740 47348
rect 17836 46786 17892 46798
rect 17836 46734 17838 46786
rect 17890 46734 17892 46786
rect 17388 46676 17444 46686
rect 17388 46674 17556 46676
rect 17388 46622 17390 46674
rect 17442 46622 17556 46674
rect 17388 46620 17556 46622
rect 17388 46610 17444 46620
rect 17500 45780 17556 46620
rect 17836 45892 17892 46734
rect 18508 46676 18564 46686
rect 19068 46676 19124 47628
rect 18508 46674 19124 46676
rect 18508 46622 18510 46674
rect 18562 46622 19124 46674
rect 18508 46620 19124 46622
rect 20188 47236 20244 47852
rect 21420 47236 21476 48750
rect 23100 48804 23156 48814
rect 21868 48690 21924 48702
rect 22316 48692 22372 48702
rect 21868 48638 21870 48690
rect 21922 48638 21924 48690
rect 21644 47236 21700 47246
rect 21420 47180 21644 47236
rect 17948 45892 18004 45902
rect 17836 45890 18004 45892
rect 17836 45838 17950 45890
rect 18002 45838 18004 45890
rect 17836 45836 18004 45838
rect 17500 45778 17668 45780
rect 17500 45726 17502 45778
rect 17554 45726 17668 45778
rect 17500 45724 17668 45726
rect 17500 45714 17556 45724
rect 4476 45388 4740 45398
rect 4532 45332 4580 45388
rect 4636 45332 4684 45388
rect 4476 45322 4740 45332
rect 17500 45332 17556 45342
rect 17164 44884 17220 44894
rect 17164 44790 17220 44828
rect 17500 44882 17556 45276
rect 17500 44830 17502 44882
rect 17554 44830 17556 44882
rect 17500 44818 17556 44830
rect 17612 44884 17668 45724
rect 17948 45332 18004 45836
rect 17948 45266 18004 45276
rect 18284 45892 18340 45902
rect 18508 45892 18564 46620
rect 19836 46396 20100 46406
rect 19892 46340 19940 46396
rect 19996 46340 20044 46396
rect 19836 46330 20100 46340
rect 18284 45890 18564 45892
rect 18284 45838 18286 45890
rect 18338 45838 18564 45890
rect 18284 45836 18564 45838
rect 17612 44818 17668 44828
rect 18060 44884 18116 44894
rect 18284 44884 18340 45836
rect 20188 45332 20244 47180
rect 20636 47124 20692 47134
rect 20524 46676 20580 46686
rect 20636 46676 20692 47068
rect 20524 46674 20692 46676
rect 20524 46622 20526 46674
rect 20578 46622 20692 46674
rect 20524 46620 20692 46622
rect 21644 47010 21700 47180
rect 21644 46958 21646 47010
rect 21698 46958 21700 47010
rect 20524 46610 20580 46620
rect 21644 46562 21700 46958
rect 21644 46510 21646 46562
rect 21698 46510 21700 46562
rect 21644 46498 21700 46510
rect 21868 47012 21924 48638
rect 22092 48690 22708 48692
rect 22092 48638 22318 48690
rect 22370 48638 22708 48690
rect 22092 48636 22708 48638
rect 22092 48018 22148 48636
rect 22316 48626 22372 48636
rect 22092 47966 22094 48018
rect 22146 47966 22148 48018
rect 22092 47954 22148 47966
rect 20524 46116 20580 46126
rect 20524 45892 20580 46060
rect 20188 45266 20244 45276
rect 20300 45890 20580 45892
rect 20300 45838 20526 45890
rect 20578 45838 20580 45890
rect 20300 45836 20580 45838
rect 18116 44828 18340 44884
rect 18060 43764 18116 44828
rect 20300 44658 20356 45836
rect 20524 45826 20580 45836
rect 21756 45778 21812 45790
rect 21756 45726 21758 45778
rect 21810 45726 21812 45778
rect 21308 45332 21364 45342
rect 21308 44770 21364 45276
rect 21308 44718 21310 44770
rect 21362 44718 21364 44770
rect 21308 44706 21364 44718
rect 20300 44606 20302 44658
rect 20354 44606 20356 44658
rect 19836 44380 20100 44390
rect 19892 44324 19940 44380
rect 19996 44324 20044 44380
rect 19836 44314 20100 44324
rect 20300 44210 20356 44606
rect 20300 44158 20302 44210
rect 20354 44158 20356 44210
rect 20300 44098 20356 44158
rect 20300 44046 20302 44098
rect 20354 44046 20356 44098
rect 18060 43698 18116 43708
rect 19628 43876 19684 43886
rect 19628 43764 19684 43820
rect 19852 43764 19908 43774
rect 19628 43762 19908 43764
rect 19628 43710 19854 43762
rect 19906 43710 19908 43762
rect 19628 43708 19908 43710
rect 4476 43372 4740 43382
rect 4532 43316 4580 43372
rect 4636 43316 4684 43372
rect 4476 43306 4740 43316
rect 7532 42866 7588 42878
rect 7532 42814 7534 42866
rect 7586 42814 7588 42866
rect 7196 42642 7252 42654
rect 7196 42590 7198 42642
rect 7250 42590 7252 42642
rect 6860 42084 6916 42094
rect 7196 42084 7252 42590
rect 6860 42082 7252 42084
rect 6860 42030 6862 42082
rect 6914 42030 7252 42082
rect 6860 42028 7252 42030
rect 4060 41858 4116 41870
rect 4060 41806 4062 41858
rect 4114 41806 4116 41858
rect 1820 41748 1876 41758
rect 1708 41692 1820 41748
rect 1708 40404 1764 41692
rect 1820 41654 1876 41692
rect 3724 41748 3780 41758
rect 1820 40850 1876 40862
rect 1820 40798 1822 40850
rect 1874 40798 1876 40850
rect 1820 40516 1876 40798
rect 1820 40450 1876 40460
rect 2380 40850 2436 40862
rect 2380 40798 2382 40850
rect 2434 40798 2436 40850
rect 1708 40068 1764 40348
rect 2380 40404 2436 40798
rect 3724 40740 3780 41692
rect 3724 40674 3780 40684
rect 2380 40338 2436 40348
rect 2716 40516 2772 40526
rect 1820 40068 1876 40078
rect 1708 40066 1988 40068
rect 1708 40014 1822 40066
rect 1874 40014 1988 40066
rect 1708 40012 1988 40014
rect 1820 40002 1876 40012
rect 1820 38836 1876 38846
rect 1708 38834 1876 38836
rect 1708 38782 1822 38834
rect 1874 38782 1876 38834
rect 1708 38780 1876 38782
rect 1708 36932 1764 38780
rect 1820 38770 1876 38780
rect 1820 38052 1876 38062
rect 1932 38052 1988 40012
rect 2156 39842 2212 39854
rect 2156 39790 2158 39842
rect 2210 39790 2212 39842
rect 2156 38948 2212 39790
rect 2716 39842 2772 40460
rect 4060 40404 4116 41806
rect 4620 41860 4676 41870
rect 4620 41766 4676 41804
rect 6188 41860 6244 41870
rect 4476 41356 4740 41366
rect 4532 41300 4580 41356
rect 4636 41300 4684 41356
rect 4476 41290 4740 41300
rect 6188 41188 6244 41804
rect 5852 41186 6244 41188
rect 5852 41134 6190 41186
rect 6242 41134 6244 41186
rect 5852 41132 6244 41134
rect 4620 40740 4676 40750
rect 4620 40628 4676 40684
rect 4620 40626 4900 40628
rect 4620 40574 4622 40626
rect 4674 40574 4900 40626
rect 4620 40572 4900 40574
rect 4620 40562 4676 40572
rect 4060 40338 4116 40348
rect 2716 39790 2718 39842
rect 2770 39790 2772 39842
rect 2716 39778 2772 39790
rect 4844 40066 4900 40572
rect 4844 40014 4846 40066
rect 4898 40014 4900 40066
rect 4476 39340 4740 39350
rect 4532 39284 4580 39340
rect 4636 39284 4684 39340
rect 4476 39274 4740 39284
rect 2380 38948 2436 38958
rect 2156 38892 2380 38948
rect 2380 38834 2436 38892
rect 2380 38782 2382 38834
rect 2434 38782 2436 38834
rect 2380 38770 2436 38782
rect 4620 38612 4676 38622
rect 4844 38612 4900 40014
rect 4956 40626 5012 40638
rect 4956 40574 4958 40626
rect 5010 40574 5012 40626
rect 4956 39620 5012 40574
rect 5740 40626 5796 40638
rect 5740 40574 5742 40626
rect 5794 40574 5796 40626
rect 5628 40516 5684 40526
rect 5628 40422 5684 40460
rect 5740 40180 5796 40574
rect 5292 40124 5796 40180
rect 5292 40066 5348 40124
rect 5292 40014 5294 40066
rect 5346 40014 5348 40066
rect 5292 40002 5348 40014
rect 5740 39844 5796 39854
rect 5852 39844 5908 41132
rect 6188 41122 6244 41132
rect 6300 41636 6356 41646
rect 6300 40850 6356 41580
rect 6300 40798 6302 40850
rect 6354 40798 6356 40850
rect 6300 40786 6356 40798
rect 6860 40628 6916 42028
rect 7196 41636 7252 41646
rect 7196 41542 7252 41580
rect 6860 40562 6916 40572
rect 6300 40516 6356 40526
rect 5740 39842 5908 39844
rect 5740 39790 5742 39842
rect 5794 39790 5908 39842
rect 5740 39788 5908 39790
rect 6076 40404 6132 40414
rect 5740 39778 5796 39788
rect 4956 39554 5012 39564
rect 6076 39170 6132 40348
rect 6300 39842 6356 40460
rect 7532 40516 7588 42814
rect 8092 42866 8148 42878
rect 8092 42814 8094 42866
rect 8146 42814 8148 42866
rect 8092 41972 8148 42814
rect 9772 42644 9828 42654
rect 8092 41906 8148 41916
rect 8988 41972 9044 41982
rect 8988 40850 9044 41916
rect 9660 41972 9716 41982
rect 9660 41878 9716 41916
rect 9772 41970 9828 42588
rect 9772 41918 9774 41970
rect 9826 41918 9828 41970
rect 9772 41906 9828 41918
rect 10220 42642 10276 42654
rect 10220 42590 10222 42642
rect 10274 42590 10276 42642
rect 8988 40798 8990 40850
rect 9042 40798 9044 40850
rect 8988 40786 9044 40798
rect 9548 41524 9604 41534
rect 9548 40852 9604 41468
rect 9548 40850 9828 40852
rect 9548 40798 9550 40850
rect 9602 40798 9828 40850
rect 9548 40796 9828 40798
rect 9548 40786 9604 40796
rect 7980 40626 8036 40638
rect 7980 40574 7982 40626
rect 8034 40574 8036 40626
rect 7532 40450 7588 40460
rect 7868 40516 7924 40526
rect 7868 40422 7924 40460
rect 7980 40068 8036 40574
rect 8652 40628 8708 40638
rect 7980 40002 8036 40012
rect 8540 40068 8596 40078
rect 8652 40068 8708 40572
rect 8540 40066 8708 40068
rect 8540 40014 8542 40066
rect 8594 40014 8708 40066
rect 8540 40012 8708 40014
rect 8540 40002 8596 40012
rect 6300 39790 6302 39842
rect 6354 39790 6356 39842
rect 6300 39778 6356 39790
rect 6076 39118 6078 39170
rect 6130 39118 6132 39170
rect 6076 39106 6132 39118
rect 6188 39620 6244 39630
rect 5628 38948 5684 38958
rect 5628 38854 5684 38892
rect 6188 38834 6244 39564
rect 6188 38782 6190 38834
rect 6242 38782 6244 38834
rect 6188 38770 6244 38782
rect 4956 38724 5012 38734
rect 4956 38630 5012 38668
rect 5740 38724 5796 38734
rect 5740 38630 5796 38668
rect 8652 38724 8708 40012
rect 8876 40068 8932 40078
rect 8876 39974 8932 40012
rect 9772 39842 9828 40796
rect 10220 40628 10276 42590
rect 10668 42644 10724 42654
rect 10668 42550 10724 42588
rect 19292 41972 19348 41982
rect 19292 41878 19348 41916
rect 19516 41970 19572 41982
rect 19516 41918 19518 41970
rect 19570 41918 19572 41970
rect 11004 41860 11060 41870
rect 11004 41766 11060 41804
rect 12124 41860 12180 41870
rect 10892 41524 10948 41534
rect 10892 41430 10948 41468
rect 12124 41074 12180 41804
rect 19516 41636 19572 41918
rect 19628 41748 19684 43708
rect 19852 43698 19908 43708
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19628 41692 19908 41748
rect 19516 41570 19572 41580
rect 12124 41022 12126 41074
rect 12178 41022 12180 41074
rect 12124 41010 12180 41022
rect 19852 40964 19908 41692
rect 19852 40870 19908 40908
rect 20188 40964 20244 40974
rect 16604 40850 16660 40862
rect 16604 40798 16606 40850
rect 16658 40798 16660 40850
rect 10220 40562 10276 40572
rect 11676 40626 11732 40638
rect 11676 40574 11678 40626
rect 11730 40574 11732 40626
rect 11676 40292 11732 40574
rect 16156 40628 16212 40638
rect 16604 40628 16660 40798
rect 18284 40852 18340 40862
rect 16156 40626 16660 40628
rect 16156 40574 16158 40626
rect 16210 40574 16660 40626
rect 16156 40572 16660 40574
rect 16156 40562 16212 40572
rect 11676 40236 11844 40292
rect 11788 40068 11844 40236
rect 11788 40002 11844 40012
rect 12572 40068 12628 40078
rect 9772 39790 9774 39842
rect 9826 39790 9828 39842
rect 9772 39778 9828 39790
rect 10332 39842 10388 39854
rect 10332 39790 10334 39842
rect 10386 39790 10388 39842
rect 9660 39620 9716 39630
rect 9660 38834 9716 39564
rect 10332 39620 10388 39790
rect 10332 39554 10388 39564
rect 9660 38782 9662 38834
rect 9714 38782 9716 38834
rect 9660 38770 9716 38782
rect 10220 38948 10276 38958
rect 10220 38834 10276 38892
rect 10220 38782 10222 38834
rect 10274 38782 10276 38834
rect 4620 38610 4900 38612
rect 4620 38558 4622 38610
rect 4674 38558 4900 38610
rect 4620 38556 4900 38558
rect 4620 38546 4676 38556
rect 2268 38052 2324 38062
rect 1820 38050 2324 38052
rect 1820 37998 1822 38050
rect 1874 37998 2270 38050
rect 2322 37998 2324 38050
rect 1820 37996 2324 37998
rect 1820 37986 1876 37996
rect 1932 37602 1988 37614
rect 1932 37550 1934 37602
rect 1986 37550 1988 37602
rect 1932 37042 1988 37550
rect 1932 36990 1934 37042
rect 1986 36990 1988 37042
rect 1932 36978 1988 36990
rect 1820 36932 1876 36942
rect 1708 36876 1820 36932
rect 1820 36866 1876 36876
rect 2268 36596 2324 37996
rect 4844 38052 4900 38556
rect 6636 38612 6692 38622
rect 8652 38612 8708 38668
rect 8876 38612 8932 38622
rect 9324 38612 9380 38622
rect 8652 38610 9380 38612
rect 8652 38558 8878 38610
rect 8930 38558 9326 38610
rect 9378 38558 9380 38610
rect 8652 38556 9380 38558
rect 4844 37986 4900 37996
rect 5740 38052 5796 38062
rect 5740 37958 5796 37996
rect 6300 38052 6356 38062
rect 2604 37826 2660 37838
rect 2604 37774 2606 37826
rect 2658 37774 2660 37826
rect 2604 37714 2660 37774
rect 2604 37662 2606 37714
rect 2658 37662 2660 37714
rect 2604 37650 2660 37662
rect 3052 37826 3108 37838
rect 3052 37774 3054 37826
rect 3106 37774 3108 37826
rect 2716 37490 2772 37502
rect 2716 37438 2718 37490
rect 2770 37438 2772 37490
rect 2716 36932 2772 37438
rect 2716 36866 2772 36876
rect 3052 36708 3108 37774
rect 3612 37826 3668 37838
rect 3612 37774 3614 37826
rect 3666 37774 3668 37826
rect 3612 36820 3668 37774
rect 6188 37602 6244 37614
rect 6188 37550 6190 37602
rect 6242 37550 6244 37602
rect 4476 37324 4740 37334
rect 4532 37268 4580 37324
rect 4636 37268 4684 37324
rect 4476 37258 4740 37268
rect 3612 36754 3668 36764
rect 4508 36932 4564 36942
rect 4508 36818 4564 36876
rect 6076 36930 6132 36942
rect 6076 36878 6078 36930
rect 6130 36878 6132 36930
rect 4508 36766 4510 36818
rect 4562 36766 4564 36818
rect 4508 36754 4564 36766
rect 5068 36820 5124 36830
rect 5068 36726 5124 36764
rect 6076 36820 6132 36878
rect 6076 36754 6132 36764
rect 6188 36818 6244 37550
rect 6188 36766 6190 36818
rect 6242 36766 6244 36818
rect 6188 36754 6244 36766
rect 3052 36642 3108 36652
rect 3836 36708 3892 36718
rect 5628 36708 5684 36718
rect 3892 36652 4004 36708
rect 3836 36642 3892 36652
rect 1820 36594 2996 36596
rect 1820 36542 2270 36594
rect 2322 36542 2996 36594
rect 1820 36540 2996 36542
rect 1820 36034 1876 36540
rect 2268 36530 2324 36540
rect 1820 35982 1822 36034
rect 1874 35982 1876 36034
rect 1820 35970 1876 35982
rect 2940 36036 2996 36540
rect 3052 36036 3108 36046
rect 2940 36034 3332 36036
rect 2940 35982 3054 36034
rect 3106 35982 3332 36034
rect 2940 35980 3332 35982
rect 3052 35970 3108 35980
rect 3276 34020 3332 35980
rect 3388 35810 3444 35822
rect 3388 35758 3390 35810
rect 3442 35758 3444 35810
rect 3388 35140 3444 35758
rect 3948 35810 4004 36652
rect 5628 36614 5684 36652
rect 5740 36596 5796 36606
rect 5740 36594 6132 36596
rect 5740 36542 5742 36594
rect 5794 36542 6132 36594
rect 5740 36540 6132 36542
rect 5740 36530 5796 36540
rect 3948 35758 3950 35810
rect 4002 35758 4004 35810
rect 3948 35746 4004 35758
rect 4172 36372 4228 36382
rect 3388 35074 3444 35084
rect 4172 34692 4228 36316
rect 6076 35812 6132 36540
rect 6188 36036 6244 36046
rect 6300 36036 6356 37996
rect 6636 38052 6692 38556
rect 8876 38546 8932 38556
rect 6636 37986 6692 37996
rect 9324 36932 9380 38556
rect 10220 37826 10276 38782
rect 12460 38612 12516 38622
rect 12572 38612 12628 40012
rect 12908 39844 12964 39854
rect 13468 39844 13524 39854
rect 12908 39842 13524 39844
rect 12908 39790 12910 39842
rect 12962 39790 13470 39842
rect 13522 39790 13524 39842
rect 12908 39788 13524 39790
rect 12908 39778 12964 39788
rect 13468 39778 13524 39788
rect 16604 39732 16660 40572
rect 17276 40626 17332 40638
rect 17276 40574 17278 40626
rect 17330 40574 17332 40626
rect 17164 39956 17220 39966
rect 16828 39732 16884 39742
rect 16604 39730 16884 39732
rect 16604 39678 16830 39730
rect 16882 39678 16884 39730
rect 16604 39676 16884 39678
rect 13356 39620 13412 39630
rect 13356 39526 13412 39564
rect 13468 38948 13524 38958
rect 13468 38854 13524 38892
rect 12796 38724 12852 38734
rect 12796 38630 12852 38668
rect 13580 38724 13636 38734
rect 13580 38630 13636 38668
rect 16828 38724 16884 39676
rect 17164 39058 17220 39900
rect 17164 39006 17166 39058
rect 17218 39006 17220 39058
rect 17164 38994 17220 39006
rect 12460 38610 12628 38612
rect 12460 38558 12462 38610
rect 12514 38558 12628 38610
rect 12460 38556 12628 38558
rect 12460 38546 12516 38556
rect 12572 38052 12628 38556
rect 16828 38610 16884 38668
rect 16828 38558 16830 38610
rect 16882 38558 16884 38610
rect 13020 38052 13076 38062
rect 12460 38050 13076 38052
rect 12460 37998 13022 38050
rect 13074 37998 13076 38050
rect 12460 37996 13076 37998
rect 10220 37774 10222 37826
rect 10274 37774 10276 37826
rect 10220 37762 10276 37774
rect 10780 37826 10836 37838
rect 10780 37774 10782 37826
rect 10834 37774 10836 37826
rect 9884 37714 9940 37726
rect 9884 37662 9886 37714
rect 9938 37662 9940 37714
rect 9324 36838 9380 36876
rect 9660 37604 9716 37614
rect 9660 36818 9716 37548
rect 9660 36766 9662 36818
rect 9714 36766 9716 36818
rect 9660 36754 9716 36766
rect 9884 36932 9940 37662
rect 10780 37604 10836 37774
rect 10780 37538 10836 37548
rect 6188 36034 6356 36036
rect 6188 35982 6190 36034
rect 6242 35982 6356 36034
rect 6188 35980 6356 35982
rect 6188 35970 6244 35980
rect 9884 35924 9940 36876
rect 10220 36818 10276 36830
rect 10220 36766 10222 36818
rect 10274 36766 10276 36818
rect 10220 36484 10276 36766
rect 12460 36594 12516 37996
rect 12460 36542 12462 36594
rect 12514 36542 12516 36594
rect 12460 36530 12516 36542
rect 12796 36596 12852 36606
rect 12796 36502 12852 36540
rect 10220 36418 10276 36428
rect 11340 36484 11396 36494
rect 9884 35858 9940 35868
rect 11004 35924 11060 35934
rect 11004 35830 11060 35868
rect 6524 35812 6580 35822
rect 6076 35810 6580 35812
rect 6076 35758 6526 35810
rect 6578 35758 6580 35810
rect 6076 35756 6580 35758
rect 6524 35746 6580 35756
rect 11340 35810 11396 36428
rect 13020 35924 13076 37996
rect 13356 37828 13412 37838
rect 13916 37828 13972 37838
rect 13356 37826 13972 37828
rect 13356 37774 13358 37826
rect 13410 37774 13918 37826
rect 13970 37774 13972 37826
rect 13356 37772 13972 37774
rect 13356 37762 13412 37772
rect 13916 37762 13972 37772
rect 16828 37714 16884 38558
rect 16828 37662 16830 37714
rect 16882 37662 16884 37714
rect 13804 37604 13860 37614
rect 13804 37510 13860 37548
rect 16716 36932 16772 36942
rect 16716 36838 16772 36876
rect 16828 36708 16884 37662
rect 16716 36652 16884 36708
rect 13580 36596 13636 36606
rect 13580 36502 13636 36540
rect 16380 36596 16436 36606
rect 16716 36596 16772 36652
rect 16380 36594 16772 36596
rect 16380 36542 16382 36594
rect 16434 36542 16772 36594
rect 16380 36540 16772 36542
rect 13468 36484 13524 36494
rect 13468 36390 13524 36428
rect 13020 35858 13076 35868
rect 14140 36034 14196 36046
rect 14140 35982 14142 36034
rect 14194 35982 14196 36034
rect 14140 35924 14196 35982
rect 14140 35858 14196 35868
rect 15260 35924 15316 35934
rect 11340 35758 11342 35810
rect 11394 35758 11396 35810
rect 11340 35746 11396 35758
rect 11900 35810 11956 35822
rect 11900 35758 11902 35810
rect 11954 35758 11956 35810
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 5628 35140 5684 35150
rect 5628 35046 5684 35084
rect 6300 35140 6356 35150
rect 4172 34626 4228 34636
rect 3724 34580 3780 34590
rect 3332 33964 3444 34020
rect 3276 33926 3332 33964
rect 3388 31780 3444 33964
rect 3724 34018 3780 34524
rect 5740 34580 5796 34590
rect 5740 34486 5796 34524
rect 3724 33966 3726 34018
rect 3778 33966 3780 34018
rect 3724 33954 3780 33966
rect 4060 34020 4116 34030
rect 4060 33926 4116 33964
rect 5740 33796 5796 33806
rect 4476 33292 4740 33302
rect 4532 33236 4580 33292
rect 4636 33236 4684 33292
rect 4476 33226 4740 33236
rect 5740 33122 5796 33740
rect 6300 33794 6356 35084
rect 11900 35140 11956 35758
rect 14476 35586 14532 35598
rect 14476 35534 14478 35586
rect 14530 35534 14532 35586
rect 11900 35074 11956 35084
rect 13468 35140 13524 35150
rect 13468 35046 13524 35084
rect 13580 34578 13636 34590
rect 13580 34526 13582 34578
rect 13634 34526 13636 34578
rect 13580 34020 13636 34526
rect 14476 34020 14532 35534
rect 13580 33964 14532 34020
rect 11900 33908 11956 33918
rect 11900 33906 12964 33908
rect 11900 33854 11902 33906
rect 11954 33854 12964 33906
rect 11900 33852 12964 33854
rect 11900 33842 11956 33852
rect 6300 33742 6302 33794
rect 6354 33742 6356 33794
rect 6300 33730 6356 33742
rect 6412 33796 6468 33806
rect 5740 33070 5742 33122
rect 5794 33070 5796 33122
rect 5740 33058 5796 33070
rect 3836 32564 3892 32574
rect 3836 31890 3892 32508
rect 5628 32564 5684 32574
rect 5628 32470 5684 32508
rect 6076 32562 6132 32574
rect 6076 32510 6078 32562
rect 6130 32510 6132 32562
rect 3836 31838 3838 31890
rect 3890 31838 3892 31890
rect 3836 31826 3892 31838
rect 4172 32002 4228 32014
rect 4172 31950 4174 32002
rect 4226 31950 4228 32002
rect 3388 31686 3444 31724
rect 4172 31780 4228 31950
rect 1820 30772 1876 30782
rect 1820 30770 1988 30772
rect 1820 30718 1822 30770
rect 1874 30718 1988 30770
rect 1820 30716 1988 30718
rect 1820 30706 1876 30716
rect 1820 29988 1876 29998
rect 1708 29932 1820 29988
rect 1708 27860 1764 29932
rect 1820 29894 1876 29932
rect 1820 28754 1876 28766
rect 1820 28702 1822 28754
rect 1874 28702 1876 28754
rect 1820 28082 1876 28702
rect 1932 28532 1988 30716
rect 2380 30770 2436 30782
rect 2380 30718 2382 30770
rect 2434 30718 2436 30770
rect 2380 30660 2436 30718
rect 2380 30594 2436 30604
rect 3724 30772 3780 30782
rect 2828 29988 2884 29998
rect 2828 29894 2884 29932
rect 3724 29986 3780 30716
rect 3724 29934 3726 29986
rect 3778 29934 3780 29986
rect 3724 29922 3780 29934
rect 4060 30548 4116 30558
rect 4172 30548 4228 31724
rect 4476 31276 4740 31286
rect 4532 31220 4580 31276
rect 4636 31220 4684 31276
rect 4476 31210 4740 31220
rect 5628 30770 5684 30782
rect 5628 30718 5630 30770
rect 5682 30718 5684 30770
rect 5516 30660 5572 30670
rect 5628 30660 5684 30718
rect 6076 30772 6132 32510
rect 6188 32450 6244 32462
rect 6188 32398 6190 32450
rect 6242 32398 6244 32450
rect 6188 31948 6244 32398
rect 6188 31892 6356 31948
rect 6300 31780 6356 31892
rect 6076 30706 6132 30716
rect 6188 31444 6244 31454
rect 6188 30770 6244 31388
rect 6188 30718 6190 30770
rect 6242 30718 6244 30770
rect 6188 30706 6244 30718
rect 5572 30604 5684 30660
rect 5516 30594 5572 30604
rect 4116 30492 4228 30548
rect 4620 30548 4676 30558
rect 4060 29988 4116 30492
rect 4620 30454 4676 30492
rect 4956 30546 5012 30558
rect 4956 30494 4958 30546
rect 5010 30494 5012 30546
rect 3276 29762 3332 29774
rect 3276 29710 3278 29762
rect 3330 29710 3332 29762
rect 3164 29426 3220 29438
rect 3164 29374 3166 29426
rect 3218 29374 3220 29426
rect 2380 28756 2436 28766
rect 2380 28662 2436 28700
rect 1932 28466 1988 28476
rect 3164 28532 3220 29374
rect 3164 28466 3220 28476
rect 1820 28030 1822 28082
rect 1874 28030 1876 28082
rect 1820 28018 1876 28030
rect 2380 28084 2436 28094
rect 2604 28084 2660 28094
rect 2380 28082 2660 28084
rect 2380 28030 2382 28082
rect 2434 28030 2606 28082
rect 2658 28030 2660 28082
rect 2380 28028 2660 28030
rect 1820 27860 1876 27870
rect 2268 27860 2324 27870
rect 1708 27858 2324 27860
rect 1708 27806 1822 27858
rect 1874 27806 2270 27858
rect 2322 27806 2324 27858
rect 1708 27804 2324 27806
rect 1708 25956 1764 27804
rect 1820 27794 1876 27804
rect 2268 27794 2324 27804
rect 1820 26740 1876 26750
rect 1820 26738 2324 26740
rect 1820 26686 1822 26738
rect 1874 26686 2324 26738
rect 1820 26684 2324 26686
rect 1820 26674 1876 26684
rect 1820 25956 1876 25966
rect 1708 25900 1820 25956
rect 1708 23940 1764 25900
rect 1820 25862 1876 25900
rect 2268 25620 2324 26684
rect 2380 26738 2436 28028
rect 2604 28018 2660 28028
rect 3164 27972 3220 27982
rect 3276 27972 3332 29710
rect 4060 28532 4116 29932
rect 4956 29540 5012 30494
rect 4956 29474 5012 29484
rect 4476 29260 4740 29270
rect 4532 29204 4580 29260
rect 4636 29204 4684 29260
rect 4476 29194 4740 29204
rect 5628 29090 5684 30604
rect 6300 29762 6356 31724
rect 6412 31778 6468 33740
rect 6860 33796 6916 33806
rect 6860 33702 6916 33740
rect 12124 33682 12180 33694
rect 12124 33630 12126 33682
rect 12178 33630 12180 33682
rect 9772 32788 9828 32798
rect 10108 32788 10164 32798
rect 9772 32786 10164 32788
rect 9772 32734 9774 32786
rect 9826 32734 10110 32786
rect 10162 32734 10164 32786
rect 9772 32732 10164 32734
rect 7532 32340 7588 32350
rect 6412 31726 6414 31778
rect 6466 31726 6468 31778
rect 6412 31714 6468 31726
rect 6972 31780 7028 31790
rect 6972 31686 7028 31724
rect 7420 31780 7476 31790
rect 7420 31686 7476 31724
rect 6300 29710 6302 29762
rect 6354 29710 6356 29762
rect 6300 29698 6356 29710
rect 6860 31444 6916 31454
rect 6860 29762 6916 31388
rect 7308 31444 7364 31454
rect 7308 31350 7364 31388
rect 7532 31444 7588 32284
rect 8876 32004 8932 32042
rect 8652 31892 8932 31948
rect 9772 32004 9828 32732
rect 10108 32722 10164 32732
rect 10892 32564 10948 32574
rect 10892 32470 10948 32508
rect 9772 31938 9828 31948
rect 9884 32002 9940 32014
rect 9884 31950 9886 32002
rect 9938 31950 9940 32002
rect 9884 31948 9940 31950
rect 12124 31948 12180 33630
rect 12236 33572 12292 33582
rect 12236 33478 12292 33516
rect 12908 33010 12964 33852
rect 12908 32958 12910 33010
rect 12962 32958 12964 33010
rect 9884 31892 10388 31948
rect 7532 31378 7588 31388
rect 8540 31668 8596 31678
rect 8652 31668 8708 31892
rect 10332 31890 10388 31892
rect 10332 31838 10334 31890
rect 10386 31838 10388 31890
rect 10332 31826 10388 31838
rect 10444 31890 10500 31902
rect 10444 31838 10446 31890
rect 10498 31838 10500 31890
rect 8540 31666 8708 31668
rect 8540 31614 8542 31666
rect 8594 31614 8708 31666
rect 8540 31612 8708 31614
rect 8764 31780 8820 31790
rect 8540 31108 8596 31612
rect 8316 31052 8596 31108
rect 7308 30548 7364 30558
rect 7308 29986 7364 30492
rect 7308 29934 7310 29986
rect 7362 29934 7364 29986
rect 7308 29922 7364 29934
rect 8316 30548 8372 31052
rect 8764 30994 8820 31724
rect 8988 31444 9044 31454
rect 8988 31442 9940 31444
rect 8988 31390 8990 31442
rect 9042 31390 9940 31442
rect 8988 31388 9940 31390
rect 8988 31378 9044 31388
rect 8764 30942 8766 30994
rect 8818 30942 8820 30994
rect 8764 30930 8820 30942
rect 9884 30770 9940 31388
rect 9884 30718 9886 30770
rect 9938 30718 9940 30770
rect 9884 30706 9940 30718
rect 9996 30996 10052 31006
rect 6860 29710 6862 29762
rect 6914 29710 6916 29762
rect 6860 29698 6916 29710
rect 5628 29038 5630 29090
rect 5682 29038 5684 29090
rect 5628 29026 5684 29038
rect 5740 29540 5796 29550
rect 5740 28754 5796 29484
rect 5740 28702 5742 28754
rect 5794 28702 5796 28754
rect 5740 28690 5796 28702
rect 6188 28756 6244 28766
rect 4956 28644 5012 28654
rect 4956 28550 5012 28588
rect 6076 28644 6132 28654
rect 6076 28550 6132 28588
rect 6188 28644 6244 28700
rect 6748 28756 6804 28766
rect 6188 28642 6356 28644
rect 6188 28590 6190 28642
rect 6242 28590 6356 28642
rect 6188 28588 6356 28590
rect 6188 28578 6244 28588
rect 4508 28532 4564 28542
rect 3164 27970 3332 27972
rect 3164 27918 3166 27970
rect 3218 27918 3332 27970
rect 3164 27916 3332 27918
rect 3612 28530 4564 28532
rect 3612 28478 4510 28530
rect 4562 28478 4564 28530
rect 3612 28476 4564 28478
rect 3612 27970 3668 28476
rect 3612 27918 3614 27970
rect 3666 27918 3668 27970
rect 3164 27906 3220 27916
rect 3612 27906 3668 27918
rect 2716 27746 2772 27758
rect 2716 27694 2718 27746
rect 2770 27694 2772 27746
rect 2716 26852 2772 27694
rect 2716 26786 2772 26796
rect 2380 26686 2382 26738
rect 2434 26686 2436 26738
rect 2380 26674 2436 26686
rect 4284 26516 4340 28476
rect 4508 28466 4564 28476
rect 5740 28532 5796 28542
rect 5740 27746 5796 28476
rect 5740 27694 5742 27746
rect 5794 27694 5796 27746
rect 5740 27682 5796 27694
rect 6300 27746 6356 28588
rect 6300 27694 6302 27746
rect 6354 27694 6356 27746
rect 6300 27682 6356 27694
rect 6748 27636 6804 28700
rect 6748 27570 6804 27580
rect 4476 27244 4740 27254
rect 4532 27188 4580 27244
rect 4636 27188 4684 27244
rect 4476 27178 4740 27188
rect 4956 26852 5012 26862
rect 4956 26758 5012 26796
rect 8316 26852 8372 30492
rect 9996 30100 10052 30940
rect 9996 30034 10052 30044
rect 10444 29650 10500 31838
rect 11788 31892 12292 31948
rect 10556 30548 10612 30558
rect 10556 30454 10612 30492
rect 11116 30548 11172 30558
rect 11116 29762 11172 30492
rect 11676 30436 11732 30446
rect 11564 30434 11732 30436
rect 11564 30382 11678 30434
rect 11730 30382 11732 30434
rect 11564 30380 11732 30382
rect 11564 29876 11620 30380
rect 11676 30370 11732 30380
rect 11676 30212 11732 30222
rect 11676 29986 11732 30156
rect 11788 30098 11844 31892
rect 12236 31890 12292 31892
rect 12236 31838 12238 31890
rect 12290 31838 12292 31890
rect 12236 31826 12292 31838
rect 12908 31892 12964 32958
rect 14028 33572 14084 33582
rect 14028 32786 14084 33516
rect 14028 32734 14030 32786
rect 14082 32734 14084 32786
rect 14028 32722 14084 32734
rect 13580 32676 13636 32686
rect 13468 32564 13524 32574
rect 13468 32470 13524 32508
rect 13580 32562 13636 32620
rect 13580 32510 13582 32562
rect 13634 32510 13636 32562
rect 13580 32498 13636 32510
rect 13916 32450 13972 32462
rect 13916 32398 13918 32450
rect 13970 32398 13972 32450
rect 13916 31948 13972 32398
rect 14140 32004 14196 32042
rect 12908 31826 12964 31836
rect 13804 31892 13860 31902
rect 13916 31892 14084 31948
rect 14140 31938 14196 31948
rect 14252 31948 14308 33964
rect 15260 32788 15316 35868
rect 16380 35924 16436 36540
rect 16380 35858 16436 35868
rect 16380 35700 16436 35710
rect 16380 35606 16436 35644
rect 16828 35698 16884 35710
rect 16828 35646 16830 35698
rect 16882 35646 16884 35698
rect 16828 35140 16884 35646
rect 16604 34692 16660 34702
rect 16604 34598 16660 34636
rect 16268 34578 16324 34590
rect 16268 34526 16270 34578
rect 16322 34526 16324 34578
rect 16268 33908 16324 34526
rect 16828 34018 16884 35084
rect 17276 35138 17332 40574
rect 18172 39956 18228 39966
rect 17724 39954 18228 39956
rect 17724 39902 18174 39954
rect 18226 39902 18228 39954
rect 17724 39900 18228 39902
rect 17500 39844 17556 39854
rect 17500 39842 17668 39844
rect 17500 39790 17502 39842
rect 17554 39790 17668 39842
rect 17500 39788 17668 39790
rect 17500 39778 17556 39788
rect 17612 38724 17668 39788
rect 17612 37826 17668 38668
rect 17612 37774 17614 37826
rect 17666 37774 17668 37826
rect 17612 37762 17668 37774
rect 17724 36146 17780 39900
rect 18172 39890 18228 39900
rect 17724 36094 17726 36146
rect 17778 36094 17780 36146
rect 17724 36082 17780 36094
rect 18172 37156 18228 37166
rect 18172 35924 18228 37100
rect 17276 35086 17278 35138
rect 17330 35086 17332 35138
rect 17276 35074 17332 35086
rect 17612 35922 18228 35924
rect 17612 35870 18174 35922
rect 18226 35870 18228 35922
rect 17612 35868 18228 35870
rect 17612 35698 17668 35868
rect 18172 35858 18228 35868
rect 17612 35646 17614 35698
rect 17666 35646 17668 35698
rect 17612 34916 17668 35646
rect 17724 35700 17780 35710
rect 17780 35644 17892 35700
rect 17724 35634 17780 35644
rect 16940 34860 17668 34916
rect 17724 35138 17780 35150
rect 17724 35086 17726 35138
rect 17778 35086 17780 35138
rect 16940 34356 16996 34860
rect 17724 34690 17780 35086
rect 17724 34638 17726 34690
rect 17778 34638 17780 34690
rect 17052 34580 17108 34590
rect 17724 34580 17780 34638
rect 17052 34578 17780 34580
rect 17052 34526 17054 34578
rect 17106 34526 17780 34578
rect 17052 34524 17780 34526
rect 17052 34514 17108 34524
rect 16940 34300 17220 34356
rect 16828 33966 16830 34018
rect 16882 33966 16884 34018
rect 16828 33954 16884 33966
rect 16380 33908 16436 33918
rect 16268 33852 16380 33908
rect 16380 33814 16436 33852
rect 16380 33684 16436 33694
rect 15708 32788 15764 32798
rect 15260 32786 15764 32788
rect 15260 32734 15262 32786
rect 15314 32734 15710 32786
rect 15762 32734 15764 32786
rect 15260 32732 15764 32734
rect 15260 32722 15316 32732
rect 14252 31892 14868 31948
rect 12908 31554 12964 31566
rect 12908 31502 12910 31554
rect 12962 31502 12964 31554
rect 12908 30884 12964 31502
rect 12460 30772 12516 30782
rect 12460 30678 12516 30716
rect 12124 30548 12180 30558
rect 12124 30454 12180 30492
rect 12908 30324 12964 30828
rect 13804 30660 13860 31836
rect 14028 30884 14084 31892
rect 14812 31890 14868 31892
rect 14812 31838 14814 31890
rect 14866 31838 14868 31890
rect 14812 31826 14868 31838
rect 15372 31892 15428 31902
rect 15372 31798 15428 31836
rect 15148 31778 15204 31790
rect 15148 31726 15150 31778
rect 15202 31726 15204 31778
rect 14364 31668 14420 31678
rect 14364 31574 14420 31612
rect 14924 30884 14980 30894
rect 14028 30828 14196 30884
rect 14028 30660 14084 30670
rect 13804 30658 14084 30660
rect 13804 30606 14030 30658
rect 14082 30606 14084 30658
rect 13804 30604 14084 30606
rect 12348 30268 12964 30324
rect 13244 30548 13300 30558
rect 11788 30046 11790 30098
rect 11842 30046 11844 30098
rect 11788 30034 11844 30046
rect 12124 30100 12180 30110
rect 12124 30006 12180 30044
rect 11676 29934 11678 29986
rect 11730 29934 11732 29986
rect 11676 29922 11732 29934
rect 11116 29710 11118 29762
rect 11170 29710 11172 29762
rect 11116 29698 11172 29710
rect 11228 29764 11284 29774
rect 11564 29764 11620 29820
rect 11228 29762 11620 29764
rect 11228 29710 11230 29762
rect 11282 29710 11620 29762
rect 11228 29708 11620 29710
rect 11228 29698 11284 29708
rect 10444 29598 10446 29650
rect 10498 29598 10500 29650
rect 10444 29586 10500 29598
rect 12348 28754 12404 30268
rect 12572 29876 12628 29886
rect 12572 29782 12628 29820
rect 13132 29874 13188 29886
rect 13132 29822 13134 29874
rect 13186 29822 13188 29874
rect 13132 29204 13188 29822
rect 13244 29874 13300 30492
rect 14028 30548 14084 30604
rect 14028 30482 14084 30492
rect 14140 30324 14196 30828
rect 14924 30790 14980 30828
rect 14700 30658 14756 30670
rect 14700 30606 14702 30658
rect 14754 30606 14756 30658
rect 14364 30548 14420 30558
rect 14700 30548 14756 30606
rect 14364 30546 14532 30548
rect 14364 30494 14366 30546
rect 14418 30494 14532 30546
rect 14364 30492 14532 30494
rect 14364 30482 14420 30492
rect 14140 30258 14196 30268
rect 13244 29822 13246 29874
rect 13298 29822 13300 29874
rect 13244 29810 13300 29822
rect 14364 29762 14420 29774
rect 14364 29710 14366 29762
rect 14418 29710 14420 29762
rect 13132 29138 13188 29148
rect 13916 29426 13972 29438
rect 13916 29374 13918 29426
rect 13970 29374 13972 29426
rect 12348 28702 12350 28754
rect 12402 28702 12404 28754
rect 12348 28690 12404 28702
rect 12908 29092 12964 29102
rect 12908 28754 12964 29036
rect 12908 28702 12910 28754
rect 12962 28702 12964 28754
rect 12908 28690 12964 28702
rect 12236 28644 12292 28654
rect 11564 28642 12292 28644
rect 11564 28590 12238 28642
rect 12290 28590 12292 28642
rect 11564 28588 12292 28590
rect 11564 27746 11620 28588
rect 12236 28578 12292 28588
rect 12460 28644 12516 28654
rect 12124 27748 12180 27758
rect 12460 27748 12516 28588
rect 13468 28644 13524 28654
rect 13692 28644 13748 28654
rect 13468 28550 13524 28588
rect 13580 28588 13692 28644
rect 13580 28530 13636 28588
rect 13692 28578 13748 28588
rect 13580 28478 13582 28530
rect 13634 28478 13636 28530
rect 13580 28466 13636 28478
rect 11564 27694 11566 27746
rect 11618 27694 11620 27746
rect 11564 27682 11620 27694
rect 11788 27746 12516 27748
rect 11788 27694 12126 27746
rect 12178 27694 12516 27746
rect 11788 27692 12516 27694
rect 12796 28418 12852 28430
rect 12796 28366 12798 28418
rect 12850 28366 12852 28418
rect 11228 27634 11284 27646
rect 11228 27582 11230 27634
rect 11282 27582 11284 27634
rect 8316 26786 8372 26796
rect 9324 26852 9380 26862
rect 10108 26852 10164 26862
rect 9380 26796 9604 26852
rect 9324 26758 9380 26796
rect 4508 26516 4564 26526
rect 4284 26514 5012 26516
rect 4284 26462 4510 26514
rect 4562 26462 5012 26514
rect 4284 26460 5012 26462
rect 4508 26450 4564 26460
rect 2716 25956 2772 25966
rect 2716 25862 2772 25900
rect 4956 25956 5012 26460
rect 4956 25954 5124 25956
rect 4956 25902 4958 25954
rect 5010 25902 5124 25954
rect 4956 25900 5124 25902
rect 4956 25890 5012 25900
rect 1820 25396 1876 25406
rect 1820 24724 1876 25340
rect 2268 24724 2324 25564
rect 3052 25730 3108 25742
rect 3052 25678 3054 25730
rect 3106 25678 3108 25730
rect 2380 24724 2436 24734
rect 1820 24722 2212 24724
rect 1820 24670 1822 24722
rect 1874 24670 2212 24722
rect 1820 24668 2212 24670
rect 2268 24722 2436 24724
rect 2268 24670 2382 24722
rect 2434 24670 2436 24722
rect 2268 24668 2436 24670
rect 1820 24658 1876 24668
rect 1820 23940 1876 23950
rect 1708 23884 1820 23940
rect 1708 21812 1764 23884
rect 1820 23846 1876 23884
rect 1932 23604 1988 23614
rect 1820 22708 1876 22718
rect 1932 22708 1988 23548
rect 1820 22706 1988 22708
rect 1820 22654 1822 22706
rect 1874 22654 1988 22706
rect 1820 22652 1988 22654
rect 2156 22708 2212 24668
rect 2380 24658 2436 24668
rect 2492 24388 2548 24398
rect 2268 24386 2548 24388
rect 2268 24334 2494 24386
rect 2546 24334 2548 24386
rect 2268 24332 2548 24334
rect 2268 23938 2324 24332
rect 2492 24322 2548 24332
rect 3052 24386 3108 25678
rect 3612 25732 3668 25742
rect 4060 25732 4116 25742
rect 3612 25730 3892 25732
rect 3612 25678 3614 25730
rect 3666 25678 3892 25730
rect 3612 25676 3892 25678
rect 3612 25666 3668 25676
rect 3052 24334 3054 24386
rect 3106 24334 3108 24386
rect 3052 24322 3108 24334
rect 3164 25394 3220 25406
rect 3164 25342 3166 25394
rect 3218 25342 3220 25394
rect 2268 23886 2270 23938
rect 2322 23886 2324 23938
rect 2268 23874 2324 23886
rect 2604 23940 2660 23950
rect 2604 23846 2660 23884
rect 3164 23604 3220 25342
rect 3500 25396 3556 25406
rect 3500 25302 3556 25340
rect 3836 24164 3892 25676
rect 4060 25730 5012 25732
rect 4060 25678 4062 25730
rect 4114 25678 5012 25730
rect 4060 25676 5012 25678
rect 4060 25666 4116 25676
rect 3948 25620 4004 25630
rect 3948 25526 4004 25564
rect 4620 25508 4676 25518
rect 4620 25506 4900 25508
rect 4620 25454 4622 25506
rect 4674 25454 4900 25506
rect 4620 25452 4900 25454
rect 4620 25442 4676 25452
rect 4476 25228 4740 25238
rect 4532 25172 4580 25228
rect 4636 25172 4684 25228
rect 4476 25162 4740 25172
rect 4844 24724 4900 25452
rect 4956 24946 5012 25676
rect 4956 24894 4958 24946
rect 5010 24894 5012 24946
rect 4956 24882 5012 24894
rect 4844 24658 4900 24668
rect 4620 24500 4676 24510
rect 5068 24500 5124 25900
rect 5740 25732 5796 25742
rect 5740 25060 5796 25676
rect 7196 25732 7252 25742
rect 7196 25638 7252 25676
rect 7756 25730 7812 25742
rect 7756 25678 7758 25730
rect 7810 25678 7812 25730
rect 6188 25620 6244 25630
rect 4620 24498 5068 24500
rect 4620 24446 4622 24498
rect 4674 24446 5068 24498
rect 4620 24444 5068 24446
rect 4620 24434 4676 24444
rect 5068 24406 5124 24444
rect 5404 25058 5796 25060
rect 5404 25006 5742 25058
rect 5794 25006 5796 25058
rect 5404 25004 5796 25006
rect 3836 24108 5012 24164
rect 3164 23538 3220 23548
rect 4844 23714 4900 23726
rect 4844 23662 4846 23714
rect 4898 23662 4900 23714
rect 4844 23604 4900 23662
rect 4844 23538 4900 23548
rect 4476 23212 4740 23222
rect 4532 23156 4580 23212
rect 4636 23156 4684 23212
rect 4476 23146 4740 23156
rect 4956 22930 5012 24108
rect 5404 23714 5460 25004
rect 5740 24994 5796 25004
rect 5852 25284 5908 25294
rect 5628 24724 5684 24734
rect 5628 24630 5684 24668
rect 5852 23938 5908 25228
rect 6188 24946 6244 25564
rect 7756 25396 7812 25678
rect 8204 25730 8260 25742
rect 8204 25678 8206 25730
rect 8258 25678 8260 25730
rect 8092 25396 8148 25406
rect 7756 25394 8148 25396
rect 7756 25342 8094 25394
rect 8146 25342 8148 25394
rect 7756 25340 8148 25342
rect 6188 24894 6190 24946
rect 6242 24894 6244 24946
rect 6188 24882 6244 24894
rect 5852 23886 5854 23938
rect 5906 23886 5908 23938
rect 5852 23874 5908 23886
rect 6188 24500 6244 24510
rect 6188 23938 6244 24444
rect 6524 24500 6580 24510
rect 6524 24406 6580 24444
rect 6188 23886 6190 23938
rect 6242 23886 6244 23938
rect 5404 23662 5406 23714
rect 5458 23662 5460 23714
rect 5404 23650 5460 23662
rect 4956 22878 4958 22930
rect 5010 22878 5012 22930
rect 4956 22866 5012 22878
rect 4620 22820 4676 22830
rect 2380 22708 2436 22718
rect 2156 22706 2436 22708
rect 2156 22654 2382 22706
rect 2434 22654 2436 22706
rect 2156 22652 2436 22654
rect 1820 22642 1876 22652
rect 2380 22642 2436 22652
rect 4620 22482 4676 22764
rect 5740 22820 5796 22830
rect 6188 22820 6244 23886
rect 8092 23716 8148 25340
rect 8204 25284 8260 25678
rect 8764 25732 8820 25742
rect 8764 25638 8820 25676
rect 8204 25218 8260 25228
rect 8876 25394 8932 25406
rect 8876 25342 8878 25394
rect 8930 25342 8932 25394
rect 8764 24724 8820 24734
rect 8876 24724 8932 25342
rect 9324 24724 9380 24734
rect 8764 24722 9044 24724
rect 8764 24670 8766 24722
rect 8818 24670 9044 24722
rect 8764 24668 9044 24670
rect 8764 24658 8820 24668
rect 8428 23716 8484 23726
rect 8092 23714 8484 23716
rect 8092 23662 8430 23714
rect 8482 23662 8484 23714
rect 8092 23660 8484 23662
rect 8428 23650 8484 23660
rect 8988 23714 9044 24668
rect 9324 24630 9380 24668
rect 9548 24500 9604 26796
rect 9772 26628 9828 26638
rect 9772 26534 9828 26572
rect 10108 26516 10164 26796
rect 11228 26852 11284 27582
rect 11228 26786 11284 26796
rect 11452 26628 11508 26638
rect 10108 26514 10612 26516
rect 10108 26462 10110 26514
rect 10162 26462 10612 26514
rect 10108 26460 10612 26462
rect 10108 26450 10164 26460
rect 10556 25954 10612 26460
rect 10556 25902 10558 25954
rect 10610 25902 10612 25954
rect 10556 25890 10612 25902
rect 11004 26404 11060 26414
rect 11004 25954 11060 26348
rect 11004 25902 11006 25954
rect 11058 25902 11060 25954
rect 11004 25890 11060 25902
rect 11452 25954 11508 26572
rect 11452 25902 11454 25954
rect 11506 25902 11508 25954
rect 11452 25890 11508 25902
rect 11788 25730 11844 27692
rect 12124 27682 12180 27692
rect 12796 26852 12852 28366
rect 13916 28308 13972 29374
rect 14028 28756 14084 28766
rect 14028 28662 14084 28700
rect 13916 28242 13972 28252
rect 14252 27970 14308 27982
rect 14252 27918 14254 27970
rect 14306 27918 14308 27970
rect 12460 26796 12796 26852
rect 12348 26740 12404 26750
rect 11788 25678 11790 25730
rect 11842 25678 11844 25730
rect 11788 25666 11844 25678
rect 12236 26738 12404 26740
rect 12236 26686 12350 26738
rect 12402 26686 12404 26738
rect 12236 26684 12404 26686
rect 9660 25396 9716 25406
rect 9660 24722 9716 25340
rect 10892 25394 10948 25406
rect 10892 25342 10894 25394
rect 10946 25342 10948 25394
rect 9660 24670 9662 24722
rect 9714 24670 9716 24722
rect 9660 24658 9716 24670
rect 10220 24724 10276 24734
rect 10220 24630 10276 24668
rect 10892 24724 10948 25342
rect 11340 25396 11396 25406
rect 11340 25302 11396 25340
rect 12124 25396 12180 25406
rect 12236 25396 12292 26684
rect 12348 26674 12404 26684
rect 12348 25732 12404 25742
rect 12460 25732 12516 26796
rect 12796 26786 12852 26796
rect 13468 26852 13524 26862
rect 12908 26740 12964 26750
rect 12348 25730 12516 25732
rect 12348 25678 12350 25730
rect 12402 25678 12516 25730
rect 12348 25676 12516 25678
rect 12796 26404 12852 26414
rect 12348 25666 12404 25676
rect 12180 25340 12292 25396
rect 12124 25330 12180 25340
rect 12796 24946 12852 26348
rect 12908 25956 12964 26684
rect 13468 26738 13524 26796
rect 13468 26686 13470 26738
rect 13522 26686 13524 26738
rect 13468 26674 13524 26686
rect 14028 26740 14084 26750
rect 14028 26646 14084 26684
rect 14252 26740 14308 27918
rect 13580 26516 13636 26526
rect 12908 25900 13524 25956
rect 13468 25058 13524 25900
rect 13468 25006 13470 25058
rect 13522 25006 13524 25058
rect 13468 24994 13524 25006
rect 12796 24894 12798 24946
rect 12850 24894 12852 24946
rect 12796 24882 12852 24894
rect 10892 24658 10948 24668
rect 13580 24722 13636 26460
rect 14252 25956 14308 26684
rect 14364 26404 14420 29710
rect 14476 29652 14532 30492
rect 14700 30482 14756 30492
rect 15036 30434 15092 30446
rect 15036 30382 15038 30434
rect 15090 30382 15092 30434
rect 15036 30100 15092 30382
rect 15036 30034 15092 30044
rect 14924 29876 14980 29886
rect 14924 29782 14980 29820
rect 15036 29652 15092 29662
rect 15148 29652 15204 31726
rect 15708 31780 15764 32732
rect 16380 32674 16436 33628
rect 16380 32622 16382 32674
rect 16434 32622 16436 32674
rect 16380 32610 16436 32622
rect 16940 33012 16996 33022
rect 16940 32002 16996 32956
rect 16940 31950 16942 32002
rect 16994 31950 16996 32002
rect 16940 31938 16996 31950
rect 15708 31714 15764 31724
rect 16380 31780 16436 31790
rect 16380 31686 16436 31724
rect 16268 30436 16324 30446
rect 15932 30100 15988 30110
rect 15932 29762 15988 30044
rect 16268 29986 16324 30380
rect 16268 29934 16270 29986
rect 16322 29934 16324 29986
rect 16268 29922 16324 29934
rect 15932 29710 15934 29762
rect 15986 29710 15988 29762
rect 15932 29698 15988 29710
rect 16156 29874 16212 29886
rect 16156 29822 16158 29874
rect 16210 29822 16212 29874
rect 14476 29650 15204 29652
rect 14476 29598 15038 29650
rect 15090 29598 15204 29650
rect 14476 29596 15204 29598
rect 15036 29586 15092 29596
rect 14924 29092 14980 29102
rect 14476 28642 14532 28654
rect 14476 28590 14478 28642
rect 14530 28590 14532 28642
rect 14476 26628 14532 28590
rect 14700 28644 14756 28654
rect 14700 27970 14756 28588
rect 14700 27918 14702 27970
rect 14754 27918 14756 27970
rect 14700 27906 14756 27918
rect 14476 26562 14532 26572
rect 14364 26338 14420 26348
rect 14588 25956 14644 25966
rect 14252 25954 14644 25956
rect 14252 25902 14590 25954
rect 14642 25902 14644 25954
rect 14252 25900 14644 25902
rect 13580 24670 13582 24722
rect 13634 24670 13636 24722
rect 13580 24658 13636 24670
rect 9548 23940 9604 24444
rect 12348 24500 12404 24510
rect 12348 24406 12404 24444
rect 14028 24500 14084 24510
rect 14028 24406 14084 24444
rect 14588 24500 14644 25900
rect 14924 25954 14980 29036
rect 15148 28868 15204 29596
rect 15484 29652 15540 29662
rect 15484 29090 15540 29596
rect 15484 29038 15486 29090
rect 15538 29038 15540 29090
rect 15484 29026 15540 29038
rect 16156 28868 16212 29822
rect 16380 29764 16436 29774
rect 16380 29670 16436 29708
rect 16940 28980 16996 28990
rect 16940 28886 16996 28924
rect 16604 28868 16660 28878
rect 15148 28866 15764 28868
rect 15148 28814 15150 28866
rect 15202 28814 15764 28866
rect 15148 28812 15764 28814
rect 16156 28812 16604 28868
rect 15148 28802 15204 28812
rect 15036 28756 15092 28766
rect 15036 28642 15092 28700
rect 15036 28590 15038 28642
rect 15090 28590 15092 28642
rect 15036 28578 15092 28590
rect 15484 27746 15540 27758
rect 15484 27694 15486 27746
rect 15538 27694 15540 27746
rect 15036 27410 15092 27422
rect 15036 27358 15038 27410
rect 15090 27358 15092 27410
rect 15036 26964 15092 27358
rect 15036 26898 15092 26908
rect 15484 26516 15540 27694
rect 15708 27746 15764 28812
rect 16604 28774 16660 28812
rect 15932 28644 15988 28654
rect 15932 28550 15988 28588
rect 16492 28644 16548 28654
rect 16492 28550 16548 28588
rect 16044 27860 16100 27870
rect 16044 27766 16100 27804
rect 15708 27694 15710 27746
rect 15762 27694 15764 27746
rect 15708 27682 15764 27694
rect 15484 26450 15540 26460
rect 16156 26740 16212 26750
rect 16156 26514 16212 26684
rect 16156 26462 16158 26514
rect 16210 26462 16212 26514
rect 16156 26450 16212 26462
rect 16604 26516 16660 26526
rect 16604 26422 16660 26460
rect 14924 25902 14926 25954
rect 14978 25902 14980 25954
rect 14924 25890 14980 25902
rect 16828 25620 16884 25630
rect 16268 24724 16324 24734
rect 16268 24630 16324 24668
rect 16716 24724 16772 24734
rect 16828 24724 16884 25564
rect 16716 24722 16884 24724
rect 16716 24670 16718 24722
rect 16770 24670 16884 24722
rect 16716 24668 16884 24670
rect 14588 24434 14644 24444
rect 9660 23940 9716 23950
rect 9548 23938 9716 23940
rect 9548 23886 9662 23938
rect 9714 23886 9716 23938
rect 9548 23884 9716 23886
rect 9660 23874 9716 23884
rect 8988 23662 8990 23714
rect 9042 23662 9044 23714
rect 8988 23650 9044 23662
rect 16716 23604 16772 24668
rect 16828 23604 16884 23614
rect 16716 23548 16828 23604
rect 16828 23510 16884 23548
rect 5796 22818 6244 22820
rect 5796 22766 6190 22818
rect 6242 22766 6244 22818
rect 5796 22764 6244 22766
rect 5740 22726 5796 22764
rect 6188 22754 6244 22764
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 4620 22418 4676 22430
rect 15708 22594 15764 22606
rect 15708 22542 15710 22594
rect 15762 22542 15764 22594
rect 15260 22372 15316 22382
rect 15260 22278 15316 22316
rect 15708 21924 15764 22542
rect 16268 22594 16324 22606
rect 16268 22542 16270 22594
rect 16322 22542 16324 22594
rect 15820 21924 15876 21934
rect 15708 21922 15876 21924
rect 15708 21870 15822 21922
rect 15874 21870 15876 21922
rect 15708 21868 15876 21870
rect 15820 21858 15876 21868
rect 1820 21812 1876 21822
rect 2268 21812 2324 21822
rect 1708 21810 2324 21812
rect 1708 21758 1822 21810
rect 1874 21758 2270 21810
rect 2322 21758 2324 21810
rect 1708 21756 2324 21758
rect 1820 21746 1876 21756
rect 2268 21746 2324 21756
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 16268 20804 16324 22542
rect 16380 22596 16436 22606
rect 16940 22596 16996 22606
rect 16380 22594 16996 22596
rect 16380 22542 16382 22594
rect 16434 22542 16942 22594
rect 16994 22542 16996 22594
rect 16380 22540 16996 22542
rect 16380 22530 16436 22540
rect 16940 21924 16996 22540
rect 16940 21858 16996 21868
rect 16380 21700 16436 21710
rect 16828 21700 16884 21710
rect 16380 21698 16884 21700
rect 16380 21646 16382 21698
rect 16434 21646 16830 21698
rect 16882 21646 16884 21698
rect 16380 21644 16884 21646
rect 16380 21634 16436 21644
rect 16268 20738 16324 20748
rect 14700 20690 14756 20702
rect 14700 20638 14702 20690
rect 14754 20638 14756 20690
rect 14700 20244 14756 20638
rect 15260 20244 15316 20254
rect 14700 20178 14756 20188
rect 15148 20132 15316 20188
rect 16828 20244 16884 21644
rect 16940 20804 16996 20814
rect 16940 20710 16996 20748
rect 4476 19180 4740 19190
rect 4532 19124 4580 19180
rect 4636 19124 4684 19180
rect 4476 19114 4740 19124
rect 15148 18674 15204 20132
rect 16716 19908 16772 19918
rect 16716 19814 16772 19852
rect 15148 18622 15150 18674
rect 15202 18622 15204 18674
rect 15148 18610 15204 18622
rect 16828 19682 16884 20188
rect 17164 20188 17220 34300
rect 17724 33908 17780 34524
rect 17500 33852 17780 33908
rect 17388 31780 17444 31790
rect 17388 29652 17444 31724
rect 17388 29586 17444 29596
rect 17388 29092 17444 29102
rect 17388 28754 17444 29036
rect 17388 28702 17390 28754
rect 17442 28702 17444 28754
rect 17388 28690 17444 28702
rect 17500 25956 17556 33852
rect 17836 33796 17892 35644
rect 18172 35140 18228 35150
rect 18284 35140 18340 40796
rect 19292 40852 19348 40862
rect 19292 40758 19348 40796
rect 19836 40348 20100 40358
rect 19892 40292 19940 40348
rect 19996 40292 20044 40348
rect 19836 40282 20100 40292
rect 20188 40068 20244 40908
rect 20300 40962 20356 44046
rect 20636 44658 20692 44670
rect 20636 44606 20638 44658
rect 20690 44606 20692 44658
rect 20636 42868 20692 44606
rect 21756 44660 21812 45726
rect 21756 44594 21812 44604
rect 21868 44770 21924 46956
rect 22428 46900 22484 46910
rect 22092 46674 22148 46686
rect 22092 46622 22094 46674
rect 22146 46622 22148 46674
rect 22092 46562 22148 46622
rect 22092 46510 22094 46562
rect 22146 46510 22148 46562
rect 22092 46498 22148 46510
rect 22428 46562 22484 46844
rect 22428 46510 22430 46562
rect 22482 46510 22484 46562
rect 22428 46498 22484 46510
rect 22652 46116 22708 48636
rect 23100 48130 23156 48748
rect 23100 48078 23102 48130
rect 23154 48078 23156 48130
rect 23100 48066 23156 48078
rect 23660 48802 23716 48814
rect 23660 48750 23662 48802
rect 23714 48750 23716 48802
rect 23548 47794 23604 47806
rect 23548 47742 23550 47794
rect 23602 47742 23604 47794
rect 22876 47012 22932 47022
rect 22876 46898 22932 46956
rect 23548 47012 23604 47742
rect 23660 47124 23716 48750
rect 23996 48804 24052 48814
rect 24332 48804 24388 48814
rect 23996 48802 24164 48804
rect 23996 48750 23998 48802
rect 24050 48750 24164 48802
rect 23996 48748 24164 48750
rect 23996 48738 24052 48748
rect 23660 47058 23716 47068
rect 23996 47794 24052 47806
rect 23996 47742 23998 47794
rect 24050 47742 24052 47794
rect 23548 46946 23604 46956
rect 22876 46846 22878 46898
rect 22930 46846 22932 46898
rect 22876 46834 22932 46846
rect 23996 46900 24052 47742
rect 23996 46834 24052 46844
rect 22652 46022 22708 46060
rect 23324 46116 23380 46126
rect 23324 46022 23380 46060
rect 23772 45778 23828 45790
rect 23772 45726 23774 45778
rect 23826 45726 23828 45778
rect 23772 45666 23828 45726
rect 23772 45614 23774 45666
rect 23826 45614 23828 45666
rect 23772 45602 23828 45614
rect 21868 44718 21870 44770
rect 21922 44718 21924 44770
rect 21196 44210 21252 44222
rect 21196 44158 21198 44210
rect 21250 44158 21252 44210
rect 21196 44098 21252 44158
rect 21196 44046 21198 44098
rect 21250 44046 21252 44098
rect 21196 44034 21252 44046
rect 21644 44100 21700 44110
rect 21868 44100 21924 44718
rect 21644 44098 21924 44100
rect 21644 44046 21646 44098
rect 21698 44046 21924 44098
rect 21644 44044 21924 44046
rect 23772 44660 23828 44670
rect 20636 42802 20692 42812
rect 20748 43762 20804 43774
rect 20748 43710 20750 43762
rect 20802 43710 20804 43762
rect 20748 43538 20804 43710
rect 21532 43764 21588 43774
rect 21644 43708 21700 44044
rect 21532 43652 21812 43708
rect 20748 43486 20750 43538
rect 20802 43486 20804 43538
rect 20412 42642 20468 42654
rect 20412 42590 20414 42642
rect 20466 42590 20468 42642
rect 20412 41748 20468 42590
rect 20468 41692 20580 41748
rect 20412 41682 20468 41692
rect 20300 40910 20302 40962
rect 20354 40910 20356 40962
rect 20300 40852 20356 40910
rect 20300 40786 20356 40796
rect 20412 41076 20468 41086
rect 20188 40002 20244 40012
rect 20188 39844 20244 39854
rect 20412 39844 20468 41020
rect 20188 39842 20468 39844
rect 20188 39790 20190 39842
rect 20242 39790 20468 39842
rect 20188 39788 20468 39790
rect 19852 38834 19908 38846
rect 19852 38782 19854 38834
rect 19906 38782 19908 38834
rect 19852 38724 19908 38782
rect 19852 38658 19908 38668
rect 19180 38612 19236 38622
rect 18844 38610 19236 38612
rect 18844 38558 19182 38610
rect 19234 38558 19236 38610
rect 18844 38556 19236 38558
rect 18396 37938 18452 37950
rect 18396 37886 18398 37938
rect 18450 37886 18452 37938
rect 18396 36148 18452 37886
rect 18732 36596 18788 36606
rect 18732 36502 18788 36540
rect 18844 36372 18900 38556
rect 19180 38546 19236 38556
rect 20188 38612 20244 39788
rect 20524 38668 20580 41692
rect 20748 41636 20804 43486
rect 21644 43538 21700 43550
rect 21644 43486 21646 43538
rect 21698 43486 21700 43538
rect 21644 42978 21700 43486
rect 21644 42926 21646 42978
rect 21698 42926 21700 42978
rect 21644 42914 21700 42926
rect 21644 41972 21700 41982
rect 21644 41878 21700 41916
rect 21756 41860 21812 43652
rect 23436 43652 23492 43662
rect 23100 42868 23156 42878
rect 23100 42774 23156 42812
rect 23436 42866 23492 43596
rect 23436 42814 23438 42866
rect 23490 42814 23492 42866
rect 23436 42802 23492 42814
rect 23772 42866 23828 44604
rect 24108 43652 24164 48748
rect 24332 48710 24388 48748
rect 25228 48804 25284 48814
rect 25228 48710 25284 48748
rect 25788 48804 25844 48814
rect 31948 48804 32004 48814
rect 25788 48802 25956 48804
rect 25788 48750 25790 48802
rect 25842 48750 25956 48802
rect 25788 48748 25956 48750
rect 25788 48738 25844 48748
rect 24668 48692 24724 48702
rect 24444 48690 24724 48692
rect 24444 48638 24670 48690
rect 24722 48638 24724 48690
rect 24444 48636 24724 48638
rect 24220 46900 24276 46910
rect 24220 46116 24276 46844
rect 24220 46022 24276 46060
rect 24220 44660 24276 44670
rect 24220 44658 24388 44660
rect 24220 44606 24222 44658
rect 24274 44606 24388 44658
rect 24220 44604 24388 44606
rect 24220 44594 24276 44604
rect 24108 43586 24164 43596
rect 24220 44210 24276 44222
rect 24220 44158 24222 44210
rect 24274 44158 24276 44210
rect 24220 44098 24276 44158
rect 24220 44046 24222 44098
rect 24274 44046 24276 44098
rect 23772 42814 23774 42866
rect 23826 42814 23828 42866
rect 23772 42802 23828 42814
rect 22092 42642 22148 42654
rect 22092 42590 22094 42642
rect 22146 42590 22148 42642
rect 21980 42196 22036 42206
rect 21868 41860 21924 41870
rect 21756 41804 21868 41860
rect 21868 41794 21924 41804
rect 20748 41570 20804 41580
rect 21980 41748 22036 42140
rect 21532 41524 21588 41534
rect 21532 41522 21700 41524
rect 21532 41470 21534 41522
rect 21586 41470 21700 41522
rect 21532 41468 21700 41470
rect 21532 41458 21588 41468
rect 21308 40852 21364 40862
rect 20748 40740 20804 40750
rect 20748 40646 20804 40684
rect 21308 40068 21364 40796
rect 21532 40738 21588 40750
rect 21532 40686 21534 40738
rect 21586 40686 21588 40738
rect 21308 40066 21476 40068
rect 21308 40014 21310 40066
rect 21362 40014 21476 40066
rect 21308 40012 21476 40014
rect 21308 40002 21364 40012
rect 20860 39956 20916 39966
rect 20860 39862 20916 39900
rect 21420 39732 21476 40012
rect 21532 39956 21588 40686
rect 21644 40068 21700 41468
rect 21868 40740 21924 40750
rect 21980 40740 22036 41692
rect 22092 41972 22148 42590
rect 24108 42642 24164 42654
rect 24108 42590 24110 42642
rect 24162 42590 24164 42642
rect 22092 41076 22148 41916
rect 22764 42196 22820 42206
rect 22764 41970 22820 42140
rect 22764 41918 22766 41970
rect 22818 41918 22820 41970
rect 22764 41906 22820 41918
rect 24108 41972 24164 42590
rect 24108 41906 24164 41916
rect 22092 41010 22148 41020
rect 22316 41860 22372 41870
rect 21868 40738 22036 40740
rect 21868 40686 21870 40738
rect 21922 40686 22036 40738
rect 21868 40684 22036 40686
rect 22316 40740 22372 41804
rect 22764 41636 22820 41646
rect 22764 40850 22820 41580
rect 22764 40798 22766 40850
rect 22818 40798 22820 40850
rect 22764 40786 22820 40798
rect 23884 41636 23940 41646
rect 21868 40674 21924 40684
rect 22316 40646 22372 40684
rect 23884 40404 23940 41580
rect 24220 40852 24276 44046
rect 24332 43876 24388 44604
rect 24332 43810 24388 43820
rect 24444 43708 24500 48636
rect 24668 48626 24724 48636
rect 25900 47010 25956 48748
rect 26460 48692 26516 48702
rect 26460 48690 27188 48692
rect 26460 48638 26462 48690
rect 26514 48638 27188 48690
rect 26460 48636 27188 48638
rect 26460 48626 26516 48636
rect 26460 48242 26516 48254
rect 26460 48190 26462 48242
rect 26514 48190 26516 48242
rect 26460 48130 26516 48190
rect 26460 48078 26462 48130
rect 26514 48078 26516 48130
rect 26460 48066 26516 48078
rect 26012 48020 26068 48030
rect 26012 47926 26068 47964
rect 25900 46958 25902 47010
rect 25954 46958 25956 47010
rect 25900 46946 25956 46958
rect 26908 47794 26964 47806
rect 26908 47742 26910 47794
rect 26962 47742 26964 47794
rect 26908 47012 26964 47742
rect 26908 46946 26964 46956
rect 27020 47570 27076 47582
rect 27020 47518 27022 47570
rect 27074 47518 27076 47570
rect 25116 46674 25172 46686
rect 25116 46622 25118 46674
rect 25170 46622 25172 46674
rect 24556 46228 24612 46238
rect 24556 44882 24612 46172
rect 25116 46228 25172 46622
rect 25116 46162 25172 46172
rect 26460 46228 26516 46238
rect 25452 46116 25508 46126
rect 25508 46060 25732 46116
rect 25452 46022 25508 46060
rect 25228 46002 25284 46014
rect 25228 45950 25230 46002
rect 25282 45950 25284 46002
rect 24556 44830 24558 44882
rect 24610 44830 24612 44882
rect 24556 44210 24612 44830
rect 24556 44158 24558 44210
rect 24610 44158 24612 44210
rect 24556 44146 24612 44158
rect 24668 45780 24724 45790
rect 25228 45780 25284 45950
rect 24668 45778 25228 45780
rect 24668 45726 24670 45778
rect 24722 45726 25228 45778
rect 24668 45724 25228 45726
rect 24668 45666 24724 45724
rect 25228 45686 25284 45724
rect 24668 45614 24670 45666
rect 24722 45614 24724 45666
rect 24220 40786 24276 40796
rect 24332 43652 24500 43708
rect 24668 44098 24724 45614
rect 24668 44046 24670 44098
rect 24722 44046 24724 44098
rect 24668 43708 24724 44046
rect 25340 44658 25396 44670
rect 25340 44606 25342 44658
rect 25394 44606 25396 44658
rect 24556 43652 24612 43662
rect 24668 43652 25172 43708
rect 21644 40002 21700 40012
rect 23660 40348 23940 40404
rect 23660 40066 23716 40348
rect 24108 40292 24164 40302
rect 23660 40014 23662 40066
rect 23714 40014 23716 40066
rect 21532 39890 21588 39900
rect 22540 39956 22596 39966
rect 22540 39862 22596 39900
rect 21644 39842 21700 39854
rect 21644 39790 21646 39842
rect 21698 39790 21700 39842
rect 21644 39732 21700 39790
rect 21420 39676 21700 39732
rect 19836 38332 20100 38342
rect 19892 38276 19940 38332
rect 19996 38276 20044 38332
rect 19836 38266 20100 38276
rect 20188 37156 20244 38556
rect 20188 37090 20244 37100
rect 20412 38612 20580 38668
rect 20636 38722 20692 38734
rect 20636 38670 20638 38722
rect 20690 38670 20692 38722
rect 20636 38612 20692 38670
rect 20412 37602 20468 38612
rect 20636 38546 20692 38556
rect 20860 38612 20916 38622
rect 20412 37550 20414 37602
rect 20466 37550 20468 37602
rect 20188 36932 20244 36942
rect 20188 36838 20244 36876
rect 19516 36818 19572 36830
rect 19516 36766 19518 36818
rect 19570 36766 19572 36818
rect 19516 36708 19572 36766
rect 19516 36642 19572 36652
rect 20412 36596 20468 37550
rect 20860 38050 20916 38556
rect 20860 37998 20862 38050
rect 20914 37998 20916 38050
rect 20748 36820 20804 36830
rect 20636 36596 20692 36606
rect 20412 36594 20692 36596
rect 20412 36542 20638 36594
rect 20690 36542 20692 36594
rect 20412 36540 20692 36542
rect 18396 36082 18452 36092
rect 18732 36316 18900 36372
rect 19836 36316 20100 36326
rect 18620 35922 18676 35934
rect 18620 35870 18622 35922
rect 18674 35870 18676 35922
rect 18620 35700 18676 35870
rect 18620 35634 18676 35644
rect 18172 35138 18340 35140
rect 18172 35086 18174 35138
rect 18226 35086 18340 35138
rect 18172 35084 18340 35086
rect 18732 35138 18788 36316
rect 19892 36260 19940 36316
rect 19996 36260 20044 36316
rect 19836 36250 20100 36260
rect 19180 36148 19236 36158
rect 19180 36054 19236 36092
rect 19628 36148 19684 36158
rect 18732 35086 18734 35138
rect 18786 35086 18788 35138
rect 18172 35074 18228 35084
rect 18732 35074 18788 35086
rect 18844 36036 18900 36046
rect 18844 35922 18900 35980
rect 18844 35870 18846 35922
rect 18898 35870 18900 35922
rect 18396 34916 18452 34926
rect 18844 34916 18900 35870
rect 19628 35810 19684 36092
rect 20636 36148 20692 36540
rect 20636 36082 20692 36092
rect 20748 36146 20804 36764
rect 20860 36708 20916 37998
rect 21644 38052 21700 39676
rect 23660 38836 23716 40014
rect 23660 38770 23716 38780
rect 23772 40068 23828 40078
rect 23772 38834 23828 40012
rect 23772 38782 23774 38834
rect 23826 38782 23828 38834
rect 23772 38770 23828 38782
rect 24108 38834 24164 40236
rect 24108 38782 24110 38834
rect 24162 38782 24164 38834
rect 24108 38770 24164 38782
rect 21644 37986 21700 37996
rect 23100 38052 23156 38062
rect 23100 37958 23156 37996
rect 23772 38052 23828 38062
rect 23828 37996 23940 38052
rect 23772 37958 23828 37996
rect 21420 37716 21476 37726
rect 21868 37716 21924 37726
rect 21420 37714 21588 37716
rect 21420 37662 21422 37714
rect 21474 37662 21588 37714
rect 21420 37660 21588 37662
rect 21420 37650 21476 37660
rect 20860 36642 20916 36652
rect 21196 36596 21252 36606
rect 21196 36502 21252 36540
rect 20748 36094 20750 36146
rect 20802 36094 20804 36146
rect 19628 35758 19630 35810
rect 19682 35758 19684 35810
rect 19628 35140 19684 35758
rect 18396 34914 18900 34916
rect 18396 34862 18398 34914
rect 18450 34862 18900 34914
rect 18396 34860 18900 34862
rect 19292 35084 19684 35140
rect 19852 36036 19908 36046
rect 18396 34850 18452 34860
rect 18172 34690 18228 34702
rect 18172 34638 18174 34690
rect 18226 34638 18228 34690
rect 18172 33908 18228 34638
rect 19180 34690 19236 34702
rect 19180 34638 19182 34690
rect 19234 34638 19236 34690
rect 18172 33842 18228 33852
rect 18844 33908 18900 33918
rect 18844 33814 18900 33852
rect 17724 33740 17892 33796
rect 18284 33794 18340 33806
rect 18284 33742 18286 33794
rect 18338 33742 18340 33794
rect 17724 33682 17780 33740
rect 17948 33684 18004 33694
rect 17724 33630 17726 33682
rect 17778 33630 17780 33682
rect 17724 33618 17780 33630
rect 17836 33628 17948 33684
rect 17836 33570 17892 33628
rect 17948 33618 18004 33628
rect 17836 33518 17838 33570
rect 17890 33518 17892 33570
rect 17836 33506 17892 33518
rect 18284 32564 18340 33742
rect 19180 33796 19236 34638
rect 18956 33684 19012 33694
rect 18956 33590 19012 33628
rect 18396 32786 18452 32798
rect 18396 32734 18398 32786
rect 18450 32734 18452 32786
rect 18396 32564 18452 32734
rect 18060 32508 18452 32564
rect 19068 32674 19124 32686
rect 19068 32622 19070 32674
rect 19122 32622 19124 32674
rect 17724 32004 17780 32014
rect 17612 30658 17668 30670
rect 17612 30606 17614 30658
rect 17666 30606 17668 30658
rect 17612 28980 17668 30606
rect 17612 28914 17668 28924
rect 17724 28868 17780 31948
rect 17948 30772 18004 30782
rect 18060 30772 18116 32508
rect 18620 32452 18676 32462
rect 18172 32450 18676 32452
rect 18172 32398 18622 32450
rect 18674 32398 18676 32450
rect 18172 32396 18676 32398
rect 18172 32002 18228 32396
rect 18620 32386 18676 32396
rect 18172 31950 18174 32002
rect 18226 31950 18228 32002
rect 18172 31938 18228 31950
rect 19068 31668 19124 32622
rect 17948 30770 18116 30772
rect 17948 30718 17950 30770
rect 18002 30718 18116 30770
rect 17948 30716 18116 30718
rect 18620 30772 18676 30782
rect 17948 30706 18004 30716
rect 18620 30678 18676 30716
rect 18284 30658 18340 30670
rect 18284 30606 18286 30658
rect 18338 30606 18340 30658
rect 18284 29764 18340 30606
rect 19068 30658 19124 31612
rect 19068 30606 19070 30658
rect 19122 30606 19124 30658
rect 19068 30594 19124 30606
rect 19180 30436 19236 33740
rect 19068 30380 19236 30436
rect 18284 29708 18788 29764
rect 18060 29652 18116 29662
rect 18060 29558 18116 29596
rect 17724 28754 17780 28812
rect 17724 28702 17726 28754
rect 17778 28702 17780 28754
rect 17724 28690 17780 28702
rect 18396 29538 18452 29550
rect 18396 29486 18398 29538
rect 18450 29486 18452 29538
rect 18396 28756 18452 29486
rect 18732 29090 18788 29708
rect 18732 29038 18734 29090
rect 18786 29038 18788 29090
rect 18732 29026 18788 29038
rect 18396 28690 18452 28700
rect 18508 28980 18564 28990
rect 17948 28642 18004 28654
rect 17948 28590 17950 28642
rect 18002 28590 18004 28642
rect 17948 28084 18004 28590
rect 17948 28018 18004 28028
rect 18508 28082 18564 28924
rect 18508 28030 18510 28082
rect 18562 28030 18564 28082
rect 18508 28018 18564 28030
rect 18956 28420 19012 28430
rect 18956 27860 19012 28364
rect 18956 27766 19012 27804
rect 17500 25900 17668 25956
rect 17500 25730 17556 25742
rect 17500 25678 17502 25730
rect 17554 25678 17556 25730
rect 17500 24724 17556 25678
rect 17500 23716 17556 24668
rect 17612 24836 17668 25900
rect 17836 25730 17892 25742
rect 17836 25678 17838 25730
rect 17890 25678 17892 25730
rect 17836 25620 17892 25678
rect 17836 25554 17892 25564
rect 17612 23826 17668 24780
rect 17612 23774 17614 23826
rect 17666 23774 17668 23826
rect 17612 23762 17668 23774
rect 17948 24724 18004 24734
rect 17500 23650 17556 23660
rect 17948 23714 18004 24668
rect 19068 24724 19124 30380
rect 19180 29204 19236 29214
rect 19180 28642 19236 29148
rect 19180 28590 19182 28642
rect 19234 28590 19236 28642
rect 19180 28532 19236 28590
rect 19180 28466 19236 28476
rect 19068 23940 19124 24668
rect 18956 23884 19068 23940
rect 18508 23716 18564 23726
rect 17948 23662 17950 23714
rect 18002 23662 18004 23714
rect 17948 23650 18004 23662
rect 18396 23714 18564 23716
rect 18396 23662 18510 23714
rect 18562 23662 18564 23714
rect 18396 23660 18564 23662
rect 18396 23604 18452 23660
rect 18508 23650 18564 23660
rect 18844 23716 18900 23726
rect 18844 23622 18900 23660
rect 18396 22596 18452 23548
rect 17836 22540 18396 22596
rect 17836 21810 17892 22540
rect 18396 22530 18452 22540
rect 17836 21758 17838 21810
rect 17890 21758 17892 21810
rect 17836 21746 17892 21758
rect 17948 21924 18004 21934
rect 17948 21476 18004 21868
rect 18284 21924 18340 21934
rect 18956 21924 19012 23884
rect 19068 23874 19124 23884
rect 18284 21830 18340 21868
rect 18844 21868 19012 21924
rect 18620 21812 18676 21822
rect 18620 21718 18676 21756
rect 17164 20132 17668 20188
rect 16828 19630 16830 19682
rect 16882 19630 16884 19682
rect 16828 17892 16884 19630
rect 16828 17890 17556 17892
rect 16828 17838 16830 17890
rect 16882 17838 17556 17890
rect 16828 17836 17556 17838
rect 16828 17826 16884 17836
rect 4476 17164 4740 17174
rect 4532 17108 4580 17164
rect 4636 17108 4684 17164
rect 4476 17098 4740 17108
rect 4476 15148 4740 15158
rect 4532 15092 4580 15148
rect 4636 15092 4684 15148
rect 4476 15082 4740 15092
rect 17500 14644 17556 17836
rect 17612 15652 17668 20132
rect 17724 19794 17780 19806
rect 17724 19742 17726 19794
rect 17778 19742 17780 19794
rect 17724 18788 17780 19742
rect 17948 19682 18004 21420
rect 18172 19908 18228 19918
rect 18172 19794 18228 19852
rect 18172 19742 18174 19794
rect 18226 19742 18228 19794
rect 18172 19730 18228 19742
rect 17948 19630 17950 19682
rect 18002 19630 18004 19682
rect 17948 19618 18004 19630
rect 18844 19684 18900 21868
rect 19180 21812 19236 21822
rect 19180 20802 19236 21756
rect 19180 20750 19182 20802
rect 19234 20750 19236 20802
rect 19180 20468 19236 20750
rect 19180 20402 19236 20412
rect 18956 19684 19012 19694
rect 18844 19682 19012 19684
rect 18844 19630 18958 19682
rect 19010 19630 19012 19682
rect 18844 19628 19012 19630
rect 18620 19348 18676 19358
rect 18620 19254 18676 19292
rect 17836 18788 17892 18798
rect 17724 18786 17892 18788
rect 17724 18734 17838 18786
rect 17890 18734 17892 18786
rect 17724 18732 17892 18734
rect 17836 18722 17892 18732
rect 17724 17668 17780 17678
rect 17724 17666 17892 17668
rect 17724 17614 17726 17666
rect 17778 17614 17892 17666
rect 17724 17612 17892 17614
rect 17724 17602 17780 17612
rect 17724 15652 17780 15662
rect 17612 15596 17724 15652
rect 17724 15558 17780 15596
rect 17836 14756 17892 17612
rect 18732 17556 18788 17566
rect 18956 17556 19012 19628
rect 19292 19684 19348 35084
rect 19852 34914 19908 35980
rect 20748 36036 20804 36094
rect 20748 35970 20804 35980
rect 19852 34862 19854 34914
rect 19906 34862 19908 34914
rect 19852 34850 19908 34862
rect 20188 35922 20244 35934
rect 20188 35870 20190 35922
rect 20242 35870 20244 35922
rect 20188 35140 20244 35870
rect 20300 35812 20356 35822
rect 21084 35812 21140 35822
rect 20300 35810 21140 35812
rect 20300 35758 20302 35810
rect 20354 35758 21086 35810
rect 21138 35758 21140 35810
rect 20300 35756 21140 35758
rect 20300 35746 20356 35756
rect 19628 34692 19684 34702
rect 19628 34020 19684 34636
rect 19836 34300 20100 34310
rect 19892 34244 19940 34300
rect 19996 34244 20044 34300
rect 19836 34234 20100 34244
rect 19852 34020 19908 34030
rect 19628 34018 19908 34020
rect 19628 33966 19854 34018
rect 19906 33966 19908 34018
rect 19628 33964 19908 33966
rect 19852 33954 19908 33964
rect 20188 34020 20244 35084
rect 20748 35028 20804 35038
rect 20860 35028 20916 35756
rect 21084 35746 21140 35756
rect 21420 35700 21476 35710
rect 21420 35140 21476 35644
rect 21532 35700 21588 37660
rect 21868 37714 22036 37716
rect 21868 37662 21870 37714
rect 21922 37662 22036 37714
rect 21868 37660 22036 37662
rect 21868 37650 21924 37660
rect 21644 36932 21700 36942
rect 21644 36818 21700 36876
rect 21644 36766 21646 36818
rect 21698 36766 21700 36818
rect 21644 36754 21700 36766
rect 21868 36820 21924 36830
rect 21868 36726 21924 36764
rect 21980 36708 22036 37660
rect 23100 36932 23156 36942
rect 23100 36838 23156 36876
rect 23884 36818 23940 37996
rect 24220 37716 24276 37726
rect 24220 36932 24276 37660
rect 24220 36838 24276 36876
rect 23884 36766 23886 36818
rect 23938 36766 23940 36818
rect 23884 36754 23940 36766
rect 22092 36708 22148 36718
rect 21980 36706 22148 36708
rect 21980 36654 22094 36706
rect 22146 36654 22148 36706
rect 21980 36652 22148 36654
rect 21868 36596 21924 36606
rect 21868 35810 21924 36540
rect 21868 35758 21870 35810
rect 21922 35758 21924 35810
rect 21868 35746 21924 35758
rect 21532 35698 21700 35700
rect 21532 35646 21534 35698
rect 21586 35646 21700 35698
rect 21532 35644 21700 35646
rect 21532 35634 21588 35644
rect 21420 35084 21588 35140
rect 20524 35026 21140 35028
rect 20524 34974 20750 35026
rect 20802 34974 21140 35026
rect 20524 34972 21140 34974
rect 20412 34804 20468 34814
rect 20412 34710 20468 34748
rect 20188 33954 20244 33964
rect 20188 33796 20244 33806
rect 20188 33702 20244 33740
rect 19740 33684 19796 33694
rect 19516 33012 19572 33022
rect 19516 32674 19572 32956
rect 19740 32898 19796 33628
rect 19740 32846 19742 32898
rect 19794 32846 19796 32898
rect 19740 32834 19796 32846
rect 19516 32622 19518 32674
rect 19570 32622 19572 32674
rect 19516 32610 19572 32622
rect 20188 32786 20244 32798
rect 20188 32734 20190 32786
rect 20242 32734 20244 32786
rect 19836 32284 20100 32294
rect 19892 32228 19940 32284
rect 19996 32228 20044 32284
rect 19836 32218 20100 32228
rect 20188 32004 20244 32734
rect 20300 32676 20356 32686
rect 20300 32582 20356 32620
rect 20412 32676 20468 32686
rect 20524 32676 20580 34972
rect 20748 34962 20804 34972
rect 21084 34244 21140 34972
rect 21420 34914 21476 34926
rect 21420 34862 21422 34914
rect 21474 34862 21476 34914
rect 21308 34802 21364 34814
rect 21308 34750 21310 34802
rect 21362 34750 21364 34802
rect 21308 34692 21364 34750
rect 21308 34626 21364 34636
rect 21084 34188 21364 34244
rect 20860 34020 20916 34030
rect 20860 33926 20916 33964
rect 20972 33908 21028 33918
rect 20972 33814 21028 33852
rect 21308 33906 21364 34188
rect 21308 33854 21310 33906
rect 21362 33854 21364 33906
rect 21308 33842 21364 33854
rect 21420 33684 21476 34862
rect 21532 34804 21588 35084
rect 21532 34710 21588 34748
rect 21644 34916 21700 35644
rect 21644 33796 21700 34860
rect 21980 34916 22036 34926
rect 21756 34690 21812 34702
rect 21756 34638 21758 34690
rect 21810 34638 21812 34690
rect 21756 34020 21812 34638
rect 21980 34690 22036 34860
rect 21980 34638 21982 34690
rect 22034 34638 22036 34690
rect 21812 33964 21924 34020
rect 21756 33954 21812 33964
rect 21644 33740 21812 33796
rect 20636 32788 20692 32798
rect 20636 32694 20692 32732
rect 20412 32674 20580 32676
rect 20412 32622 20414 32674
rect 20466 32622 20580 32674
rect 20412 32620 20580 32622
rect 20412 32610 20468 32620
rect 20188 31938 20244 31948
rect 19516 31892 19572 31902
rect 19516 29876 19572 31836
rect 21308 31890 21364 31902
rect 21308 31838 21310 31890
rect 21362 31838 21364 31890
rect 20860 31780 20916 31790
rect 20636 31778 20916 31780
rect 20636 31726 20862 31778
rect 20914 31726 20916 31778
rect 20636 31724 20916 31726
rect 20188 31668 20244 31678
rect 20188 31574 20244 31612
rect 20412 31444 20468 31454
rect 20412 31442 20580 31444
rect 20412 31390 20414 31442
rect 20466 31390 20580 31442
rect 20412 31388 20580 31390
rect 20412 31378 20468 31388
rect 19740 30660 19796 30670
rect 19628 30658 19796 30660
rect 19628 30606 19742 30658
rect 19794 30606 19796 30658
rect 19628 30604 19796 30606
rect 19628 30100 19684 30604
rect 19740 30594 19796 30604
rect 20412 30548 20468 30558
rect 20412 30454 20468 30492
rect 19836 30268 20100 30278
rect 19892 30212 19940 30268
rect 19996 30212 20044 30268
rect 19836 30202 20100 30212
rect 19628 30034 19684 30044
rect 20412 29988 20468 29998
rect 20524 29988 20580 31388
rect 20412 29986 20580 29988
rect 20412 29934 20414 29986
rect 20466 29934 20580 29986
rect 20412 29932 20580 29934
rect 20412 29922 20468 29932
rect 19516 29820 19684 29876
rect 19628 29204 19684 29820
rect 19516 28756 19572 28766
rect 19404 28084 19460 28094
rect 19404 27858 19460 28028
rect 19404 27806 19406 27858
rect 19458 27806 19460 27858
rect 19404 27412 19460 27806
rect 19516 27746 19572 28700
rect 19628 28642 19684 29148
rect 19852 28980 19908 28990
rect 19852 28866 19908 28924
rect 20636 28980 20692 31724
rect 20860 31714 20916 31724
rect 21308 31444 21364 31838
rect 21420 31778 21476 33628
rect 21644 33572 21700 33582
rect 21644 33478 21700 33516
rect 21756 32898 21812 33740
rect 21756 32846 21758 32898
rect 21810 32846 21812 32898
rect 21756 32834 21812 32846
rect 21868 32788 21924 33964
rect 21980 33906 22036 34638
rect 21980 33854 21982 33906
rect 22034 33854 22036 33906
rect 21980 33842 22036 33854
rect 22092 33012 22148 36652
rect 23548 36596 23604 36606
rect 23548 36502 23604 36540
rect 23996 36596 24052 36606
rect 23884 35924 23940 35934
rect 23436 35922 23940 35924
rect 23436 35870 23886 35922
rect 23938 35870 23940 35922
rect 23436 35868 23940 35870
rect 22876 34804 22932 34814
rect 22876 34710 22932 34748
rect 23324 34804 23380 34814
rect 23324 34710 23380 34748
rect 22428 34692 22484 34702
rect 22428 34598 22484 34636
rect 22316 34578 22372 34590
rect 22316 34526 22318 34578
rect 22370 34526 22372 34578
rect 22316 34356 22372 34526
rect 22204 33796 22260 33806
rect 22316 33796 22372 34300
rect 22764 34578 22820 34590
rect 22764 34526 22766 34578
rect 22818 34526 22820 34578
rect 22764 34132 22820 34526
rect 22540 34076 22820 34132
rect 23212 34132 23268 34142
rect 22204 33794 22372 33796
rect 22204 33742 22206 33794
rect 22258 33742 22372 33794
rect 22204 33740 22372 33742
rect 22428 33908 22484 33918
rect 22540 33908 22596 34076
rect 22428 33906 22596 33908
rect 22428 33854 22430 33906
rect 22482 33854 22596 33906
rect 22428 33852 22596 33854
rect 22652 33908 22708 33918
rect 22204 33730 22260 33740
rect 22092 32946 22148 32956
rect 22204 33570 22260 33582
rect 22204 33518 22206 33570
rect 22258 33518 22260 33570
rect 22092 32788 22148 32798
rect 21868 32786 22148 32788
rect 21868 32734 22094 32786
rect 22146 32734 22148 32786
rect 21868 32732 22148 32734
rect 22092 32722 22148 32732
rect 22204 32788 22260 33518
rect 22204 32722 22260 32732
rect 22428 32564 22484 33852
rect 22652 33814 22708 33852
rect 23212 33684 23268 34076
rect 23436 34130 23492 35868
rect 23884 35858 23940 35868
rect 23772 34692 23828 34702
rect 23772 34598 23828 34636
rect 23436 34078 23438 34130
rect 23490 34078 23492 34130
rect 23436 34066 23492 34078
rect 23660 33908 23716 33918
rect 22428 32498 22484 32508
rect 23100 33682 23268 33684
rect 23100 33630 23214 33682
rect 23266 33630 23268 33682
rect 23100 33628 23268 33630
rect 21420 31726 21422 31778
rect 21474 31726 21476 31778
rect 21420 31714 21476 31726
rect 22876 31892 22932 31902
rect 21308 31378 21364 31388
rect 22204 31666 22260 31678
rect 22204 31614 22206 31666
rect 22258 31614 22260 31666
rect 22204 31444 22260 31614
rect 22204 31378 22260 31388
rect 22876 30884 22932 31836
rect 22988 31444 23044 31454
rect 23100 31444 23156 33628
rect 23212 33618 23268 33628
rect 23548 33684 23604 33694
rect 23548 32786 23604 33628
rect 23548 32734 23550 32786
rect 23602 32734 23604 32786
rect 23548 32722 23604 32734
rect 23660 32674 23716 33852
rect 23884 33908 23940 33918
rect 23996 33908 24052 36540
rect 24332 34244 24388 43652
rect 24556 40292 24612 43596
rect 24668 43428 24724 43438
rect 24668 42866 24724 43372
rect 24668 42814 24670 42866
rect 24722 42814 24724 42866
rect 24668 42802 24724 42814
rect 25116 41972 25172 43652
rect 25228 42868 25284 42878
rect 25340 42868 25396 44606
rect 25228 42866 25396 42868
rect 25228 42814 25230 42866
rect 25282 42814 25396 42866
rect 25228 42812 25396 42814
rect 25676 44098 25732 46060
rect 26460 46114 26516 46172
rect 26460 46062 26462 46114
rect 26514 46062 26516 46114
rect 26460 46050 26516 46062
rect 25676 44046 25678 44098
rect 25730 44046 25732 44098
rect 25676 43764 25732 44046
rect 26012 44658 26068 44670
rect 26012 44606 26014 44658
rect 26066 44606 26068 44658
rect 26012 43708 26068 44606
rect 27020 43876 27076 47518
rect 27132 46116 27188 48636
rect 27244 48242 27300 48254
rect 27244 48190 27246 48242
rect 27298 48190 27300 48242
rect 27244 47122 27300 48190
rect 27692 48242 27748 48254
rect 27692 48190 27694 48242
rect 27746 48190 27748 48242
rect 27692 47906 27748 48190
rect 27692 47854 27694 47906
rect 27746 47854 27748 47906
rect 27692 47842 27748 47854
rect 28140 48020 28196 48030
rect 27356 47794 27412 47806
rect 27356 47742 27358 47794
rect 27410 47742 27412 47794
rect 27356 47570 27412 47742
rect 27356 47518 27358 47570
rect 27410 47518 27412 47570
rect 27356 47506 27412 47518
rect 27244 47070 27246 47122
rect 27298 47070 27300 47122
rect 27244 47010 27300 47070
rect 27244 46958 27246 47010
rect 27298 46958 27300 47010
rect 27244 46946 27300 46958
rect 27804 47122 27860 47134
rect 27804 47070 27806 47122
rect 27858 47070 27860 47122
rect 27692 46674 27748 46686
rect 27692 46622 27694 46674
rect 27746 46622 27748 46674
rect 27356 46228 27412 46238
rect 27244 46116 27300 46126
rect 27132 46114 27300 46116
rect 27132 46062 27246 46114
rect 27298 46062 27300 46114
rect 27132 46060 27300 46062
rect 27244 46050 27300 46060
rect 25228 42802 25284 42812
rect 25340 41972 25396 41982
rect 25116 41970 25396 41972
rect 25116 41918 25342 41970
rect 25394 41918 25396 41970
rect 25116 41916 25396 41918
rect 25116 41860 25172 41916
rect 25116 41794 25172 41804
rect 24556 40226 24612 40236
rect 24668 41748 24724 41758
rect 24668 40066 24724 41692
rect 24668 40014 24670 40066
rect 24722 40014 24724 40066
rect 24668 39956 24724 40014
rect 24444 39732 24500 39742
rect 24444 38834 24500 39676
rect 24444 38782 24446 38834
rect 24498 38782 24500 38834
rect 24444 38770 24500 38782
rect 24668 37714 24724 39900
rect 24780 40404 24836 40414
rect 24780 38834 24836 40348
rect 24780 38782 24782 38834
rect 24834 38782 24836 38834
rect 24780 38770 24836 38782
rect 25228 38276 25284 41916
rect 25340 41906 25396 41916
rect 25564 41858 25620 41870
rect 25564 41806 25566 41858
rect 25618 41806 25620 41858
rect 25564 41636 25620 41806
rect 25676 41748 25732 43708
rect 25900 43652 26068 43708
rect 26124 43764 26180 43802
rect 26124 43698 26180 43708
rect 27020 43708 27076 43820
rect 27244 45780 27300 45790
rect 27244 44098 27300 45724
rect 27244 44046 27246 44098
rect 27298 44046 27300 44098
rect 27020 43652 27188 43708
rect 25900 42754 25956 43652
rect 27132 42980 27188 43652
rect 27244 43652 27300 44046
rect 27356 44882 27412 46172
rect 27692 46228 27748 46622
rect 27692 46162 27748 46172
rect 27356 44830 27358 44882
rect 27410 44830 27412 44882
rect 27356 43708 27412 44830
rect 27804 45890 27860 47070
rect 28140 47012 28196 47964
rect 28476 48020 28532 48030
rect 28476 47926 28532 47964
rect 31052 47682 31108 47694
rect 31052 47630 31054 47682
rect 31106 47630 31108 47682
rect 28476 47122 28532 47134
rect 28476 47070 28478 47122
rect 28530 47070 28532 47122
rect 28476 47012 28532 47070
rect 28588 47012 28644 47022
rect 28140 47010 28308 47012
rect 28140 46958 28142 47010
rect 28194 46958 28308 47010
rect 28140 46956 28308 46958
rect 28476 47010 28644 47012
rect 28476 46958 28590 47010
rect 28642 46958 28644 47010
rect 28476 46956 28644 46958
rect 28140 46946 28196 46956
rect 28252 46788 28308 46956
rect 28588 46900 28644 46956
rect 28588 46834 28644 46844
rect 29372 46900 29428 46910
rect 29372 46806 29428 46844
rect 29820 46898 29876 46910
rect 29820 46846 29822 46898
rect 29874 46846 29876 46898
rect 28252 46004 28308 46732
rect 29820 46788 29876 46846
rect 29820 46722 29876 46732
rect 30604 46228 30660 46238
rect 30604 46114 30660 46172
rect 30604 46062 30606 46114
rect 30658 46062 30660 46114
rect 30604 46050 30660 46062
rect 27804 45838 27806 45890
rect 27858 45838 27860 45890
rect 27804 44660 27860 45838
rect 27804 44594 27860 44604
rect 28140 46002 28308 46004
rect 28140 45950 28254 46002
rect 28306 45950 28308 46002
rect 28140 45948 28308 45950
rect 28140 44770 28196 45948
rect 28252 45938 28308 45948
rect 31052 46004 31108 47630
rect 31948 46452 32004 48748
rect 32508 48804 32564 48814
rect 33068 48804 33124 48814
rect 32508 48802 33124 48804
rect 32508 48750 32510 48802
rect 32562 48750 33070 48802
rect 33122 48750 33124 48802
rect 32508 48748 33124 48750
rect 32508 48738 32564 48748
rect 32060 47794 32116 47806
rect 32620 47796 32676 47806
rect 32060 47742 32062 47794
rect 32114 47742 32116 47794
rect 32060 47012 32116 47742
rect 32060 46676 32116 46956
rect 32508 47794 32676 47796
rect 32508 47742 32622 47794
rect 32674 47742 32676 47794
rect 32508 47740 32676 47742
rect 32172 46900 32228 46910
rect 32172 46898 32452 46900
rect 32172 46846 32174 46898
rect 32226 46846 32452 46898
rect 32172 46844 32452 46846
rect 32172 46834 32228 46844
rect 32060 46610 32116 46620
rect 31948 46396 32340 46452
rect 32284 46228 32340 46396
rect 32060 46172 32284 46228
rect 31052 45938 31108 45948
rect 31948 46116 32004 46126
rect 31948 46002 32004 46060
rect 31948 45950 31950 46002
rect 32002 45950 32004 46002
rect 31948 45938 32004 45950
rect 31500 45892 31556 45902
rect 31500 45798 31556 45836
rect 28140 44718 28142 44770
rect 28194 44718 28196 44770
rect 28028 43762 28084 43774
rect 28028 43710 28030 43762
rect 28082 43710 28084 43762
rect 27356 43652 27748 43708
rect 27244 43586 27300 43596
rect 27244 42980 27300 42990
rect 27132 42924 27244 42980
rect 27244 42886 27300 42924
rect 27692 42978 27748 43652
rect 27692 42926 27694 42978
rect 27746 42926 27748 42978
rect 27692 42914 27748 42926
rect 25900 42702 25902 42754
rect 25954 42702 25956 42754
rect 25900 42690 25956 42702
rect 28028 42868 28084 43710
rect 26796 42642 26852 42654
rect 26796 42590 26798 42642
rect 26850 42590 26852 42642
rect 26796 42196 26852 42590
rect 26796 42130 26852 42140
rect 27468 41972 27524 41982
rect 27468 41878 27524 41916
rect 27916 41970 27972 41982
rect 27916 41918 27918 41970
rect 27970 41918 27972 41970
rect 25676 41682 25732 41692
rect 26796 41858 26852 41870
rect 26796 41806 26798 41858
rect 26850 41806 26852 41858
rect 26796 41748 26852 41806
rect 27132 41860 27188 41870
rect 27132 41748 27188 41804
rect 26852 41692 27188 41748
rect 26796 41682 26852 41692
rect 25564 41570 25620 41580
rect 27020 41524 27076 41534
rect 26908 41522 27076 41524
rect 26908 41470 27022 41522
rect 27074 41470 27076 41522
rect 26908 41468 27076 41470
rect 25452 41076 25508 41086
rect 25452 40850 25508 41020
rect 25452 40798 25454 40850
rect 25506 40798 25508 40850
rect 25452 40786 25508 40798
rect 25788 40852 25844 40862
rect 25788 40758 25844 40796
rect 26572 40514 26628 40526
rect 26572 40462 26574 40514
rect 26626 40462 26628 40514
rect 26348 39956 26404 39966
rect 26348 39862 26404 39900
rect 25452 39732 25508 39742
rect 25452 39638 25508 39676
rect 25900 38836 25956 38846
rect 25900 38742 25956 38780
rect 25340 38724 25396 38734
rect 25340 38630 25396 38668
rect 26572 38722 26628 40462
rect 26572 38670 26574 38722
rect 26626 38670 26628 38722
rect 26572 38658 26628 38670
rect 25228 38220 25396 38276
rect 25228 38052 25284 38062
rect 25228 37938 25284 37996
rect 25228 37886 25230 37938
rect 25282 37886 25284 37938
rect 25228 37874 25284 37886
rect 25340 37828 25396 38220
rect 25564 37828 25620 37838
rect 25340 37826 25620 37828
rect 25340 37774 25566 37826
rect 25618 37774 25620 37826
rect 25340 37772 25620 37774
rect 24668 37662 24670 37714
rect 24722 37662 24724 37714
rect 24444 36708 24500 36718
rect 24444 35812 24500 36652
rect 24668 36596 24724 37662
rect 25564 37716 25620 37772
rect 25564 37650 25620 37660
rect 26012 36708 26068 36718
rect 26012 36614 26068 36652
rect 24668 36530 24724 36540
rect 25900 36596 25956 36606
rect 25900 35922 25956 36540
rect 25900 35870 25902 35922
rect 25954 35870 25956 35922
rect 25900 35858 25956 35870
rect 26460 36484 26516 36494
rect 26460 35922 26516 36428
rect 26460 35870 26462 35922
rect 26514 35870 26516 35922
rect 26460 35858 26516 35870
rect 24556 35812 24612 35822
rect 24444 35756 24556 35812
rect 24556 35718 24612 35756
rect 26348 35812 26404 35822
rect 25452 35476 25508 35486
rect 25116 35474 25508 35476
rect 25116 35422 25454 35474
rect 25506 35422 25508 35474
rect 25116 35420 25508 35422
rect 24892 34802 24948 34814
rect 24892 34750 24894 34802
rect 24946 34750 24948 34802
rect 24668 34580 24724 34590
rect 24332 34188 24612 34244
rect 24108 34132 24164 34142
rect 24164 34076 24388 34132
rect 24108 34066 24164 34076
rect 23884 33906 24052 33908
rect 23884 33854 23886 33906
rect 23938 33854 24052 33906
rect 23884 33852 24052 33854
rect 24332 33906 24388 34076
rect 24332 33854 24334 33906
rect 24386 33854 24388 33906
rect 23884 33842 23940 33852
rect 24332 33842 24388 33854
rect 24108 33794 24164 33806
rect 24108 33742 24110 33794
rect 24162 33742 24164 33794
rect 24108 33684 24164 33742
rect 24164 33628 24500 33684
rect 24108 33618 24164 33628
rect 24332 32788 24388 32798
rect 24332 32694 24388 32732
rect 24444 32786 24500 33628
rect 24556 32900 24612 34188
rect 24668 34132 24724 34524
rect 24668 34066 24724 34076
rect 24892 34020 24948 34750
rect 25116 34690 25172 35420
rect 25452 35410 25508 35420
rect 25676 35252 25732 35262
rect 25676 34802 25732 35196
rect 25676 34750 25678 34802
rect 25730 34750 25732 34802
rect 25676 34738 25732 34750
rect 25116 34638 25118 34690
rect 25170 34638 25172 34690
rect 25116 34626 25172 34638
rect 26012 34690 26068 34702
rect 26012 34638 26014 34690
rect 26066 34638 26068 34690
rect 24892 33954 24948 33964
rect 25228 34578 25284 34590
rect 25228 34526 25230 34578
rect 25282 34526 25284 34578
rect 25116 33794 25172 33806
rect 25116 33742 25118 33794
rect 25170 33742 25172 33794
rect 25116 33684 25172 33742
rect 25116 33618 25172 33628
rect 24556 32844 24836 32900
rect 24444 32734 24446 32786
rect 24498 32734 24500 32786
rect 24444 32722 24500 32734
rect 23660 32622 23662 32674
rect 23714 32622 23716 32674
rect 23660 32610 23716 32622
rect 23212 32564 23268 32574
rect 23212 32562 23380 32564
rect 23212 32510 23214 32562
rect 23266 32510 23380 32562
rect 23212 32508 23380 32510
rect 23212 32498 23268 32508
rect 23044 31388 23156 31444
rect 22988 31378 23044 31388
rect 22876 30882 23268 30884
rect 22876 30830 22878 30882
rect 22930 30830 23268 30882
rect 22876 30828 23268 30830
rect 22876 30818 22932 30828
rect 23212 30770 23268 30828
rect 23212 30718 23214 30770
rect 23266 30718 23268 30770
rect 23212 30706 23268 30718
rect 21420 30548 21476 30558
rect 21476 30492 21700 30548
rect 21420 30482 21476 30492
rect 21420 30100 21476 30110
rect 21420 30006 21476 30044
rect 21084 29762 21140 29774
rect 21084 29710 21086 29762
rect 21138 29710 21140 29762
rect 21084 29652 21140 29710
rect 21084 29586 21140 29596
rect 21196 29764 21252 29774
rect 20636 28886 20692 28924
rect 21196 29092 21252 29708
rect 19852 28814 19854 28866
rect 19906 28814 19908 28866
rect 19852 28802 19908 28814
rect 20300 28756 20356 28766
rect 21196 28756 21252 29036
rect 21644 29090 21700 30492
rect 21868 29876 21924 29886
rect 21868 29782 21924 29820
rect 22316 29874 22372 29886
rect 22316 29822 22318 29874
rect 22370 29822 22372 29874
rect 22092 29762 22148 29774
rect 22092 29710 22094 29762
rect 22146 29710 22148 29762
rect 21644 29038 21646 29090
rect 21698 29038 21700 29090
rect 21644 29026 21700 29038
rect 21756 29428 21812 29438
rect 21532 28980 21588 28990
rect 21308 28756 21364 28766
rect 21196 28754 21364 28756
rect 21196 28702 21310 28754
rect 21362 28702 21364 28754
rect 21196 28700 21364 28702
rect 20300 28662 20356 28700
rect 21308 28690 21364 28700
rect 19628 28590 19630 28642
rect 19682 28590 19684 28642
rect 19628 28578 19684 28590
rect 21532 28642 21588 28924
rect 21756 28754 21812 29372
rect 22092 28980 22148 29710
rect 22092 28914 22148 28924
rect 21756 28702 21758 28754
rect 21810 28702 21812 28754
rect 21756 28690 21812 28702
rect 22316 28868 22372 29822
rect 21532 28590 21534 28642
rect 21586 28590 21588 28642
rect 21532 28578 21588 28590
rect 22316 28308 22372 28812
rect 22988 29762 23044 29774
rect 22988 29710 22990 29762
rect 23042 29710 23044 29762
rect 22988 28756 23044 29710
rect 23100 29764 23156 29774
rect 23100 29670 23156 29708
rect 22988 28690 23044 28700
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 22316 28242 22372 28252
rect 19836 28186 20100 28196
rect 19516 27694 19518 27746
rect 19570 27694 19572 27746
rect 19516 27682 19572 27694
rect 19516 27412 19572 27422
rect 19404 27356 19516 27412
rect 19516 27346 19572 27356
rect 22204 26628 22260 26638
rect 20748 26516 20804 26526
rect 20636 26514 20804 26516
rect 20636 26462 20750 26514
rect 20802 26462 20804 26514
rect 20636 26460 20804 26462
rect 19836 26236 20100 26246
rect 19892 26180 19940 26236
rect 19996 26180 20044 26236
rect 19836 26170 20100 26180
rect 19964 25732 20020 25742
rect 19404 24836 19460 24846
rect 19964 24836 20020 25676
rect 20524 25284 20580 25294
rect 20524 24946 20580 25228
rect 20524 24894 20526 24946
rect 20578 24894 20580 24946
rect 20524 24882 20580 24894
rect 19460 24780 19684 24836
rect 19404 24742 19460 24780
rect 19628 22036 19684 24780
rect 19964 24770 20020 24780
rect 19836 24220 20100 24230
rect 19892 24164 19940 24220
rect 19996 24164 20044 24220
rect 19836 24154 20100 24164
rect 20300 23716 20356 23726
rect 20188 22596 20244 22606
rect 19836 22204 20100 22214
rect 19892 22148 19940 22204
rect 19996 22148 20044 22204
rect 19836 22138 20100 22148
rect 19628 21980 19908 22036
rect 19852 20804 19908 21980
rect 20188 20804 20244 22540
rect 20300 22482 20356 23660
rect 20636 22820 20692 26460
rect 20748 26450 20804 26460
rect 21420 26514 21476 26526
rect 21420 26462 21422 26514
rect 21474 26462 21476 26514
rect 20748 25732 20804 25742
rect 21196 25732 21252 25742
rect 20748 25730 21252 25732
rect 20748 25678 20750 25730
rect 20802 25678 21198 25730
rect 21250 25678 21252 25730
rect 20748 25676 21252 25678
rect 20748 25666 20804 25676
rect 21196 25666 21252 25676
rect 21420 25732 21476 26462
rect 21868 26514 21924 26526
rect 21868 26462 21870 26514
rect 21922 26462 21924 26514
rect 21868 26180 21924 26462
rect 21924 26124 22036 26180
rect 21868 26114 21924 26124
rect 21420 25666 21476 25676
rect 21532 25730 21588 25742
rect 21532 25678 21534 25730
rect 21586 25678 21588 25730
rect 21420 25396 21476 25406
rect 21308 25340 21420 25396
rect 21308 23940 21364 25340
rect 21420 25330 21476 25340
rect 21420 24948 21476 24958
rect 21420 24722 21476 24892
rect 21420 24670 21422 24722
rect 21474 24670 21476 24722
rect 21420 24658 21476 24670
rect 21420 23940 21476 23950
rect 21308 23938 21476 23940
rect 21308 23886 21422 23938
rect 21474 23886 21476 23938
rect 21308 23884 21476 23886
rect 21420 23874 21476 23884
rect 20748 22820 20804 22830
rect 20636 22818 20804 22820
rect 20636 22766 20750 22818
rect 20802 22766 20804 22818
rect 20636 22764 20804 22766
rect 20636 22596 20692 22764
rect 20748 22754 20804 22764
rect 20636 22530 20692 22540
rect 21308 22594 21364 22606
rect 21308 22542 21310 22594
rect 21362 22542 21364 22594
rect 20300 22430 20302 22482
rect 20354 22430 20356 22482
rect 20300 21700 20356 22430
rect 20524 21924 20580 21934
rect 21308 21924 21364 22542
rect 21532 22596 21588 25678
rect 21868 25730 21924 25742
rect 21868 25678 21870 25730
rect 21922 25678 21924 25730
rect 21868 25396 21924 25678
rect 21868 25330 21924 25340
rect 21980 24948 22036 26124
rect 22204 25954 22260 26572
rect 23324 26180 23380 32508
rect 23884 32562 23940 32574
rect 23884 32510 23886 32562
rect 23938 32510 23940 32562
rect 23884 30660 23940 32510
rect 24108 32562 24164 32574
rect 24108 32510 24110 32562
rect 24162 32510 24164 32562
rect 24108 31444 24164 32510
rect 24668 32564 24724 32574
rect 24668 32470 24724 32508
rect 24220 31892 24276 31902
rect 24220 31798 24276 31836
rect 24668 31780 24724 31790
rect 24668 31686 24724 31724
rect 24556 31444 24612 31454
rect 24108 31442 24612 31444
rect 24108 31390 24558 31442
rect 24610 31390 24612 31442
rect 24108 31388 24612 31390
rect 23996 30660 24052 30670
rect 23884 30658 24052 30660
rect 23884 30606 23998 30658
rect 24050 30606 24052 30658
rect 23884 30604 24052 30606
rect 23996 30594 24052 30604
rect 24220 30436 24276 30446
rect 24220 29762 24276 30380
rect 24556 30212 24612 31388
rect 24556 30146 24612 30156
rect 24220 29710 24222 29762
rect 24274 29710 24276 29762
rect 24108 29426 24164 29438
rect 24108 29374 24110 29426
rect 24162 29374 24164 29426
rect 24108 28644 24164 29374
rect 24220 28756 24276 29710
rect 24444 29988 24500 29998
rect 24444 29762 24500 29932
rect 24444 29710 24446 29762
rect 24498 29710 24500 29762
rect 24444 29698 24500 29710
rect 24668 29876 24724 29886
rect 24668 29762 24724 29820
rect 24668 29710 24670 29762
rect 24722 29710 24724 29762
rect 24668 29698 24724 29710
rect 24444 28756 24500 28766
rect 24220 28754 24500 28756
rect 24220 28702 24446 28754
rect 24498 28702 24500 28754
rect 24220 28700 24500 28702
rect 24444 28690 24500 28700
rect 24668 28754 24724 28766
rect 24668 28702 24670 28754
rect 24722 28702 24724 28754
rect 24108 28578 24164 28588
rect 24332 28532 24388 28542
rect 24332 28438 24388 28476
rect 24556 27748 24612 27758
rect 23436 27300 23492 27310
rect 23436 26850 23492 27244
rect 23436 26798 23438 26850
rect 23490 26798 23492 26850
rect 23436 26786 23492 26798
rect 24556 26850 24612 27692
rect 24668 27524 24724 28702
rect 24668 27458 24724 27468
rect 24556 26798 24558 26850
rect 24610 26798 24612 26850
rect 24556 26786 24612 26798
rect 23324 26114 23380 26124
rect 23548 26626 23604 26638
rect 23548 26574 23550 26626
rect 23602 26574 23604 26626
rect 22204 25902 22206 25954
rect 22258 25902 22260 25954
rect 22204 25890 22260 25902
rect 21980 24882 22036 24892
rect 22764 25730 22820 25742
rect 22764 25678 22766 25730
rect 22818 25678 22820 25730
rect 22764 25620 22820 25678
rect 21980 24724 22036 24734
rect 21980 24630 22036 24668
rect 22316 24500 22372 24510
rect 22092 24050 22148 24062
rect 22092 23998 22094 24050
rect 22146 23998 22148 24050
rect 22092 23940 22148 23998
rect 22092 23846 22148 23884
rect 21756 22708 21812 22718
rect 21644 22596 21700 22606
rect 21756 22596 21812 22652
rect 22316 22706 22372 24444
rect 22540 23604 22596 23614
rect 22540 23510 22596 23548
rect 22316 22654 22318 22706
rect 22370 22654 22372 22706
rect 22316 22642 22372 22654
rect 21532 22594 21812 22596
rect 21532 22542 21646 22594
rect 21698 22542 21812 22594
rect 21532 22540 21812 22542
rect 21980 22594 22036 22606
rect 21980 22542 21982 22594
rect 22034 22542 22036 22594
rect 21644 22530 21700 22540
rect 20524 21922 21364 21924
rect 20524 21870 20526 21922
rect 20578 21870 21364 21922
rect 20524 21868 21364 21870
rect 21980 21924 22036 22542
rect 22764 22594 22820 25564
rect 23324 25730 23380 25742
rect 23324 25678 23326 25730
rect 23378 25678 23380 25730
rect 23324 25284 23380 25678
rect 23324 25218 23380 25228
rect 22988 24948 23044 24958
rect 22988 24050 23044 24892
rect 23548 24500 23604 26574
rect 24108 26628 24164 26638
rect 24108 26534 24164 26572
rect 23996 25844 24052 25854
rect 23996 25842 24164 25844
rect 23996 25790 23998 25842
rect 24050 25790 24164 25842
rect 23996 25788 24164 25790
rect 23996 25778 24052 25788
rect 24108 24834 24164 25788
rect 24780 25396 24836 32844
rect 24892 32564 24948 32574
rect 24892 32470 24948 32508
rect 25116 32562 25172 32574
rect 25116 32510 25118 32562
rect 25170 32510 25172 32562
rect 25116 31108 25172 32510
rect 25228 32116 25284 34526
rect 25452 34578 25508 34590
rect 25452 34526 25454 34578
rect 25506 34526 25508 34578
rect 25340 34356 25396 34366
rect 25340 34018 25396 34300
rect 25340 33966 25342 34018
rect 25394 33966 25396 34018
rect 25340 33954 25396 33966
rect 25452 33908 25508 34526
rect 25788 33908 25844 33918
rect 25452 33852 25788 33908
rect 25788 33814 25844 33852
rect 26012 33796 26068 34638
rect 26124 34690 26180 34702
rect 26124 34638 26126 34690
rect 26178 34638 26180 34690
rect 26124 34580 26180 34638
rect 26124 34514 26180 34524
rect 26236 34020 26292 34030
rect 25900 33794 26068 33796
rect 25900 33742 26014 33794
rect 26066 33742 26068 33794
rect 25900 33740 26068 33742
rect 25564 33682 25620 33694
rect 25564 33630 25566 33682
rect 25618 33630 25620 33682
rect 25340 32788 25396 32798
rect 25340 32564 25396 32732
rect 25564 32788 25620 33630
rect 25900 33124 25956 33740
rect 26012 33730 26068 33740
rect 26124 33964 26236 34020
rect 25564 32722 25620 32732
rect 25676 33068 25956 33124
rect 25564 32564 25620 32574
rect 25676 32564 25732 33068
rect 25900 32900 25956 32910
rect 25900 32676 25956 32844
rect 25900 32582 25956 32620
rect 25340 32562 25732 32564
rect 25340 32510 25566 32562
rect 25618 32510 25732 32562
rect 25340 32508 25732 32510
rect 26012 32564 26068 32574
rect 25564 32498 25620 32508
rect 25228 32050 25284 32060
rect 26012 32002 26068 32508
rect 26012 31950 26014 32002
rect 26066 31950 26068 32002
rect 26012 31938 26068 31950
rect 25228 31892 25284 31902
rect 25228 31778 25284 31836
rect 25228 31726 25230 31778
rect 25282 31726 25284 31778
rect 25228 31714 25284 31726
rect 26012 31780 26068 31790
rect 25116 31042 25172 31052
rect 26012 30996 26068 31724
rect 26012 30902 26068 30940
rect 25788 30324 25844 30334
rect 25676 29986 25732 29998
rect 25676 29934 25678 29986
rect 25730 29934 25732 29986
rect 25676 29876 25732 29934
rect 25676 29650 25732 29820
rect 25676 29598 25678 29650
rect 25730 29598 25732 29650
rect 25676 29586 25732 29598
rect 25228 29428 25284 29438
rect 25228 29334 25284 29372
rect 24892 28754 24948 28766
rect 24892 28702 24894 28754
rect 24946 28702 24948 28754
rect 24892 28084 24948 28702
rect 25452 28756 25508 28766
rect 24892 28018 24948 28028
rect 25116 28642 25172 28654
rect 25116 28590 25118 28642
rect 25170 28590 25172 28642
rect 24780 25330 24836 25340
rect 24892 26514 24948 26526
rect 24892 26462 24894 26514
rect 24946 26462 24948 26514
rect 24108 24782 24110 24834
rect 24162 24782 24164 24834
rect 24108 24770 24164 24782
rect 24556 25172 24612 25182
rect 24108 24500 24164 24510
rect 23548 24434 23604 24444
rect 23772 24444 24108 24500
rect 22988 23998 22990 24050
rect 23042 23998 23044 24050
rect 22988 23938 23044 23998
rect 22988 23886 22990 23938
rect 23042 23886 23044 23938
rect 22988 23874 23044 23886
rect 23212 23940 23268 23950
rect 22764 22542 22766 22594
rect 22818 22542 22820 22594
rect 22764 22530 22820 22542
rect 22652 22034 22708 22046
rect 22652 21982 22654 22034
rect 22706 21982 22708 22034
rect 22092 21924 22148 21934
rect 21980 21922 22148 21924
rect 21980 21870 22094 21922
rect 22146 21870 22148 21922
rect 21980 21868 22148 21870
rect 20524 21858 20580 21868
rect 22092 21858 22148 21868
rect 20748 21700 20804 21710
rect 20300 21644 20748 21700
rect 20300 20804 20356 20814
rect 20188 20802 20356 20804
rect 20188 20750 20302 20802
rect 20354 20750 20356 20802
rect 20188 20748 20356 20750
rect 19852 20710 19908 20748
rect 20300 20580 20356 20748
rect 20188 20468 20244 20478
rect 19836 20188 20100 20198
rect 19892 20132 19940 20188
rect 19996 20132 20044 20188
rect 19836 20122 20100 20132
rect 19628 19796 19684 19806
rect 19628 19702 19684 19740
rect 19292 19590 19348 19628
rect 20188 19570 20244 20412
rect 20300 20188 20356 20524
rect 20748 20802 20804 21644
rect 21196 21700 21252 21710
rect 21196 21606 21252 21644
rect 20748 20750 20750 20802
rect 20802 20750 20804 20802
rect 20748 20468 20804 20750
rect 21420 20692 21476 20702
rect 21420 20598 21476 20636
rect 22540 20692 22596 20702
rect 20748 20402 20804 20412
rect 21644 20580 21700 20590
rect 21644 20188 21700 20524
rect 20300 20132 20804 20188
rect 21644 20132 21812 20188
rect 20300 19796 20356 20132
rect 20300 19730 20356 19740
rect 20188 19518 20190 19570
rect 20242 19518 20244 19570
rect 19836 18172 20100 18182
rect 19892 18116 19940 18172
rect 19996 18116 20044 18172
rect 19836 18106 20100 18116
rect 18732 17554 19012 17556
rect 18732 17502 18734 17554
rect 18786 17502 19012 17554
rect 18732 17500 19012 17502
rect 18732 16884 18788 17500
rect 18732 16818 18788 16828
rect 19516 16884 19572 16894
rect 19292 14866 19348 14878
rect 19292 14814 19294 14866
rect 19346 14814 19348 14866
rect 16828 13748 16884 13758
rect 16828 13654 16884 13692
rect 17500 13634 17556 14588
rect 17500 13582 17502 13634
rect 17554 13582 17556 13634
rect 17500 13570 17556 13582
rect 17612 14700 17836 14756
rect 4476 13132 4740 13142
rect 4532 13076 4580 13132
rect 4636 13076 4684 13132
rect 4476 13066 4740 13076
rect 17500 12628 17556 12638
rect 17612 12628 17668 14700
rect 17836 14690 17892 14700
rect 19180 14756 19236 14766
rect 19180 14662 19236 14700
rect 18396 14420 18452 14430
rect 18396 13758 18452 14364
rect 19180 13860 19236 13870
rect 19292 13860 19348 14814
rect 19180 13858 19348 13860
rect 19180 13806 19182 13858
rect 19234 13806 19348 13858
rect 19180 13804 19348 13806
rect 19180 13794 19236 13804
rect 18284 13748 18340 13758
rect 18396 13748 18461 13758
rect 18340 13746 18461 13748
rect 18340 13694 18407 13746
rect 18459 13694 18461 13746
rect 18340 13692 18461 13694
rect 18284 13682 18340 13692
rect 18405 13682 18461 13692
rect 19292 12850 19348 13804
rect 19516 13636 19572 16828
rect 20188 16772 20244 19518
rect 20748 18786 20804 20132
rect 20748 18734 20750 18786
rect 20802 18734 20804 18786
rect 20748 18722 20804 18734
rect 20300 16772 20356 16782
rect 20188 16770 20356 16772
rect 20188 16718 20302 16770
rect 20354 16718 20356 16770
rect 20188 16716 20356 16718
rect 21756 16772 21812 20132
rect 22540 20020 22596 20636
rect 22092 19572 22148 19582
rect 21868 16772 21924 16782
rect 21756 16716 21868 16772
rect 20300 16706 20356 16716
rect 21868 16706 21924 16716
rect 22092 16770 22148 19516
rect 22092 16718 22094 16770
rect 22146 16718 22148 16770
rect 22092 16660 22148 16718
rect 19836 16156 20100 16166
rect 19892 16100 19940 16156
rect 19996 16100 20044 16156
rect 19836 16090 20100 16100
rect 19740 15764 19796 15774
rect 19740 15670 19796 15708
rect 19852 15652 19908 15662
rect 19628 14644 19684 14654
rect 19628 14550 19684 14588
rect 19852 14306 19908 15596
rect 22092 15652 22148 16604
rect 22540 16770 22596 19964
rect 22652 18450 22708 21982
rect 22764 21812 22820 21822
rect 23212 21812 23268 23884
rect 23436 23604 23492 23614
rect 23436 23510 23492 23548
rect 23436 22594 23492 22606
rect 23436 22542 23438 22594
rect 23490 22542 23492 22594
rect 23436 22034 23492 22542
rect 23436 21982 23438 22034
rect 23490 21982 23492 22034
rect 23436 21970 23492 21982
rect 22764 21810 23268 21812
rect 22764 21758 22766 21810
rect 22818 21758 23214 21810
rect 23266 21758 23268 21810
rect 22764 21756 23268 21758
rect 22764 21700 22820 21756
rect 23212 21746 23268 21756
rect 22764 21634 22820 21644
rect 23212 20692 23268 20702
rect 23212 19682 23268 20636
rect 23660 20692 23716 20702
rect 23660 20598 23716 20636
rect 23212 19630 23214 19682
rect 23266 19630 23268 19682
rect 23212 19618 23268 19630
rect 22764 19572 22820 19582
rect 22764 19478 22820 19516
rect 22652 18398 22654 18450
rect 22706 18398 22708 18450
rect 22652 17890 22708 18398
rect 22652 17838 22654 17890
rect 22706 17838 22708 17890
rect 22652 17826 22708 17838
rect 23660 17554 23716 17566
rect 23660 17502 23662 17554
rect 23714 17502 23716 17554
rect 22540 16718 22542 16770
rect 22594 16718 22596 16770
rect 22540 16548 22596 16718
rect 22988 16772 23044 16782
rect 22988 16678 23044 16716
rect 23212 16772 23268 16782
rect 22540 16482 22596 16492
rect 23212 15874 23268 16716
rect 23660 16772 23716 17502
rect 23660 16706 23716 16716
rect 23436 16548 23492 16558
rect 23212 15822 23214 15874
rect 23266 15822 23268 15874
rect 23212 15810 23268 15822
rect 23324 16492 23436 16548
rect 22092 15586 22148 15596
rect 20188 15426 20244 15438
rect 20188 15374 20190 15426
rect 20242 15374 20244 15426
rect 20188 14868 20244 15374
rect 20188 14774 20244 14812
rect 20748 15092 20804 15102
rect 20076 14532 20132 14542
rect 19964 14530 20356 14532
rect 19964 14478 20078 14530
rect 20130 14478 20356 14530
rect 19964 14476 20356 14478
rect 19964 14420 20020 14476
rect 20076 14438 20132 14476
rect 19964 14354 20020 14364
rect 19852 14254 19854 14306
rect 19906 14254 19908 14306
rect 19852 14242 19908 14254
rect 20076 14308 20132 14318
rect 20076 14306 20244 14308
rect 20076 14254 20078 14306
rect 20130 14254 20244 14306
rect 20076 14252 20244 14254
rect 20076 14242 20132 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13972 20244 14252
rect 20076 13916 20244 13972
rect 20076 13746 20132 13916
rect 20076 13694 20078 13746
rect 20130 13694 20132 13746
rect 20076 13682 20132 13694
rect 19740 13636 19796 13646
rect 19516 13634 19796 13636
rect 19516 13582 19742 13634
rect 19794 13582 19796 13634
rect 19516 13580 19796 13582
rect 20300 13636 20356 14476
rect 20412 13636 20468 13646
rect 20300 13634 20468 13636
rect 20300 13582 20414 13634
rect 20466 13582 20468 13634
rect 20300 13580 20468 13582
rect 19292 12798 19294 12850
rect 19346 12798 19348 12850
rect 19292 12786 19348 12798
rect 17500 12626 17668 12628
rect 17500 12574 17502 12626
rect 17554 12574 17668 12626
rect 17500 12572 17668 12574
rect 17500 12562 17556 12572
rect 18956 12516 19012 12526
rect 19740 12516 19796 13580
rect 18956 12514 19796 12516
rect 18956 12462 18958 12514
rect 19010 12462 19796 12514
rect 18956 12460 19796 12462
rect 18620 11620 18676 11630
rect 4476 11116 4740 11126
rect 4532 11060 4580 11116
rect 4636 11060 4684 11116
rect 4476 11050 4740 11060
rect 18172 9828 18228 9838
rect 18172 9734 18228 9772
rect 18620 9602 18676 11564
rect 18956 10724 19012 12460
rect 19836 12124 20100 12134
rect 19892 12068 19940 12124
rect 19996 12068 20044 12124
rect 19836 12058 20100 12068
rect 20412 11732 20468 13580
rect 20524 11732 20580 11742
rect 20412 11730 20580 11732
rect 20412 11678 20526 11730
rect 20578 11678 20580 11730
rect 20412 11676 20580 11678
rect 19740 11620 19796 11630
rect 19740 11526 19796 11564
rect 19404 11508 19460 11518
rect 18956 10658 19012 10668
rect 19068 11452 19404 11508
rect 18620 9550 18622 9602
rect 18674 9550 18676 9602
rect 18620 9538 18676 9550
rect 19068 9828 19124 11452
rect 19404 11414 19460 11452
rect 20524 11508 20580 11676
rect 20300 10946 20356 10958
rect 20300 10894 20302 10946
rect 20354 10894 20356 10946
rect 20300 10722 20356 10894
rect 20300 10670 20302 10722
rect 20354 10670 20356 10722
rect 19836 10108 20100 10118
rect 19892 10052 19940 10108
rect 19996 10052 20044 10108
rect 19836 10042 20100 10052
rect 20300 10052 20356 10670
rect 20524 10500 20580 11452
rect 20748 10946 20804 15036
rect 21420 15092 21476 15102
rect 21420 14532 21476 15036
rect 21420 14438 21476 14476
rect 22204 14530 22260 14542
rect 22204 14478 22206 14530
rect 22258 14478 22260 14530
rect 21756 14420 21812 14430
rect 21868 14420 21924 14430
rect 22204 14420 22260 14478
rect 22876 14530 22932 14542
rect 22876 14478 22878 14530
rect 22930 14478 22932 14530
rect 21812 14418 22260 14420
rect 21812 14366 21870 14418
rect 21922 14366 22260 14418
rect 21812 14364 22260 14366
rect 22540 14420 22596 14430
rect 20972 13636 21028 13646
rect 20972 13542 21028 13580
rect 21756 13636 21812 14364
rect 21868 14354 21924 14364
rect 22540 14326 22596 14364
rect 21308 12516 21364 12526
rect 21756 12516 21812 13580
rect 22428 12740 22484 12750
rect 22876 12740 22932 14478
rect 23212 14530 23268 14542
rect 23212 14478 23214 14530
rect 23266 14478 23268 14530
rect 23212 13412 23268 14478
rect 23324 14532 23380 16492
rect 23436 16454 23492 16492
rect 23660 15876 23716 15886
rect 23660 15782 23716 15820
rect 23772 14644 23828 24444
rect 24108 24434 24164 24444
rect 24556 23940 24612 25116
rect 24892 24836 24948 26462
rect 24780 24780 24948 24836
rect 25116 24836 25172 28590
rect 25340 28420 25396 28430
rect 25340 28326 25396 28364
rect 25340 28084 25396 28094
rect 25340 27990 25396 28028
rect 25452 27634 25508 28700
rect 25788 28642 25844 30268
rect 25900 29988 25956 29998
rect 26124 29988 26180 33964
rect 26236 33954 26292 33964
rect 26348 34020 26404 35756
rect 26572 35700 26628 35710
rect 26572 35698 26740 35700
rect 26572 35646 26574 35698
rect 26626 35646 26740 35698
rect 26572 35644 26740 35646
rect 26572 35634 26628 35644
rect 26684 34804 26740 35644
rect 26908 35252 26964 41468
rect 27020 41458 27076 41468
rect 27132 40964 27188 41692
rect 27132 40962 27300 40964
rect 27132 40910 27134 40962
rect 27186 40910 27300 40962
rect 27132 40908 27300 40910
rect 27132 40898 27188 40908
rect 27244 37940 27300 40908
rect 27916 40404 27972 41918
rect 28028 41076 28084 42812
rect 28140 43652 28196 44718
rect 29148 44996 29204 45006
rect 28252 44660 28308 44670
rect 28252 44566 28308 44604
rect 28700 44660 28756 44670
rect 28700 44098 28756 44604
rect 28700 44046 28702 44098
rect 28754 44046 28756 44098
rect 28700 43988 28756 44046
rect 29036 43988 29092 43998
rect 28700 43932 29036 43988
rect 28700 43708 28756 43932
rect 29036 43894 29092 43932
rect 29148 43708 29204 44940
rect 32060 44882 32116 46172
rect 32284 46134 32340 46172
rect 32396 44996 32452 46844
rect 32508 46788 32564 47740
rect 32620 47730 32676 47740
rect 32620 47012 32676 47022
rect 32620 46898 32676 46956
rect 32620 46846 32622 46898
rect 32674 46846 32676 46898
rect 32620 46834 32676 46846
rect 33068 46900 33124 48748
rect 33068 46834 33124 46844
rect 33516 48802 33572 49086
rect 33516 48750 33518 48802
rect 33570 48750 33572 48802
rect 32508 46116 32564 46732
rect 33180 46676 33236 46686
rect 33180 46582 33236 46620
rect 32508 46050 32564 46060
rect 33516 46340 33572 48750
rect 36988 48916 37044 48926
rect 35532 48690 35588 48702
rect 35532 48638 35534 48690
rect 35586 48638 35588 48690
rect 35532 48130 35588 48638
rect 35532 48078 35534 48130
rect 35586 48078 35588 48130
rect 35196 47404 35460 47414
rect 35252 47348 35300 47404
rect 35356 47348 35404 47404
rect 35196 47338 35460 47348
rect 34188 47012 34244 47022
rect 34076 46900 34132 46910
rect 34076 46806 34132 46844
rect 33852 46674 33908 46686
rect 33852 46622 33854 46674
rect 33906 46622 33908 46674
rect 33852 46340 33908 46622
rect 33516 46284 33908 46340
rect 33068 46004 33124 46014
rect 33068 45910 33124 45948
rect 33404 45892 33460 45902
rect 33180 45890 33460 45892
rect 33180 45838 33406 45890
rect 33458 45838 33460 45890
rect 33180 45836 33460 45838
rect 32396 44930 32452 44940
rect 32620 45108 32676 45118
rect 32060 44830 32062 44882
rect 32114 44830 32116 44882
rect 30492 44770 30548 44782
rect 30492 44718 30494 44770
rect 30546 44718 30548 44770
rect 30492 44098 30548 44718
rect 30492 44046 30494 44098
rect 30546 44046 30548 44098
rect 30492 44034 30548 44046
rect 30828 44770 30884 44782
rect 30828 44718 30830 44770
rect 30882 44718 30884 44770
rect 28140 42756 28196 43596
rect 28140 42662 28196 42700
rect 28588 43652 28756 43708
rect 29036 43652 29204 43708
rect 30268 43988 30324 43998
rect 28588 42642 28644 43652
rect 29036 42980 29092 43652
rect 29036 42866 29092 42924
rect 29036 42814 29038 42866
rect 29090 42814 29092 42866
rect 29036 42802 29092 42814
rect 30268 42866 30324 43932
rect 30828 43708 30884 44718
rect 31164 44770 31220 44782
rect 31164 44718 31166 44770
rect 31218 44718 31220 44770
rect 31164 44212 31220 44718
rect 31500 44658 31556 44670
rect 31500 44606 31502 44658
rect 31554 44606 31556 44658
rect 31276 44212 31332 44222
rect 31164 44210 31332 44212
rect 31164 44158 31278 44210
rect 31330 44158 31332 44210
rect 31164 44156 31332 44158
rect 31276 44146 31332 44156
rect 31500 43708 31556 44606
rect 31724 43988 31780 43998
rect 31724 43874 31780 43932
rect 31724 43822 31726 43874
rect 31778 43822 31780 43874
rect 31724 43810 31780 43822
rect 30268 42814 30270 42866
rect 30322 42814 30324 42866
rect 30268 42802 30324 42814
rect 30380 43652 30884 43708
rect 30940 43652 31556 43708
rect 32060 43764 32116 44830
rect 32620 44882 32676 45052
rect 32620 44830 32622 44882
rect 32674 44830 32676 44882
rect 32620 44818 32676 44830
rect 32172 43988 32228 43998
rect 32172 43894 32228 43932
rect 33180 43708 33236 45836
rect 33404 45826 33460 45836
rect 32060 43698 32116 43708
rect 32396 43652 33236 43708
rect 33292 44658 33348 44670
rect 33292 44606 33294 44658
rect 33346 44606 33348 44658
rect 28588 42590 28590 42642
rect 28642 42590 28644 42642
rect 28588 41972 28644 42590
rect 29372 42754 29428 42766
rect 29372 42702 29374 42754
rect 29426 42702 29428 42754
rect 29372 42196 29428 42702
rect 29596 42756 29652 42766
rect 29652 42700 29764 42756
rect 29596 42662 29652 42700
rect 29372 42130 29428 42140
rect 29708 42084 29764 42700
rect 29708 42018 29764 42028
rect 28476 41916 28644 41972
rect 30268 41972 30324 41982
rect 28476 41860 28532 41916
rect 30268 41878 30324 41916
rect 28476 41794 28532 41804
rect 28140 41748 28196 41758
rect 28140 41654 28196 41692
rect 28812 41748 28868 41758
rect 28812 41654 28868 41692
rect 29820 41524 29876 41534
rect 28028 41010 28084 41020
rect 29708 41522 29876 41524
rect 29708 41470 29822 41522
rect 29874 41470 29876 41522
rect 29708 41468 29876 41470
rect 27916 40338 27972 40348
rect 27356 38724 27412 38734
rect 27356 38630 27412 38668
rect 27356 37940 27412 37950
rect 27244 37938 27412 37940
rect 27244 37886 27358 37938
rect 27410 37886 27412 37938
rect 27244 37884 27412 37886
rect 27356 37874 27412 37884
rect 28364 37492 28420 37502
rect 28028 37490 28420 37492
rect 28028 37438 28366 37490
rect 28418 37438 28420 37490
rect 28028 37436 28420 37438
rect 27356 36596 27412 36606
rect 27356 36502 27412 36540
rect 27916 36484 27972 36494
rect 27916 36390 27972 36428
rect 27804 35924 27860 35934
rect 27132 35922 27860 35924
rect 27132 35870 27806 35922
rect 27858 35870 27860 35922
rect 27132 35868 27860 35870
rect 27020 35812 27076 35822
rect 27020 35718 27076 35756
rect 26908 35186 26964 35196
rect 27132 35138 27188 35868
rect 27804 35858 27860 35868
rect 28028 35700 28084 37436
rect 28364 37426 28420 37436
rect 28364 36818 28420 36830
rect 28364 36766 28366 36818
rect 28418 36766 28420 36818
rect 28364 36596 28420 36766
rect 28364 36530 28420 36540
rect 29260 36596 29316 36606
rect 27804 35644 28084 35700
rect 27132 35086 27134 35138
rect 27186 35086 27188 35138
rect 27132 35074 27188 35086
rect 27580 35252 27636 35262
rect 26684 34710 26740 34748
rect 27356 34466 27412 34478
rect 27356 34414 27358 34466
rect 27410 34414 27412 34466
rect 27356 34132 27412 34414
rect 27020 34076 27412 34132
rect 26460 34020 26516 34030
rect 26348 34018 26516 34020
rect 26348 33966 26462 34018
rect 26514 33966 26516 34018
rect 26348 33964 26516 33966
rect 26348 31892 26404 33964
rect 26460 33954 26516 33964
rect 26684 34020 26740 34030
rect 26684 33794 26740 33964
rect 27020 34018 27076 34076
rect 27020 33966 27022 34018
rect 27074 33966 27076 34018
rect 27020 33954 27076 33966
rect 27356 33908 27412 33918
rect 27356 33814 27412 33852
rect 26684 33742 26686 33794
rect 26738 33742 26740 33794
rect 26684 33730 26740 33742
rect 27580 33794 27636 35196
rect 27804 34802 27860 35644
rect 29260 35588 29316 36540
rect 29484 35588 29540 35598
rect 28812 35532 29484 35588
rect 27804 34750 27806 34802
rect 27858 34750 27860 34802
rect 27804 34738 27860 34750
rect 28028 34804 28084 34814
rect 28028 34710 28084 34748
rect 28364 34690 28420 34702
rect 28364 34638 28366 34690
rect 28418 34638 28420 34690
rect 28364 34580 28420 34638
rect 28364 34514 28420 34524
rect 28812 34018 28868 35532
rect 28812 33966 28814 34018
rect 28866 33966 28868 34018
rect 28812 33954 28868 33966
rect 29260 34804 29316 34814
rect 27580 33742 27582 33794
rect 27634 33742 27636 33794
rect 27580 33730 27636 33742
rect 27916 33908 27972 33918
rect 27244 33684 27300 33694
rect 27244 33682 27412 33684
rect 27244 33630 27246 33682
rect 27298 33630 27412 33682
rect 27244 33628 27412 33630
rect 27244 33618 27300 33628
rect 26460 32116 26516 32126
rect 26516 32060 26628 32116
rect 26460 32050 26516 32060
rect 26348 31826 26404 31836
rect 25900 29874 25956 29932
rect 25900 29822 25902 29874
rect 25954 29822 25956 29874
rect 25900 29810 25956 29822
rect 26012 29932 26180 29988
rect 26460 30212 26516 30222
rect 26012 28868 26068 29932
rect 26124 29764 26180 29774
rect 26348 29764 26404 29774
rect 26124 29670 26180 29708
rect 26236 29708 26348 29764
rect 25788 28590 25790 28642
rect 25842 28590 25844 28642
rect 25788 28578 25844 28590
rect 25900 28812 26068 28868
rect 25564 28530 25620 28542
rect 25564 28478 25566 28530
rect 25618 28478 25620 28530
rect 25564 27972 25620 28478
rect 25900 28084 25956 28812
rect 26012 28644 26068 28654
rect 26236 28644 26292 29708
rect 26348 29670 26404 29708
rect 26348 29092 26404 29102
rect 26348 28998 26404 29036
rect 26460 28754 26516 30156
rect 26572 29874 26628 32060
rect 27020 30884 27076 30894
rect 26684 30658 26740 30670
rect 26684 30606 26686 30658
rect 26738 30606 26740 30658
rect 26684 30436 26740 30606
rect 27020 30658 27076 30828
rect 27356 30772 27412 33628
rect 27916 31332 27972 33852
rect 28588 33012 28644 33022
rect 28588 32898 28644 32956
rect 28588 32846 28590 32898
rect 28642 32846 28644 32898
rect 28588 32834 28644 32846
rect 28028 31556 28084 31566
rect 28028 31554 28644 31556
rect 28028 31502 28030 31554
rect 28082 31502 28644 31554
rect 28028 31500 28644 31502
rect 28028 31490 28084 31500
rect 27916 31276 28084 31332
rect 27916 31108 27972 31118
rect 27468 30772 27524 30782
rect 27356 30770 27524 30772
rect 27356 30718 27470 30770
rect 27522 30718 27524 30770
rect 27356 30716 27524 30718
rect 27468 30706 27524 30716
rect 27020 30606 27022 30658
rect 27074 30606 27076 30658
rect 27020 30594 27076 30606
rect 27244 30548 27300 30558
rect 27804 30548 27860 30558
rect 27244 30546 27412 30548
rect 27244 30494 27246 30546
rect 27298 30494 27412 30546
rect 27244 30492 27412 30494
rect 27244 30482 27300 30492
rect 26684 30370 26740 30380
rect 27020 30434 27076 30446
rect 27020 30382 27022 30434
rect 27074 30382 27076 30434
rect 27020 30100 27076 30382
rect 27020 30034 27076 30044
rect 27132 30100 27188 30110
rect 27132 30098 27300 30100
rect 27132 30046 27134 30098
rect 27186 30046 27300 30098
rect 27132 30044 27300 30046
rect 27132 30034 27188 30044
rect 26572 29822 26574 29874
rect 26626 29822 26628 29874
rect 26572 29810 26628 29822
rect 27020 29874 27076 29886
rect 27020 29822 27022 29874
rect 27074 29822 27076 29874
rect 26684 29652 26740 29662
rect 26684 29650 26852 29652
rect 26684 29598 26686 29650
rect 26738 29598 26852 29650
rect 26684 29596 26852 29598
rect 26684 29586 26740 29596
rect 26684 28756 26740 28766
rect 26460 28702 26462 28754
rect 26514 28702 26516 28754
rect 26460 28690 26516 28702
rect 26572 28754 26740 28756
rect 26572 28702 26686 28754
rect 26738 28702 26740 28754
rect 26572 28700 26740 28702
rect 26012 28642 26292 28644
rect 26012 28590 26014 28642
rect 26066 28590 26292 28642
rect 26012 28588 26292 28590
rect 26012 28578 26068 28588
rect 25564 27906 25620 27916
rect 25788 28028 25956 28084
rect 26012 28308 26068 28318
rect 25676 27748 25732 27758
rect 25676 27654 25732 27692
rect 25452 27582 25454 27634
rect 25506 27582 25508 27634
rect 25452 27570 25508 27582
rect 25788 27188 25844 28028
rect 26012 27972 26068 28252
rect 26572 27972 26628 28700
rect 26684 28690 26740 28700
rect 25900 27916 26068 27972
rect 26460 27916 26628 27972
rect 25900 27860 25956 27916
rect 26124 27860 26180 27870
rect 25900 27766 25956 27804
rect 26012 27858 26180 27860
rect 26012 27806 26126 27858
rect 26178 27806 26180 27858
rect 26012 27804 26180 27806
rect 25788 27122 25844 27132
rect 25676 26852 25732 26862
rect 25564 26180 25620 26190
rect 25564 25956 25620 26124
rect 25452 25954 25620 25956
rect 25452 25902 25566 25954
rect 25618 25902 25620 25954
rect 25452 25900 25620 25902
rect 25452 25284 25508 25900
rect 25564 25890 25620 25900
rect 25452 25218 25508 25228
rect 25564 25396 25620 25406
rect 25564 24836 25620 25340
rect 25116 24780 25284 24836
rect 24780 24388 24836 24780
rect 24892 24612 24948 24622
rect 24892 24518 24948 24556
rect 25004 24610 25060 24622
rect 25004 24558 25006 24610
rect 25058 24558 25060 24610
rect 25004 24500 25060 24558
rect 25004 24434 25060 24444
rect 24780 24332 24948 24388
rect 24556 23846 24612 23884
rect 24780 23828 24836 23838
rect 24108 23604 24164 23614
rect 24108 23510 24164 23548
rect 23884 23492 23940 23502
rect 23884 22708 23940 23436
rect 23884 21810 23940 22652
rect 24780 22706 24836 23772
rect 24892 23492 24948 24332
rect 25116 23716 25172 23726
rect 25116 23622 25172 23660
rect 24892 23426 24948 23436
rect 25228 22818 25284 24780
rect 25564 24722 25620 24780
rect 25564 24670 25566 24722
rect 25618 24670 25620 24722
rect 25564 24658 25620 24670
rect 25452 24500 25508 24510
rect 25228 22766 25230 22818
rect 25282 22766 25284 22818
rect 25228 22754 25284 22766
rect 25340 23826 25396 23838
rect 25340 23774 25342 23826
rect 25394 23774 25396 23826
rect 24780 22654 24782 22706
rect 24834 22654 24836 22706
rect 24780 22642 24836 22654
rect 25228 22596 25284 22606
rect 25228 22502 25284 22540
rect 23884 21758 23886 21810
rect 23938 21758 23940 21810
rect 23884 21746 23940 21758
rect 24108 22482 24164 22494
rect 24108 22430 24110 22482
rect 24162 22430 24164 22482
rect 24108 20188 24164 22430
rect 24892 22482 24948 22494
rect 24892 22430 24894 22482
rect 24946 22430 24948 22482
rect 24556 21700 24612 21710
rect 23996 20132 24164 20188
rect 24220 21588 24276 21598
rect 24220 20580 24276 21532
rect 24556 20914 24612 21644
rect 24668 21588 24724 21598
rect 24668 21586 24836 21588
rect 24668 21534 24670 21586
rect 24722 21534 24836 21586
rect 24668 21532 24836 21534
rect 24668 21522 24724 21532
rect 24556 20862 24558 20914
rect 24610 20862 24612 20914
rect 24556 20850 24612 20862
rect 24780 20914 24836 21532
rect 24780 20862 24782 20914
rect 24834 20862 24836 20914
rect 24780 20692 24836 20862
rect 24780 20626 24836 20636
rect 23996 19906 24052 20132
rect 23996 19854 23998 19906
rect 24050 19854 24052 19906
rect 23996 19842 24052 19854
rect 24220 18676 24276 20524
rect 23996 18674 24276 18676
rect 23996 18622 24222 18674
rect 24274 18622 24276 18674
rect 23996 18620 24276 18622
rect 23884 18002 23940 18014
rect 23884 17950 23886 18002
rect 23938 17950 23940 18002
rect 23884 16770 23940 17950
rect 23884 16718 23886 16770
rect 23938 16718 23940 16770
rect 23884 16706 23940 16718
rect 23996 16548 24052 18620
rect 24220 18610 24276 18620
rect 24332 19684 24388 19694
rect 24220 18002 24276 18014
rect 24220 17950 24222 18002
rect 24274 17950 24276 18002
rect 24220 17890 24276 17950
rect 24220 17838 24222 17890
rect 24274 17838 24276 17890
rect 24220 17826 24276 17838
rect 24220 16772 24276 16782
rect 23996 16482 24052 16492
rect 24108 16660 24164 16670
rect 24108 15874 24164 16604
rect 24220 16658 24276 16716
rect 24220 16606 24222 16658
rect 24274 16606 24276 16658
rect 24220 16594 24276 16606
rect 24108 15822 24110 15874
rect 24162 15822 24164 15874
rect 24108 15540 24164 15822
rect 24108 15474 24164 15484
rect 23884 14644 23940 14654
rect 23772 14642 23940 14644
rect 23772 14590 23886 14642
rect 23938 14590 23940 14642
rect 23772 14588 23940 14590
rect 23884 14578 23940 14588
rect 23324 13746 23380 14476
rect 23548 14530 23604 14542
rect 23548 14478 23550 14530
rect 23602 14478 23604 14530
rect 23548 14420 23604 14478
rect 23548 14354 23604 14364
rect 23324 13694 23326 13746
rect 23378 13694 23380 13746
rect 23324 13682 23380 13694
rect 23660 13412 23716 13422
rect 23212 13356 23660 13412
rect 22428 12738 22932 12740
rect 22428 12686 22430 12738
rect 22482 12686 22932 12738
rect 22428 12684 22932 12686
rect 22428 12674 22484 12684
rect 23660 12626 23716 13356
rect 23660 12574 23662 12626
rect 23714 12574 23716 12626
rect 23660 12562 23716 12574
rect 24332 12626 24388 19628
rect 24892 19348 24948 22430
rect 25340 22260 25396 23774
rect 25452 23716 25508 24444
rect 25564 23940 25620 23950
rect 25676 23940 25732 26796
rect 25900 25956 25956 25966
rect 26012 25956 26068 27804
rect 26124 27794 26180 27804
rect 26236 27860 26292 27870
rect 26236 27412 26292 27804
rect 26236 27346 26292 27356
rect 26348 27746 26404 27758
rect 26348 27694 26350 27746
rect 26402 27694 26404 27746
rect 26124 27188 26180 27198
rect 26348 27188 26404 27694
rect 26180 27132 26404 27188
rect 26124 27122 26180 27132
rect 26124 26964 26180 26974
rect 26124 26850 26180 26908
rect 26124 26798 26126 26850
rect 26178 26798 26180 26850
rect 26124 26786 26180 26798
rect 26236 25956 26292 27132
rect 26460 27076 26516 27916
rect 26460 27010 26516 27020
rect 26572 27746 26628 27758
rect 26572 27694 26574 27746
rect 26626 27694 26628 27746
rect 26348 26516 26404 26526
rect 26348 26422 26404 26460
rect 25900 25954 26068 25956
rect 25900 25902 25902 25954
rect 25954 25902 26068 25954
rect 25900 25900 26068 25902
rect 26124 25900 26292 25956
rect 25900 25890 25956 25900
rect 26124 24500 26180 25900
rect 26236 25730 26292 25742
rect 26460 25732 26516 25742
rect 26236 25678 26238 25730
rect 26290 25678 26292 25730
rect 26236 25508 26292 25678
rect 26236 25442 26292 25452
rect 26348 25730 26516 25732
rect 26348 25678 26462 25730
rect 26514 25678 26516 25730
rect 26348 25676 26516 25678
rect 26124 24434 26180 24444
rect 26236 24610 26292 24622
rect 26236 24558 26238 24610
rect 26290 24558 26292 24610
rect 26012 24386 26068 24398
rect 26012 24334 26014 24386
rect 26066 24334 26068 24386
rect 25900 23940 25956 23950
rect 25564 23938 25732 23940
rect 25564 23886 25566 23938
rect 25618 23886 25732 23938
rect 25564 23884 25732 23886
rect 25788 23884 25900 23940
rect 25564 23874 25620 23884
rect 25788 23828 25844 23884
rect 25900 23874 25956 23884
rect 25452 23650 25508 23660
rect 25676 23826 25844 23828
rect 25676 23774 25790 23826
rect 25842 23774 25844 23826
rect 25676 23772 25844 23774
rect 25564 22708 25620 22718
rect 25116 22204 25396 22260
rect 25452 22706 25620 22708
rect 25452 22654 25566 22706
rect 25618 22654 25620 22706
rect 25452 22652 25620 22654
rect 25116 21810 25172 22204
rect 25116 21758 25118 21810
rect 25170 21758 25172 21810
rect 25116 21746 25172 21758
rect 25452 21252 25508 22652
rect 25564 22642 25620 22652
rect 25676 22596 25732 23772
rect 25788 23762 25844 23772
rect 26012 23714 26068 24334
rect 26236 23828 26292 24558
rect 26348 24164 26404 25676
rect 26460 25666 26516 25676
rect 26572 24724 26628 27694
rect 26796 27748 26852 29596
rect 27020 28980 27076 29822
rect 27132 29876 27188 29886
rect 27132 29782 27188 29820
rect 27132 29204 27188 29214
rect 27244 29204 27300 30044
rect 27188 29148 27300 29204
rect 27132 29138 27188 29148
rect 27356 28980 27412 30492
rect 27468 30546 27860 30548
rect 27468 30494 27806 30546
rect 27858 30494 27860 30546
rect 27468 30492 27860 30494
rect 27468 30436 27524 30492
rect 27804 30482 27860 30492
rect 27468 29874 27524 30380
rect 27468 29822 27470 29874
rect 27522 29822 27524 29874
rect 27468 29810 27524 29822
rect 26908 28924 27860 28980
rect 26908 28754 26964 28924
rect 26908 28702 26910 28754
rect 26962 28702 26964 28754
rect 26908 28690 26964 28702
rect 27132 28754 27188 28766
rect 27132 28702 27134 28754
rect 27186 28702 27188 28754
rect 27132 28532 27188 28702
rect 27132 28466 27188 28476
rect 27244 28644 27300 28654
rect 27132 28196 27188 28206
rect 27020 28082 27076 28094
rect 27020 28030 27022 28082
rect 27074 28030 27076 28082
rect 26908 27972 26964 27982
rect 26908 27878 26964 27916
rect 27020 27860 27076 28030
rect 27020 27794 27076 27804
rect 27132 27858 27188 28140
rect 27132 27806 27134 27858
rect 27186 27806 27188 27858
rect 27132 27794 27188 27806
rect 27244 27860 27300 28588
rect 27356 28644 27412 28654
rect 27356 28642 27524 28644
rect 27356 28590 27358 28642
rect 27410 28590 27524 28642
rect 27356 28588 27524 28590
rect 27356 28578 27412 28588
rect 27356 27860 27412 27870
rect 27244 27858 27412 27860
rect 27244 27806 27358 27858
rect 27410 27806 27412 27858
rect 27244 27804 27412 27806
rect 27356 27794 27412 27804
rect 26796 27692 26908 27748
rect 26852 27636 26908 27692
rect 27020 27636 27076 27646
rect 26852 27580 26964 27636
rect 26796 27412 26852 27422
rect 26796 26964 26852 27356
rect 26796 26852 26852 26908
rect 26684 26796 26852 26852
rect 26684 26626 26740 26796
rect 26684 26574 26686 26626
rect 26738 26574 26740 26626
rect 26684 26562 26740 26574
rect 26796 26516 26852 26526
rect 26796 25956 26852 26460
rect 26908 26404 26964 27580
rect 27020 26626 27076 27580
rect 27468 26908 27524 28588
rect 27804 28530 27860 28924
rect 27804 28478 27806 28530
rect 27858 28478 27860 28530
rect 27580 28420 27636 28430
rect 27580 28326 27636 28364
rect 27804 27970 27860 28478
rect 27916 28308 27972 31052
rect 28028 29652 28084 31276
rect 28140 30996 28196 31006
rect 28140 30658 28196 30940
rect 28140 30606 28142 30658
rect 28194 30606 28196 30658
rect 28140 30436 28196 30606
rect 28140 30370 28196 30380
rect 28140 29876 28196 29886
rect 28252 29876 28308 31500
rect 28476 31108 28532 31118
rect 28476 31014 28532 31052
rect 28588 30772 28644 31500
rect 28588 30770 29204 30772
rect 28588 30718 28590 30770
rect 28642 30718 29204 30770
rect 28588 30716 29204 30718
rect 28588 30706 28644 30716
rect 29148 30658 29204 30716
rect 29148 30606 29150 30658
rect 29202 30606 29204 30658
rect 29148 30594 29204 30606
rect 29148 30436 29204 30446
rect 28140 29874 28308 29876
rect 28140 29822 28142 29874
rect 28194 29822 28308 29874
rect 28140 29820 28308 29822
rect 28476 29986 28532 29998
rect 28476 29934 28478 29986
rect 28530 29934 28532 29986
rect 28140 29810 28196 29820
rect 28364 29764 28420 29774
rect 28252 29708 28364 29764
rect 28028 29596 28196 29652
rect 28028 28868 28084 28878
rect 28028 28642 28084 28812
rect 28140 28756 28196 29596
rect 28140 28690 28196 28700
rect 28028 28590 28030 28642
rect 28082 28590 28084 28642
rect 28028 28578 28084 28590
rect 28252 28644 28308 29708
rect 28364 29698 28420 29708
rect 28476 29428 28532 29934
rect 28812 29986 28868 29998
rect 28812 29934 28814 29986
rect 28866 29934 28868 29986
rect 28812 29764 28868 29934
rect 29148 29874 29204 30380
rect 29148 29822 29150 29874
rect 29202 29822 29204 29874
rect 29148 29810 29204 29822
rect 28812 29698 28868 29708
rect 28476 29362 28532 29372
rect 28812 29428 28868 29438
rect 28252 28550 28308 28588
rect 27916 28242 27972 28252
rect 27804 27918 27806 27970
rect 27858 27918 27860 27970
rect 27804 27906 27860 27918
rect 28476 27972 28532 27982
rect 28140 27860 28196 27870
rect 28140 27766 28196 27804
rect 27356 26852 27524 26908
rect 28140 27524 28196 27534
rect 27356 26786 27412 26796
rect 28140 26850 28196 27468
rect 28476 26908 28532 27916
rect 28812 27860 28868 29372
rect 29148 28866 29204 28878
rect 29148 28814 29150 28866
rect 29202 28814 29204 28866
rect 29148 28756 29204 28814
rect 29260 28756 29316 34748
rect 29484 34802 29540 35532
rect 29708 35252 29764 41468
rect 29820 41458 29876 41468
rect 30380 40292 30436 43652
rect 30828 41972 30884 41982
rect 30940 41972 30996 43652
rect 30828 41970 30996 41972
rect 30828 41918 30830 41970
rect 30882 41918 30996 41970
rect 30828 41916 30996 41918
rect 30828 41906 30884 41916
rect 30380 40178 30436 40236
rect 30380 40126 30382 40178
rect 30434 40126 30436 40178
rect 30380 40114 30436 40126
rect 30940 41748 30996 41758
rect 31500 41748 31556 41758
rect 30996 41746 31556 41748
rect 30996 41694 31502 41746
rect 31554 41694 31556 41746
rect 30996 41692 31556 41694
rect 30716 39842 30772 39854
rect 30716 39790 30718 39842
rect 30770 39790 30772 39842
rect 30716 39732 30772 39790
rect 30716 39666 30772 39676
rect 29932 38724 29988 38734
rect 29820 35812 29876 35822
rect 29820 35718 29876 35756
rect 29708 35186 29764 35196
rect 29484 34750 29486 34802
rect 29538 34750 29540 34802
rect 29484 34738 29540 34750
rect 29372 34580 29428 34590
rect 29372 34486 29428 34524
rect 29484 33012 29540 33022
rect 29484 32674 29540 32956
rect 29820 32900 29876 32910
rect 29820 32786 29876 32844
rect 29820 32734 29822 32786
rect 29874 32734 29876 32786
rect 29820 32722 29876 32734
rect 29484 32622 29486 32674
rect 29538 32622 29540 32674
rect 29484 32610 29540 32622
rect 29932 32564 29988 38668
rect 30156 38724 30212 38734
rect 30604 38724 30660 38734
rect 30156 38722 30660 38724
rect 30156 38670 30158 38722
rect 30210 38670 30606 38722
rect 30658 38670 30660 38722
rect 30156 38668 30660 38670
rect 30156 38658 30212 38668
rect 30268 37716 30324 38668
rect 30604 38658 30660 38668
rect 30268 37650 30324 37660
rect 30604 35700 30660 35710
rect 30604 34916 30660 35644
rect 30940 35028 30996 41692
rect 31500 41682 31556 41692
rect 31836 40850 31892 40862
rect 31836 40798 31838 40850
rect 31890 40798 31892 40850
rect 31276 40628 31332 40638
rect 31836 40628 31892 40798
rect 31276 40626 31892 40628
rect 31276 40574 31278 40626
rect 31330 40574 31892 40626
rect 31276 40572 31892 40574
rect 31276 40562 31332 40572
rect 31836 40292 31892 40572
rect 31836 40226 31892 40236
rect 32060 39842 32116 39854
rect 32060 39790 32062 39842
rect 32114 39790 32116 39842
rect 31164 39732 31220 39742
rect 31724 39732 31780 39742
rect 32060 39732 32116 39790
rect 31220 39730 32116 39732
rect 31220 39678 31726 39730
rect 31778 39678 32116 39730
rect 31220 39676 32116 39678
rect 31164 39638 31220 39676
rect 31052 37716 31108 37726
rect 31052 36596 31108 37660
rect 31500 36596 31556 36606
rect 31052 36594 31556 36596
rect 31052 36542 31502 36594
rect 31554 36542 31556 36594
rect 31052 36540 31556 36542
rect 31388 35700 31444 36540
rect 31500 36530 31556 36540
rect 31388 35634 31444 35644
rect 31500 35588 31556 35598
rect 31612 35588 31668 39676
rect 31724 39666 31780 39676
rect 32396 39618 32452 43652
rect 33292 43092 33348 44606
rect 33404 43988 33460 43998
rect 33516 43988 33572 46284
rect 33740 45892 33796 45902
rect 34076 45892 34132 45902
rect 33740 45798 33796 45836
rect 33852 45890 34132 45892
rect 33852 45838 34078 45890
rect 34130 45838 34132 45890
rect 33852 45836 34132 45838
rect 33460 43932 33572 43988
rect 33628 44100 33684 44110
rect 33404 43922 33460 43932
rect 33628 43708 33684 44044
rect 33292 43026 33348 43036
rect 33404 43652 33684 43708
rect 32956 42868 33012 42878
rect 32956 42774 33012 42812
rect 33292 42868 33348 42878
rect 33404 42868 33460 43652
rect 33292 42866 33460 42868
rect 33292 42814 33294 42866
rect 33346 42814 33460 42866
rect 33292 42812 33460 42814
rect 33292 42802 33348 42812
rect 33404 42196 33460 42206
rect 33404 41748 33460 42140
rect 33852 41972 33908 45836
rect 34076 45826 34132 45836
rect 34076 44996 34132 45006
rect 34076 44902 34132 44940
rect 34188 44884 34244 46956
rect 34860 47012 34916 47022
rect 34860 46898 34916 46956
rect 34860 46846 34862 46898
rect 34914 46846 34916 46898
rect 34860 46834 34916 46846
rect 35196 46676 35252 46686
rect 34524 46228 34580 46238
rect 34524 46002 34580 46172
rect 34524 45950 34526 46002
rect 34578 45950 34580 46002
rect 34524 45938 34580 45950
rect 35196 46002 35252 46620
rect 35196 45950 35198 46002
rect 35250 45950 35252 46002
rect 35196 45938 35252 45950
rect 35196 45388 35460 45398
rect 35252 45332 35300 45388
rect 35356 45332 35404 45388
rect 35196 45322 35460 45332
rect 35308 45108 35364 45118
rect 35532 45108 35588 48078
rect 36988 47906 37044 48860
rect 39228 48916 39284 48926
rect 39564 48916 39620 48926
rect 39284 48914 39620 48916
rect 39284 48862 39566 48914
rect 39618 48862 39620 48914
rect 39284 48860 39620 48862
rect 39228 48822 39284 48860
rect 39564 48850 39620 48860
rect 38780 48804 38836 48814
rect 38780 48710 38836 48748
rect 40684 48804 40740 48814
rect 38332 48692 38388 48702
rect 38332 48598 38388 48636
rect 39004 48692 39060 48702
rect 36988 47854 36990 47906
rect 37042 47854 37044 47906
rect 36988 46900 37044 47854
rect 39004 47906 39060 48636
rect 39004 47854 39006 47906
rect 39058 47854 39060 47906
rect 39004 47842 39060 47854
rect 40348 47794 40404 47806
rect 40348 47742 40350 47794
rect 40402 47742 40404 47794
rect 36988 46834 37044 46844
rect 37548 46900 37604 46910
rect 37100 46674 37156 46686
rect 37100 46622 37102 46674
rect 37154 46622 37156 46674
rect 35644 46564 35700 46574
rect 35644 46562 35924 46564
rect 35644 46510 35646 46562
rect 35698 46510 35924 46562
rect 35644 46508 35924 46510
rect 35644 46498 35700 46508
rect 35868 46114 35924 46508
rect 35868 46062 35870 46114
rect 35922 46062 35924 46114
rect 35868 46050 35924 46062
rect 36988 45778 37044 45790
rect 36988 45726 36990 45778
rect 37042 45726 37044 45778
rect 36988 45332 37044 45726
rect 36988 45266 37044 45276
rect 35364 45052 35588 45108
rect 35308 45014 35364 45052
rect 34188 44100 34244 44828
rect 34524 44996 34580 45006
rect 34524 44884 34580 44940
rect 36092 44884 36148 44894
rect 34524 44882 34916 44884
rect 34524 44830 34526 44882
rect 34578 44830 34916 44882
rect 34524 44828 34916 44830
rect 34524 44818 34580 44828
rect 34188 44006 34244 44044
rect 33964 43092 34020 43102
rect 33964 42998 34020 43036
rect 34636 42868 34692 42878
rect 33852 41906 33908 41916
rect 34412 41972 34468 41982
rect 34412 41878 34468 41916
rect 33964 41860 34020 41870
rect 33964 41766 34020 41804
rect 33404 41746 33572 41748
rect 33404 41694 33406 41746
rect 33458 41694 33572 41746
rect 33404 41692 33572 41694
rect 33404 41682 33460 41692
rect 33180 40628 33236 40638
rect 33180 40626 33460 40628
rect 33180 40574 33182 40626
rect 33234 40574 33460 40626
rect 33180 40572 33460 40574
rect 33180 40562 33236 40572
rect 33404 39954 33460 40572
rect 33404 39902 33406 39954
rect 33458 39902 33460 39954
rect 33404 39890 33460 39902
rect 33516 39956 33572 41692
rect 34636 40962 34692 42812
rect 34636 40910 34638 40962
rect 34690 40910 34692 40962
rect 34636 40898 34692 40910
rect 34748 41524 34804 41534
rect 33516 39890 33572 39900
rect 33852 39954 33908 39966
rect 33852 39902 33854 39954
rect 33906 39902 33908 39954
rect 32396 39566 32398 39618
rect 32450 39566 32452 39618
rect 32172 38052 32228 38062
rect 31724 37938 31780 37950
rect 31724 37886 31726 37938
rect 31778 37886 31780 37938
rect 31724 36932 31780 37886
rect 32172 37938 32228 37996
rect 32172 37886 32174 37938
rect 32226 37886 32228 37938
rect 32172 37874 32228 37886
rect 31836 37826 31892 37838
rect 31836 37774 31838 37826
rect 31890 37774 31892 37826
rect 31836 37716 31892 37774
rect 32396 37716 32452 39566
rect 32956 39508 33012 39518
rect 31836 37660 32452 37716
rect 32060 36932 32116 36942
rect 31724 36930 32116 36932
rect 31724 36878 32062 36930
rect 32114 36878 32116 36930
rect 31724 36876 32116 36878
rect 32060 36866 32116 36876
rect 31836 35812 31892 35822
rect 31836 35718 31892 35756
rect 31500 35586 31668 35588
rect 31500 35534 31502 35586
rect 31554 35534 31668 35586
rect 31500 35532 31668 35534
rect 31500 35522 31556 35532
rect 30940 34972 31108 35028
rect 30268 34914 30996 34916
rect 30268 34862 30606 34914
rect 30658 34862 30996 34914
rect 30268 34860 30996 34862
rect 30268 34018 30324 34860
rect 30604 34850 30660 34860
rect 30268 33966 30270 34018
rect 30322 33966 30324 34018
rect 30268 33954 30324 33966
rect 30716 33796 30772 33806
rect 30716 33702 30772 33740
rect 30268 32788 30324 32798
rect 30324 32732 30436 32788
rect 30268 32722 30324 32732
rect 29820 32508 29988 32564
rect 30044 32674 30100 32686
rect 30044 32622 30046 32674
rect 30098 32622 30100 32674
rect 29372 31892 29428 31902
rect 29428 31836 29764 31892
rect 29372 31798 29428 31836
rect 29708 31778 29764 31836
rect 29708 31726 29710 31778
rect 29762 31726 29764 31778
rect 29708 31714 29764 31726
rect 29484 30660 29540 30670
rect 29484 30546 29540 30604
rect 29484 30494 29486 30546
rect 29538 30494 29540 30546
rect 29484 30482 29540 30494
rect 29820 30212 29876 32508
rect 30044 31948 30100 32622
rect 30380 32004 30436 32732
rect 30828 32786 30884 34860
rect 30940 34802 30996 34860
rect 30940 34750 30942 34802
rect 30994 34750 30996 34802
rect 30940 34738 30996 34750
rect 30828 32734 30830 32786
rect 30882 32734 30884 32786
rect 30828 32722 30884 32734
rect 30492 32676 30548 32686
rect 30492 32582 30548 32620
rect 30492 32004 30548 32014
rect 30380 32002 30548 32004
rect 30380 31950 30494 32002
rect 30546 31950 30548 32002
rect 30380 31948 30548 31950
rect 30044 31892 30324 31948
rect 30492 31938 30548 31948
rect 30156 30772 30212 30782
rect 30156 30712 30158 30716
rect 30210 30712 30212 30716
rect 30156 30678 30212 30712
rect 29932 30660 29988 30670
rect 29932 30566 29988 30604
rect 30044 30436 30100 30446
rect 30044 30342 30100 30380
rect 29820 30156 30212 30212
rect 29484 29092 29540 29102
rect 29484 28756 29540 29036
rect 29932 28980 29988 28990
rect 29932 28756 29988 28924
rect 29260 28700 29428 28756
rect 29148 28690 29204 28700
rect 28812 27766 28868 27804
rect 29260 28532 29316 28542
rect 29372 28532 29428 28700
rect 29484 28754 29988 28756
rect 29484 28702 29486 28754
rect 29538 28702 29934 28754
rect 29986 28702 29988 28754
rect 29484 28700 29988 28702
rect 29484 28690 29540 28700
rect 29932 28690 29988 28700
rect 29372 28476 29764 28532
rect 29260 27634 29316 28476
rect 29260 27582 29262 27634
rect 29314 27582 29316 27634
rect 29260 27524 29316 27582
rect 29260 27458 29316 27468
rect 28140 26798 28142 26850
rect 28194 26798 28196 26850
rect 28140 26786 28196 26798
rect 28364 26852 28532 26908
rect 28700 27076 28756 27086
rect 27020 26574 27022 26626
rect 27074 26574 27076 26626
rect 27020 26562 27076 26574
rect 27356 26628 27412 26666
rect 27356 26562 27412 26572
rect 27916 26626 27972 26638
rect 27916 26574 27918 26626
rect 27970 26574 27972 26626
rect 27468 26516 27524 26526
rect 27468 26422 27524 26460
rect 27356 26404 27412 26414
rect 26908 26402 27412 26404
rect 26908 26350 27358 26402
rect 27410 26350 27412 26402
rect 26908 26348 27412 26350
rect 27356 26338 27412 26348
rect 26348 24098 26404 24108
rect 26460 24668 26628 24724
rect 26684 25900 26852 25956
rect 27020 26180 27076 26190
rect 26460 23940 26516 24668
rect 26572 24500 26628 24510
rect 26572 24406 26628 24444
rect 26572 23940 26628 23950
rect 26460 23938 26628 23940
rect 26460 23886 26574 23938
rect 26626 23886 26628 23938
rect 26460 23884 26628 23886
rect 26572 23874 26628 23884
rect 26684 23940 26740 25900
rect 27020 25730 27076 26124
rect 27020 25678 27022 25730
rect 27074 25678 27076 25730
rect 27020 25666 27076 25678
rect 27804 25732 27860 25742
rect 27468 25620 27524 25630
rect 26908 25508 26964 25518
rect 26908 25414 26964 25452
rect 27020 24836 27076 24846
rect 27020 24742 27076 24780
rect 26684 23846 26740 23884
rect 27244 24612 27300 24622
rect 26348 23828 26404 23838
rect 26236 23772 26348 23828
rect 26348 23734 26404 23772
rect 26012 23662 26014 23714
rect 26066 23662 26068 23714
rect 26012 23650 26068 23662
rect 26124 23714 26180 23726
rect 26124 23662 26126 23714
rect 26178 23662 26180 23714
rect 25788 23604 25844 23614
rect 25788 22706 25844 23548
rect 25788 22654 25790 22706
rect 25842 22654 25844 22706
rect 25788 22642 25844 22654
rect 25676 22530 25732 22540
rect 26012 22594 26068 22606
rect 26012 22542 26014 22594
rect 26066 22542 26068 22594
rect 26012 22036 26068 22542
rect 26124 22372 26180 23662
rect 26908 23714 26964 23726
rect 26908 23662 26910 23714
rect 26962 23662 26964 23714
rect 26124 22306 26180 22316
rect 26348 23604 26404 23614
rect 26012 21980 26180 22036
rect 26012 21812 26068 21822
rect 25676 21810 26068 21812
rect 25676 21758 26014 21810
rect 26066 21758 26068 21810
rect 25676 21756 26068 21758
rect 25564 21700 25620 21710
rect 25564 21606 25620 21644
rect 25340 21196 25508 21252
rect 25004 20914 25060 20926
rect 25004 20862 25006 20914
rect 25058 20862 25060 20914
rect 25004 20804 25060 20862
rect 25340 20804 25396 21196
rect 25676 21140 25732 21756
rect 26012 21746 26068 21756
rect 26124 21588 26180 21980
rect 26124 21522 26180 21532
rect 26236 21586 26292 21598
rect 26236 21534 26238 21586
rect 26290 21534 26292 21586
rect 26236 21476 26292 21534
rect 26236 21410 26292 21420
rect 25452 21084 25732 21140
rect 25452 21026 25508 21084
rect 25452 20974 25454 21026
rect 25506 20974 25508 21026
rect 25452 20962 25508 20974
rect 25004 20802 25284 20804
rect 25004 20750 25006 20802
rect 25058 20750 25284 20802
rect 25004 20748 25284 20750
rect 25340 20748 25844 20804
rect 25004 20738 25060 20748
rect 25228 20580 25284 20748
rect 25340 20580 25396 20590
rect 25228 20578 25396 20580
rect 25228 20526 25342 20578
rect 25394 20526 25396 20578
rect 25228 20524 25396 20526
rect 25340 20132 25396 20524
rect 24892 19282 24948 19292
rect 25004 20076 25340 20132
rect 25004 18676 25060 20076
rect 25340 20066 25396 20076
rect 25564 20244 25620 20254
rect 25564 19906 25620 20188
rect 25788 20018 25844 20748
rect 26348 20802 26404 23548
rect 26796 21586 26852 21598
rect 26796 21534 26798 21586
rect 26850 21534 26852 21586
rect 26796 21476 26852 21534
rect 26796 21410 26852 21420
rect 26348 20750 26350 20802
rect 26402 20750 26404 20802
rect 25900 20466 25956 20478
rect 25900 20414 25902 20466
rect 25954 20414 25956 20466
rect 25900 20132 25956 20414
rect 26348 20188 26404 20750
rect 25900 20066 25956 20076
rect 26236 20132 26404 20188
rect 26908 20188 26964 23662
rect 27244 20188 27300 24556
rect 27468 24610 27524 25564
rect 27692 24724 27748 24734
rect 27804 24724 27860 25676
rect 27916 25620 27972 26574
rect 28252 26628 28308 26638
rect 28364 26628 28420 26852
rect 28476 26740 28532 26750
rect 28476 26646 28532 26684
rect 28252 26626 28420 26628
rect 28252 26574 28254 26626
rect 28306 26574 28420 26626
rect 28252 26572 28420 26574
rect 28252 26516 28308 26572
rect 28252 26450 28308 26460
rect 28364 25741 28420 25753
rect 28364 25689 28366 25741
rect 28418 25732 28420 25741
rect 28476 25732 28532 25742
rect 28418 25689 28476 25732
rect 28364 25676 28476 25689
rect 28476 25666 28532 25676
rect 28588 25730 28644 25742
rect 28588 25678 28590 25730
rect 28642 25678 28644 25730
rect 28028 25620 28084 25630
rect 27916 25618 28084 25620
rect 27916 25566 28030 25618
rect 28082 25566 28084 25618
rect 27916 25564 28084 25566
rect 27692 24722 27860 24724
rect 27692 24670 27694 24722
rect 27746 24670 27860 24722
rect 27692 24668 27860 24670
rect 27692 24658 27748 24668
rect 27468 24558 27470 24610
rect 27522 24558 27524 24610
rect 27468 24546 27524 24558
rect 27580 24386 27636 24398
rect 27580 24334 27582 24386
rect 27634 24334 27636 24386
rect 27580 23828 27636 24334
rect 27580 23762 27636 23772
rect 27804 23604 27860 23614
rect 27804 23510 27860 23548
rect 27692 23490 27748 23502
rect 27692 23438 27694 23490
rect 27746 23438 27748 23490
rect 27692 22594 27748 23438
rect 27692 22542 27694 22594
rect 27746 22542 27748 22594
rect 27692 22530 27748 22542
rect 27468 20356 27524 20366
rect 26460 20132 26516 20142
rect 26908 20132 27188 20188
rect 27244 20132 27412 20188
rect 25788 19966 25790 20018
rect 25842 19966 25844 20018
rect 25788 19954 25844 19966
rect 26236 20020 26292 20132
rect 26236 19954 26292 19964
rect 25564 19854 25566 19906
rect 25618 19854 25620 19906
rect 25564 19842 25620 19854
rect 26236 19684 26292 19694
rect 26236 19590 26292 19628
rect 25564 19572 25620 19582
rect 25564 18786 25620 19516
rect 25564 18734 25566 18786
rect 25618 18734 25620 18786
rect 25564 18722 25620 18734
rect 26460 18786 26516 20076
rect 26460 18734 26462 18786
rect 26514 18734 26516 18786
rect 26460 18722 26516 18734
rect 26796 19794 26852 19806
rect 26796 19742 26798 19794
rect 26850 19742 26852 19794
rect 24668 18674 25396 18676
rect 24668 18622 25006 18674
rect 25058 18622 25396 18674
rect 24668 18620 25396 18622
rect 24668 18002 24724 18620
rect 25004 18610 25060 18620
rect 24668 17950 24670 18002
rect 24722 17950 24724 18002
rect 24668 17890 24724 17950
rect 24668 17838 24670 17890
rect 24722 17838 24724 17890
rect 24668 17826 24724 17838
rect 25340 17778 25396 18620
rect 25340 17726 25342 17778
rect 25394 17726 25396 17778
rect 24444 16660 24500 16670
rect 24444 16566 24500 16604
rect 24780 16660 24836 16670
rect 24780 16566 24836 16604
rect 25340 16658 25396 17726
rect 26012 18564 26068 18574
rect 26012 16772 26068 18508
rect 26796 17892 26852 19742
rect 26908 19570 26964 19582
rect 26908 19518 26910 19570
rect 26962 19518 26964 19570
rect 26908 19348 26964 19518
rect 27020 19348 27076 19358
rect 26908 19346 27076 19348
rect 26908 19294 27022 19346
rect 27074 19294 27076 19346
rect 26908 19292 27076 19294
rect 27020 19282 27076 19292
rect 27132 19012 27188 20132
rect 26796 17826 26852 17836
rect 27020 18956 27188 19012
rect 27356 19346 27412 20132
rect 27468 20132 27524 20300
rect 28028 20188 28084 25564
rect 28588 25396 28644 25678
rect 28588 25330 28644 25340
rect 28700 25394 28756 27020
rect 28812 26516 28868 26526
rect 28812 25730 28868 26460
rect 28812 25678 28814 25730
rect 28866 25678 28868 25730
rect 28812 25666 28868 25678
rect 28924 26404 28980 26414
rect 28700 25342 28702 25394
rect 28754 25342 28756 25394
rect 28700 25330 28756 25342
rect 28140 25172 28196 25182
rect 28140 24834 28196 25116
rect 28924 25060 28980 26348
rect 28140 24782 28142 24834
rect 28194 24782 28196 24834
rect 28140 24612 28196 24782
rect 28812 25004 28980 25060
rect 29036 25730 29092 25742
rect 29036 25678 29038 25730
rect 29090 25678 29092 25730
rect 28140 24546 28196 24556
rect 28252 24724 28308 24734
rect 28252 23938 28308 24668
rect 28252 23886 28254 23938
rect 28306 23886 28308 23938
rect 28252 23716 28308 23886
rect 28252 23650 28308 23660
rect 28364 24500 28420 24510
rect 28364 22930 28420 24444
rect 28700 23828 28756 23838
rect 28364 22878 28366 22930
rect 28418 22878 28420 22930
rect 28364 22866 28420 22878
rect 28476 23772 28700 23828
rect 28812 23828 28868 25004
rect 29036 23940 29092 25678
rect 29484 25730 29540 28476
rect 29708 27970 29764 28476
rect 29708 27918 29710 27970
rect 29762 27918 29764 27970
rect 29708 27906 29764 27918
rect 30044 27858 30100 27870
rect 30044 27806 30046 27858
rect 30098 27806 30100 27858
rect 29708 27636 29764 27646
rect 29596 26514 29652 26526
rect 29596 26462 29598 26514
rect 29650 26462 29652 26514
rect 29596 26404 29652 26462
rect 29596 26338 29652 26348
rect 29708 25842 29764 27580
rect 30044 26740 30100 27806
rect 30156 27412 30212 30156
rect 30268 28756 30324 31892
rect 30492 31108 30548 31118
rect 30492 30772 30548 31052
rect 30492 29986 30548 30716
rect 30826 30772 30882 30782
rect 30940 30772 30996 30782
rect 30826 30770 30940 30772
rect 30826 30718 30828 30770
rect 30880 30718 30940 30770
rect 30826 30716 30940 30718
rect 30826 30706 30882 30716
rect 30940 30706 30996 30716
rect 30604 30660 30660 30670
rect 30604 30566 30660 30604
rect 30492 29934 30494 29986
rect 30546 29934 30548 29986
rect 30492 29922 30548 29934
rect 30716 30434 30772 30446
rect 30716 30382 30718 30434
rect 30770 30382 30772 30434
rect 30716 29988 30772 30382
rect 30716 29922 30772 29932
rect 30716 29092 30772 29102
rect 30268 28700 30660 28756
rect 30156 27346 30212 27356
rect 30380 28530 30436 28542
rect 30380 28478 30382 28530
rect 30434 28478 30436 28530
rect 30380 27858 30436 28478
rect 30604 27972 30660 28700
rect 30716 28642 30772 29036
rect 30716 28590 30718 28642
rect 30770 28590 30772 28642
rect 30716 28578 30772 28590
rect 31052 28084 31108 34972
rect 31276 33906 31332 33918
rect 31276 33854 31278 33906
rect 31330 33854 31332 33906
rect 31276 33796 31332 33854
rect 31276 33730 31332 33740
rect 31164 33682 31220 33694
rect 31164 33630 31166 33682
rect 31218 33630 31220 33682
rect 31164 32900 31220 33630
rect 31164 32834 31220 32844
rect 31276 32676 31332 32686
rect 31500 32676 31556 32686
rect 31332 32674 31556 32676
rect 31332 32622 31502 32674
rect 31554 32622 31556 32674
rect 31332 32620 31556 32622
rect 31276 32610 31332 32620
rect 31500 32610 31556 32620
rect 31612 32340 31668 35532
rect 31724 34580 31780 34590
rect 31724 34578 32340 34580
rect 31724 34526 31726 34578
rect 31778 34526 32340 34578
rect 31724 34524 32340 34526
rect 31724 34514 31780 34524
rect 32284 34130 32340 34524
rect 32284 34078 32286 34130
rect 32338 34078 32340 34130
rect 32284 34066 32340 34078
rect 31836 33908 31892 33918
rect 31836 33814 31892 33852
rect 32396 33684 32452 37660
rect 32396 33618 32452 33628
rect 32508 39506 33012 39508
rect 32508 39454 32958 39506
rect 33010 39454 33012 39506
rect 32508 39452 33012 39454
rect 32508 33236 32564 39452
rect 32956 39442 33012 39452
rect 33516 38612 33572 38622
rect 33180 38052 33236 38062
rect 33180 37958 33236 37996
rect 33516 37826 33572 38556
rect 33852 38610 33908 39902
rect 34076 39732 34132 39742
rect 34076 39638 34132 39676
rect 34636 39058 34692 39070
rect 34636 39006 34638 39058
rect 34690 39006 34692 39058
rect 34636 38668 34692 39006
rect 33852 38558 33854 38610
rect 33906 38558 33908 38610
rect 33852 38546 33908 38558
rect 34412 38612 34468 38622
rect 34524 38612 34692 38668
rect 34468 38556 34580 38612
rect 34412 38546 34468 38556
rect 33516 37774 33518 37826
rect 33570 37774 33572 37826
rect 32620 37492 32676 37502
rect 32620 37490 33460 37492
rect 32620 37438 32622 37490
rect 32674 37438 33460 37490
rect 32620 37436 33460 37438
rect 32620 37426 32676 37436
rect 33180 35700 33236 35710
rect 33180 35606 33236 35644
rect 31388 32284 31668 32340
rect 32172 33180 32564 33236
rect 32732 35364 32788 35374
rect 31164 30884 31220 30894
rect 31164 30790 31220 30828
rect 31276 30660 31332 30670
rect 31276 30566 31332 30604
rect 31164 29092 31220 29102
rect 31164 28866 31220 29036
rect 31164 28814 31166 28866
rect 31218 28814 31220 28866
rect 31164 28802 31220 28814
rect 31164 28084 31220 28094
rect 31052 28082 31220 28084
rect 31052 28030 31166 28082
rect 31218 28030 31220 28082
rect 31052 28028 31220 28030
rect 30716 27972 30772 27982
rect 30604 27970 30772 27972
rect 30604 27918 30718 27970
rect 30770 27918 30772 27970
rect 30604 27916 30772 27918
rect 30380 27806 30382 27858
rect 30434 27806 30436 27858
rect 30044 26674 30100 26684
rect 29708 25790 29710 25842
rect 29762 25790 29764 25842
rect 29484 25678 29486 25730
rect 29538 25678 29540 25730
rect 29484 25666 29540 25678
rect 29596 25730 29652 25742
rect 29596 25678 29598 25730
rect 29650 25678 29652 25730
rect 29372 25396 29428 25406
rect 29428 25340 29540 25396
rect 29372 25330 29428 25340
rect 29148 24780 29428 24836
rect 29148 24722 29204 24780
rect 29148 24670 29150 24722
rect 29202 24670 29204 24722
rect 29148 24658 29204 24670
rect 29372 24612 29428 24780
rect 29484 24834 29540 25340
rect 29484 24782 29486 24834
rect 29538 24782 29540 24834
rect 29484 24770 29540 24782
rect 29596 24612 29652 25678
rect 29708 24724 29764 25790
rect 30044 26516 30100 26526
rect 30044 24836 30100 26460
rect 30268 26066 30324 26078
rect 30268 26014 30270 26066
rect 30322 26014 30324 26066
rect 30268 25954 30324 26014
rect 30268 25902 30270 25954
rect 30322 25902 30324 25954
rect 30268 24948 30324 25902
rect 30380 25620 30436 27806
rect 30492 26514 30548 26526
rect 30492 26462 30494 26514
rect 30546 26462 30548 26514
rect 30492 26292 30548 26462
rect 30492 26226 30548 26236
rect 30716 25956 30772 27916
rect 30828 26738 30884 26750
rect 30828 26686 30830 26738
rect 30882 26686 30884 26738
rect 30828 26066 30884 26686
rect 30828 26014 30830 26066
rect 30882 26014 30884 26066
rect 30828 26002 30884 26014
rect 30940 26514 30996 26526
rect 30940 26462 30942 26514
rect 30994 26462 30996 26514
rect 30940 26404 30996 26462
rect 30716 25890 30772 25900
rect 30716 25732 30772 25742
rect 30940 25732 30996 26348
rect 30716 25730 30996 25732
rect 30716 25678 30718 25730
rect 30770 25678 30996 25730
rect 30716 25676 30996 25678
rect 30716 25666 30772 25676
rect 30380 25554 30436 25564
rect 31052 25172 31108 28028
rect 31164 28018 31220 28028
rect 31388 27860 31444 32284
rect 32060 30884 32116 30894
rect 32060 30790 32116 30828
rect 31500 30770 31556 30782
rect 31500 30718 31502 30770
rect 31554 30718 31556 30770
rect 31500 30436 31556 30718
rect 31836 30436 31892 30446
rect 31500 30380 31836 30436
rect 31836 29986 31892 30380
rect 31836 29934 31838 29986
rect 31890 29934 31892 29986
rect 31836 29922 31892 29934
rect 31612 29540 31668 29550
rect 31612 28866 31668 29484
rect 31612 28814 31614 28866
rect 31666 28814 31668 28866
rect 31164 27804 31444 27860
rect 31500 27860 31556 27870
rect 31164 25956 31220 27804
rect 31500 27766 31556 27804
rect 31612 27188 31668 28814
rect 32060 28532 32116 28542
rect 32060 28438 32116 28476
rect 32060 27860 32116 27870
rect 32172 27860 32228 33180
rect 32508 31554 32564 31566
rect 32508 31502 32510 31554
rect 32562 31502 32564 31554
rect 32508 30772 32564 31502
rect 32508 30706 32564 30716
rect 32620 31220 32676 31230
rect 32620 30770 32676 31164
rect 32732 30884 32788 35308
rect 33180 33460 33236 33470
rect 32732 30818 32788 30828
rect 33068 33458 33236 33460
rect 33068 33406 33182 33458
rect 33234 33406 33236 33458
rect 33068 33404 33236 33406
rect 32620 30718 32622 30770
rect 32674 30718 32676 30770
rect 32060 27858 32228 27860
rect 32060 27806 32062 27858
rect 32114 27806 32228 27858
rect 32060 27804 32228 27806
rect 32396 30324 32452 30334
rect 32396 28642 32452 30268
rect 32396 28590 32398 28642
rect 32450 28590 32452 28642
rect 32396 27860 32452 28590
rect 32060 27794 32116 27804
rect 31836 27636 31892 27646
rect 31836 27542 31892 27580
rect 31500 27132 31668 27188
rect 31724 27522 31780 27534
rect 31724 27470 31726 27522
rect 31778 27470 31780 27522
rect 31500 26908 31556 27132
rect 31276 26852 31556 26908
rect 31612 26964 31668 26974
rect 31276 26626 31332 26852
rect 31276 26574 31278 26626
rect 31330 26574 31332 26626
rect 31276 26292 31332 26574
rect 31276 26226 31332 26236
rect 31388 26628 31444 26638
rect 31164 25900 31332 25956
rect 31164 25732 31220 25742
rect 31164 25638 31220 25676
rect 31052 25106 31108 25116
rect 30268 24882 30324 24892
rect 30044 24770 30100 24780
rect 29820 24724 29876 24734
rect 29708 24668 29820 24724
rect 29820 24630 29876 24668
rect 29372 24556 29652 24612
rect 29260 24500 29316 24510
rect 29260 24406 29316 24444
rect 29708 24500 29764 24510
rect 29708 24498 30100 24500
rect 29708 24446 29710 24498
rect 29762 24446 30100 24498
rect 29708 24444 30100 24446
rect 29708 24434 29764 24444
rect 29036 23884 29428 23940
rect 28924 23828 28980 23838
rect 28812 23826 28980 23828
rect 28812 23774 28926 23826
rect 28978 23774 28980 23826
rect 28812 23772 28980 23774
rect 28476 23490 28532 23772
rect 28700 23734 28756 23772
rect 28924 23604 28980 23772
rect 29036 23716 29092 23726
rect 29036 23622 29092 23660
rect 28924 23538 28980 23548
rect 28476 23438 28478 23490
rect 28530 23438 28532 23490
rect 28476 20804 28532 23438
rect 29148 21812 29204 21822
rect 29148 21810 29316 21812
rect 29148 21758 29150 21810
rect 29202 21758 29316 21810
rect 29148 21756 29316 21758
rect 29148 21746 29204 21756
rect 28924 21586 28980 21598
rect 28924 21534 28926 21586
rect 28978 21534 28980 21586
rect 28924 21476 28980 21534
rect 28924 21410 28980 21420
rect 28588 20804 28644 20814
rect 28476 20802 29204 20804
rect 28476 20750 28590 20802
rect 28642 20750 29204 20802
rect 28476 20748 29204 20750
rect 28476 20356 28532 20748
rect 28588 20738 28644 20748
rect 29148 20690 29204 20748
rect 29148 20638 29150 20690
rect 29202 20638 29204 20690
rect 29148 20626 29204 20638
rect 28028 20132 28308 20188
rect 27468 19906 27524 20076
rect 27468 19854 27470 19906
rect 27522 19854 27524 19906
rect 27468 19842 27524 19854
rect 27356 19294 27358 19346
rect 27410 19294 27412 19346
rect 26796 17668 26852 17678
rect 26460 17666 26852 17668
rect 26460 17614 26798 17666
rect 26850 17614 26852 17666
rect 26460 17612 26852 17614
rect 26460 17554 26516 17612
rect 26796 17602 26852 17612
rect 26460 17502 26462 17554
rect 26514 17502 26516 17554
rect 26460 17490 26516 17502
rect 25340 16606 25342 16658
rect 25394 16606 25396 16658
rect 24668 15764 24724 15774
rect 25228 15764 25284 15774
rect 25340 15764 25396 16606
rect 24668 15762 25396 15764
rect 24668 15710 24670 15762
rect 24722 15710 25230 15762
rect 25282 15710 25396 15762
rect 24668 15708 25396 15710
rect 24668 15698 24724 15708
rect 25228 15698 25284 15708
rect 25228 15540 25284 15550
rect 25004 14868 25060 14878
rect 25004 14642 25060 14812
rect 25004 14590 25006 14642
rect 25058 14590 25060 14642
rect 25004 14578 25060 14590
rect 24444 14532 24500 14542
rect 24444 14530 24612 14532
rect 24444 14478 24446 14530
rect 24498 14478 24612 14530
rect 24444 14476 24612 14478
rect 24444 14466 24500 14476
rect 24444 13860 24500 13870
rect 24444 13766 24500 13804
rect 24556 13524 24612 14476
rect 25228 13860 25284 15484
rect 25340 14756 25396 15708
rect 25340 14690 25396 14700
rect 25788 16716 26012 16772
rect 25676 14418 25732 14430
rect 25676 14366 25678 14418
rect 25730 14366 25732 14418
rect 25340 13860 25396 13870
rect 25228 13858 25396 13860
rect 25228 13806 25342 13858
rect 25394 13806 25396 13858
rect 25228 13804 25396 13806
rect 25340 13748 25396 13804
rect 25676 13860 25732 14366
rect 25676 13794 25732 13804
rect 25788 13858 25844 16716
rect 26012 16706 26068 16716
rect 26796 16660 26852 16670
rect 26684 14756 26740 14766
rect 26572 14700 26684 14756
rect 25788 13806 25790 13858
rect 25842 13806 25844 13858
rect 25788 13794 25844 13806
rect 25900 14532 25956 14542
rect 25340 13682 25396 13692
rect 24892 13524 24948 13534
rect 24556 13468 24892 13524
rect 24332 12574 24334 12626
rect 24386 12574 24388 12626
rect 24332 12562 24388 12574
rect 24892 12626 24948 13468
rect 24892 12574 24894 12626
rect 24946 12574 24948 12626
rect 24892 12562 24948 12574
rect 21308 12514 21812 12516
rect 21308 12462 21310 12514
rect 21362 12462 21812 12514
rect 21308 12460 21812 12462
rect 21308 12450 21364 12460
rect 21756 11508 21812 12460
rect 23324 12514 23380 12526
rect 23324 12462 23326 12514
rect 23378 12462 23380 12514
rect 22764 11956 22820 11966
rect 22540 11954 22820 11956
rect 22540 11902 22766 11954
rect 22818 11902 22820 11954
rect 22540 11900 22820 11902
rect 22540 11618 22596 11900
rect 22764 11890 22820 11900
rect 23324 11954 23380 12462
rect 23324 11902 23326 11954
rect 23378 11902 23380 11954
rect 23324 11890 23380 11902
rect 23996 12514 24052 12526
rect 25452 12516 25508 12526
rect 23996 12462 23998 12514
rect 24050 12462 24052 12514
rect 22540 11566 22542 11618
rect 22594 11566 22596 11618
rect 22540 11554 22596 11566
rect 22988 11508 23044 11518
rect 23436 11508 23492 11518
rect 21812 11452 21924 11508
rect 21756 11442 21812 11452
rect 20748 10894 20750 10946
rect 20802 10894 20804 10946
rect 20748 10882 20804 10894
rect 21420 10724 21476 10734
rect 20748 10500 20804 10510
rect 20524 10444 20748 10500
rect 20748 10406 20804 10444
rect 20300 9986 20356 9996
rect 19068 9602 19124 9772
rect 19068 9550 19070 9602
rect 19122 9550 19124 9602
rect 19068 9538 19124 9550
rect 21308 9716 21364 9726
rect 21420 9716 21476 10668
rect 21868 10498 21924 11452
rect 23044 11506 23492 11508
rect 23044 11454 23438 11506
rect 23490 11454 23492 11506
rect 23044 11452 23492 11454
rect 22988 11414 23044 11452
rect 22876 10948 22932 10958
rect 21868 10446 21870 10498
rect 21922 10446 21924 10498
rect 21868 10434 21924 10446
rect 22316 10500 22372 10510
rect 21308 9714 21476 9716
rect 21308 9662 21310 9714
rect 21362 9662 21476 9714
rect 21308 9660 21476 9662
rect 21644 10052 21700 10062
rect 4476 9100 4740 9110
rect 4532 9044 4580 9100
rect 4636 9044 4684 9100
rect 4476 9034 4740 9044
rect 19836 8092 20100 8102
rect 19892 8036 19940 8092
rect 19996 8036 20044 8092
rect 19836 8026 20100 8036
rect 3836 7810 3892 7822
rect 3836 7758 3838 7810
rect 3890 7758 3892 7810
rect 3836 6804 3892 7758
rect 4284 7810 4340 7822
rect 4284 7758 4286 7810
rect 4338 7758 4340 7810
rect 4284 7476 4340 7758
rect 21308 7812 21364 9660
rect 21644 9602 21700 9996
rect 21644 9550 21646 9602
rect 21698 9550 21700 9602
rect 21644 8818 21700 9550
rect 21644 8766 21646 8818
rect 21698 8766 21700 8818
rect 21644 8706 21700 8766
rect 21644 8654 21646 8706
rect 21698 8654 21700 8706
rect 21644 8642 21700 8654
rect 22092 8708 22148 8718
rect 22092 8614 22148 8652
rect 22316 8428 22372 10444
rect 22876 9826 22932 10892
rect 22876 9774 22878 9826
rect 22930 9774 22932 9826
rect 22876 9762 22932 9774
rect 23436 9828 23492 11452
rect 23996 10948 24052 12462
rect 25116 12514 25508 12516
rect 25116 12462 25454 12514
rect 25506 12462 25508 12514
rect 25116 12460 25508 12462
rect 23996 10882 24052 10892
rect 24444 11620 24500 11630
rect 24444 10500 24500 11564
rect 24220 10498 24500 10500
rect 24220 10446 24446 10498
rect 24498 10446 24500 10498
rect 24220 10444 24500 10446
rect 23436 9762 23492 9772
rect 23660 9938 23716 9950
rect 23660 9886 23662 9938
rect 23714 9886 23716 9938
rect 23660 9826 23716 9886
rect 23660 9774 23662 9826
rect 23714 9774 23716 9826
rect 23660 9762 23716 9774
rect 23772 9828 23828 9838
rect 22988 8818 23044 8830
rect 22988 8766 22990 8818
rect 23042 8766 23044 8818
rect 22540 8708 22596 8718
rect 22540 8614 22596 8652
rect 22988 8706 23044 8766
rect 22988 8654 22990 8706
rect 23042 8654 23044 8706
rect 22988 8596 23044 8654
rect 23772 8708 23828 9772
rect 24220 9826 24276 10444
rect 24444 10434 24500 10444
rect 24668 11506 24724 11518
rect 24668 11454 24670 11506
rect 24722 11454 24724 11506
rect 24668 9940 24724 11454
rect 25116 10834 25172 12460
rect 25452 12450 25508 12460
rect 25116 10782 25118 10834
rect 25170 10782 25172 10834
rect 25116 10770 25172 10782
rect 25228 11732 25284 11742
rect 24668 9938 24948 9940
rect 24668 9886 24670 9938
rect 24722 9886 24948 9938
rect 24668 9884 24948 9886
rect 24668 9874 24724 9884
rect 24220 9774 24222 9826
rect 24274 9774 24276 9826
rect 24220 9762 24276 9774
rect 22988 8530 23044 8540
rect 23660 8596 23716 8606
rect 23660 8502 23716 8540
rect 23772 8594 23828 8652
rect 23772 8542 23774 8594
rect 23826 8542 23828 8594
rect 23772 8530 23828 8542
rect 23996 9716 24052 9726
rect 22876 8484 22932 8494
rect 22316 8372 22932 8428
rect 23996 8484 24052 9660
rect 24668 9716 24724 9726
rect 24668 9622 24724 9660
rect 23996 8418 24052 8428
rect 24892 8594 24948 9884
rect 25228 9716 25284 11676
rect 25900 11732 25956 14476
rect 26572 13860 26628 14700
rect 26684 14690 26740 14700
rect 26684 14532 26740 14542
rect 26796 14532 26852 16604
rect 27020 15988 27076 18956
rect 27132 18788 27188 18798
rect 27132 17780 27188 18732
rect 27356 18786 27412 19294
rect 27356 18734 27358 18786
rect 27410 18734 27412 18786
rect 27356 18722 27412 18734
rect 27804 17892 27860 17902
rect 27804 17798 27860 17836
rect 27132 17778 27300 17780
rect 27132 17726 27134 17778
rect 27186 17726 27300 17778
rect 27132 17724 27300 17726
rect 27132 17714 27188 17724
rect 27020 15922 27076 15932
rect 27132 14756 27188 14766
rect 27132 14662 27188 14700
rect 26740 14476 26852 14532
rect 26684 14438 26740 14476
rect 26684 13860 26740 13870
rect 26572 13858 26740 13860
rect 26572 13806 26686 13858
rect 26738 13806 26740 13858
rect 26572 13804 26740 13806
rect 26684 13794 26740 13804
rect 26236 13524 26292 13534
rect 26236 13430 26292 13468
rect 27020 13524 27076 13534
rect 27020 12740 27076 13468
rect 27244 13412 27300 17724
rect 27468 17668 27524 17678
rect 27468 17666 27748 17668
rect 27468 17614 27470 17666
rect 27522 17614 27748 17666
rect 27468 17612 27748 17614
rect 27468 17602 27524 17612
rect 27692 16324 27748 17612
rect 27804 16548 27860 16558
rect 27804 16454 27860 16492
rect 27692 16268 28084 16324
rect 28028 15986 28084 16268
rect 28028 15934 28030 15986
rect 28082 15934 28084 15986
rect 28028 15922 28084 15934
rect 28252 15764 28308 20132
rect 28364 19684 28420 19694
rect 28476 19684 28532 20300
rect 29260 20188 29316 21756
rect 29372 21476 29428 23884
rect 30044 21810 30100 24444
rect 30940 23828 30996 23838
rect 30940 23734 30996 23772
rect 30044 21758 30046 21810
rect 30098 21758 30100 21810
rect 30044 21746 30100 21758
rect 31276 22484 31332 25900
rect 31388 25842 31444 26572
rect 31612 26626 31668 26908
rect 31724 26908 31780 27470
rect 32396 27076 32452 27804
rect 31724 26852 31892 26908
rect 31612 26574 31614 26626
rect 31666 26574 31668 26626
rect 31612 26516 31668 26574
rect 31612 26450 31668 26460
rect 31388 25790 31390 25842
rect 31442 25790 31444 25842
rect 31388 25778 31444 25790
rect 31612 26292 31668 26302
rect 31388 25618 31444 25630
rect 31388 25566 31390 25618
rect 31442 25566 31444 25618
rect 31388 25060 31444 25566
rect 31388 24994 31444 25004
rect 31612 24834 31668 26236
rect 31724 25732 31780 25742
rect 31836 25732 31892 26852
rect 31724 25730 31892 25732
rect 31724 25678 31726 25730
rect 31778 25678 31892 25730
rect 31724 25676 31892 25678
rect 32172 25732 32228 25742
rect 31724 25666 31780 25676
rect 32172 25638 32228 25676
rect 32284 25732 32340 25742
rect 32396 25732 32452 27020
rect 32508 28532 32564 28542
rect 32620 28532 32676 30718
rect 33068 30770 33124 33404
rect 33180 33394 33236 33404
rect 33068 30718 33070 30770
rect 33122 30718 33124 30770
rect 33068 30706 33124 30718
rect 33404 30770 33460 37436
rect 33516 35810 33572 37774
rect 33516 35758 33518 35810
rect 33570 35758 33572 35810
rect 33516 35700 33572 35758
rect 33516 35634 33572 35644
rect 34076 36818 34132 36830
rect 34076 36766 34078 36818
rect 34130 36766 34132 36818
rect 34076 35700 34132 36766
rect 33628 35474 33684 35486
rect 33628 35422 33630 35474
rect 33682 35422 33684 35474
rect 33628 33906 33684 35422
rect 33740 34804 33796 34814
rect 33740 34710 33796 34748
rect 33964 34692 34020 34702
rect 34076 34692 34132 35644
rect 34748 35364 34804 41468
rect 34860 40180 34916 44828
rect 36092 44790 36148 44828
rect 36876 44884 36932 44894
rect 37100 44884 37156 46622
rect 37548 45778 37604 46844
rect 39116 46788 39172 46798
rect 38668 46786 39172 46788
rect 38668 46734 39118 46786
rect 39170 46734 39172 46786
rect 38668 46732 39172 46734
rect 37996 46674 38052 46686
rect 37996 46622 37998 46674
rect 38050 46622 38052 46674
rect 37548 45726 37550 45778
rect 37602 45726 37604 45778
rect 37548 44996 37604 45726
rect 37548 44902 37604 44940
rect 37884 45892 37940 45902
rect 37996 45892 38052 46622
rect 37884 45890 38052 45892
rect 37884 45838 37886 45890
rect 37938 45838 38052 45890
rect 37884 45836 38052 45838
rect 37884 45332 37940 45836
rect 36932 44882 37156 44884
rect 36932 44830 37102 44882
rect 37154 44830 37156 44882
rect 36932 44828 37156 44830
rect 36876 44818 36932 44828
rect 35196 43372 35460 43382
rect 35252 43316 35300 43372
rect 35356 43316 35404 43372
rect 35196 43306 35460 43316
rect 37100 43090 37156 44828
rect 37884 44882 37940 45276
rect 38668 45218 38724 46732
rect 39116 46722 39172 46732
rect 39452 46786 39508 46798
rect 39788 46788 39844 46798
rect 39452 46734 39454 46786
rect 39506 46734 39508 46786
rect 38668 45166 38670 45218
rect 38722 45166 38724 45218
rect 38668 45154 38724 45166
rect 39116 45890 39172 45902
rect 39116 45838 39118 45890
rect 39170 45838 39172 45890
rect 37996 44996 38052 45006
rect 38052 44940 38164 44996
rect 37996 44930 38052 44940
rect 37884 44830 37886 44882
rect 37938 44830 37940 44882
rect 37884 43876 37940 44830
rect 38108 44882 38164 44940
rect 38108 44830 38110 44882
rect 38162 44830 38164 44882
rect 38108 44210 38164 44830
rect 38108 44158 38110 44210
rect 38162 44158 38164 44210
rect 38108 44146 38164 44158
rect 38332 44882 38388 44894
rect 38332 44830 38334 44882
rect 38386 44830 38388 44882
rect 37996 43876 38052 43886
rect 37884 43820 37996 43876
rect 37324 43762 37380 43774
rect 37324 43710 37326 43762
rect 37378 43710 37380 43762
rect 37324 43708 37380 43710
rect 37772 43762 37828 43774
rect 37772 43710 37774 43762
rect 37826 43710 37828 43762
rect 37324 43652 37492 43708
rect 37100 43038 37102 43090
rect 37154 43038 37156 43090
rect 37100 43026 37156 43038
rect 36876 42980 36932 42990
rect 36428 42644 36484 42654
rect 36316 42642 36484 42644
rect 36316 42590 36430 42642
rect 36482 42590 36484 42642
rect 36316 42588 36484 42590
rect 35084 42082 35140 42094
rect 35084 42030 35086 42082
rect 35138 42030 35140 42082
rect 34972 40852 35028 40862
rect 35084 40852 35140 42030
rect 35756 41972 35812 41982
rect 35532 41860 35588 41870
rect 35196 41356 35460 41366
rect 35252 41300 35300 41356
rect 35356 41300 35404 41356
rect 35196 41290 35460 41300
rect 35532 40964 35588 41804
rect 35308 40962 35588 40964
rect 35308 40910 35534 40962
rect 35586 40910 35588 40962
rect 35308 40908 35588 40910
rect 35084 40796 35252 40852
rect 34972 40628 35028 40796
rect 35084 40628 35140 40638
rect 34972 40626 35140 40628
rect 34972 40574 35086 40626
rect 35138 40574 35140 40626
rect 34972 40572 35140 40574
rect 35084 40562 35140 40572
rect 35196 40292 35252 40796
rect 35196 40226 35252 40236
rect 34860 38946 34916 40124
rect 35084 40068 35140 40078
rect 35308 40068 35364 40908
rect 35532 40898 35588 40908
rect 35140 40012 35364 40068
rect 35084 39058 35140 40012
rect 35756 39844 35812 41916
rect 36316 41972 36372 42588
rect 36428 42578 36484 42588
rect 36316 41858 36372 41916
rect 36876 41970 36932 42924
rect 37100 42642 37156 42654
rect 37100 42590 37102 42642
rect 37154 42590 37156 42642
rect 37100 42530 37156 42590
rect 37100 42478 37102 42530
rect 37154 42478 37156 42530
rect 37100 42466 37156 42478
rect 36876 41918 36878 41970
rect 36930 41918 36932 41970
rect 36876 41906 36932 41918
rect 36316 41806 36318 41858
rect 36370 41806 36372 41858
rect 36316 41794 36372 41806
rect 36428 41860 36484 41870
rect 36428 41766 36484 41804
rect 37212 41634 37268 41646
rect 37212 41582 37214 41634
rect 37266 41582 37268 41634
rect 36428 40852 36484 40862
rect 36428 40758 36484 40796
rect 35980 40740 36036 40750
rect 35980 40180 36036 40684
rect 37100 40516 37156 40526
rect 35980 40114 36036 40124
rect 36988 40292 37044 40302
rect 36540 39956 36596 39966
rect 36540 39862 36596 39900
rect 35532 39842 35812 39844
rect 35532 39790 35758 39842
rect 35810 39790 35812 39842
rect 35532 39788 35812 39790
rect 35196 39340 35460 39350
rect 35252 39284 35300 39340
rect 35356 39284 35404 39340
rect 35196 39274 35460 39284
rect 35532 39172 35588 39788
rect 35756 39778 35812 39788
rect 35084 39006 35086 39058
rect 35138 39006 35140 39058
rect 35084 38994 35140 39006
rect 35308 39116 35588 39172
rect 34860 38894 34862 38946
rect 34914 38894 34916 38946
rect 34860 38882 34916 38894
rect 35308 38946 35364 39116
rect 35308 38894 35310 38946
rect 35362 38894 35364 38946
rect 35308 38882 35364 38894
rect 35532 38612 35588 39116
rect 36988 38834 37044 40236
rect 36988 38782 36990 38834
rect 37042 38782 37044 38834
rect 36988 38770 37044 38782
rect 36428 38722 36484 38734
rect 36428 38670 36430 38722
rect 36482 38670 36484 38722
rect 36428 38668 36484 38670
rect 35532 38546 35588 38556
rect 36316 38612 36484 38668
rect 36316 37716 36372 38556
rect 35196 37324 35460 37334
rect 35252 37268 35300 37324
rect 35356 37268 35404 37324
rect 35196 37258 35460 37268
rect 36316 36932 36372 37660
rect 36652 37716 36708 37726
rect 37100 37716 37156 40460
rect 37212 38836 37268 41582
rect 37324 39956 37380 39966
rect 37436 39956 37492 43652
rect 37548 43090 37604 43102
rect 37548 43038 37550 43090
rect 37602 43038 37604 43090
rect 37548 42978 37604 43038
rect 37548 42926 37550 42978
rect 37602 42926 37604 42978
rect 37548 42914 37604 42926
rect 37772 42868 37828 43710
rect 37772 42802 37828 42812
rect 37996 42642 38052 43820
rect 38108 43764 38164 43802
rect 38108 43698 38164 43708
rect 38332 43708 38388 44830
rect 39004 44210 39060 44222
rect 39004 44158 39006 44210
rect 39058 44158 39060 44210
rect 39004 44098 39060 44158
rect 39004 44046 39006 44098
rect 39058 44046 39060 44098
rect 39004 44034 39060 44046
rect 38556 43874 38612 43886
rect 38556 43822 38558 43874
rect 38610 43822 38612 43874
rect 38556 43708 38612 43822
rect 38332 43652 38724 43708
rect 38332 43090 38388 43652
rect 38332 43038 38334 43090
rect 38386 43038 38388 43090
rect 38332 43026 38388 43038
rect 38668 43650 38724 43652
rect 38668 43598 38670 43650
rect 38722 43598 38724 43650
rect 37996 42590 37998 42642
rect 38050 42590 38052 42642
rect 37996 42530 38052 42590
rect 37996 42478 37998 42530
rect 38050 42478 38052 42530
rect 37772 41860 37828 41870
rect 37996 41860 38052 42478
rect 37828 41804 38052 41860
rect 37772 41766 37828 41804
rect 37884 40740 37940 40750
rect 37380 39900 37492 39956
rect 37548 39956 37604 39966
rect 37548 39954 37716 39956
rect 37548 39902 37550 39954
rect 37602 39902 37716 39954
rect 37548 39900 37716 39902
rect 37324 39890 37380 39900
rect 37548 39890 37604 39900
rect 37212 38770 37268 38780
rect 37324 39732 37380 39742
rect 37324 39060 37380 39676
rect 37324 38834 37380 39004
rect 37324 38782 37326 38834
rect 37378 38782 37380 38834
rect 37324 38770 37380 38782
rect 37660 38834 37716 39900
rect 37884 39844 37940 40684
rect 37996 40516 38052 41804
rect 38668 42866 38724 43598
rect 39116 43650 39172 45838
rect 39452 45556 39508 46734
rect 39564 46786 39844 46788
rect 39564 46734 39790 46786
rect 39842 46734 39844 46786
rect 39564 46732 39844 46734
rect 39564 46114 39620 46732
rect 39788 46722 39844 46732
rect 40124 46676 40180 46686
rect 40124 46674 40292 46676
rect 40124 46622 40126 46674
rect 40178 46622 40292 46674
rect 40124 46620 40292 46622
rect 40124 46610 40180 46620
rect 39564 46062 39566 46114
rect 39618 46062 39620 46114
rect 39564 46050 39620 46062
rect 40124 46004 40180 46014
rect 40124 45910 40180 45948
rect 39564 45556 39620 45566
rect 39452 45500 39564 45556
rect 39564 44882 39620 45500
rect 40236 45332 40292 46620
rect 40348 46004 40404 47742
rect 40684 47572 40740 48748
rect 41356 48802 41412 48814
rect 41356 48750 41358 48802
rect 41410 48750 41412 48802
rect 41244 48690 41300 48702
rect 41244 48638 41246 48690
rect 41298 48638 41300 48690
rect 41020 47794 41076 47806
rect 41020 47742 41022 47794
rect 41074 47742 41076 47794
rect 41020 47682 41076 47742
rect 41020 47630 41022 47682
rect 41074 47630 41076 47682
rect 40796 47572 40852 47582
rect 40684 47570 40852 47572
rect 40684 47518 40798 47570
rect 40850 47518 40852 47570
rect 40684 47516 40852 47518
rect 40796 47506 40852 47516
rect 41020 46900 41076 47630
rect 41020 46834 41076 46844
rect 41244 46898 41300 48638
rect 41356 48692 41412 48750
rect 42588 48804 42644 48814
rect 42588 48710 42644 48748
rect 43148 48802 43204 48814
rect 43148 48750 43150 48802
rect 43202 48750 43204 48802
rect 41412 48636 41524 48692
rect 41356 48626 41412 48636
rect 41468 48132 41524 48636
rect 43148 48132 43204 48750
rect 43596 48804 43652 48814
rect 43652 48748 43764 48804
rect 43596 48738 43652 48748
rect 41468 48130 41860 48132
rect 41468 48078 41470 48130
rect 41522 48078 41860 48130
rect 41468 48076 41860 48078
rect 43148 48076 43428 48132
rect 41468 48066 41524 48076
rect 41580 47682 41636 47694
rect 41580 47630 41582 47682
rect 41634 47630 41636 47682
rect 41244 46846 41246 46898
rect 41298 46846 41300 46898
rect 41244 46834 41300 46846
rect 41356 47570 41412 47582
rect 41356 47518 41358 47570
rect 41410 47518 41412 47570
rect 40348 45938 40404 45948
rect 40684 46788 40740 46798
rect 40236 45266 40292 45276
rect 39564 44830 39566 44882
rect 39618 44830 39620 44882
rect 39564 44818 39620 44830
rect 39116 43598 39118 43650
rect 39170 43598 39172 43650
rect 39116 43586 39172 43598
rect 39228 44770 39284 44782
rect 39900 44772 39956 44782
rect 39228 44718 39230 44770
rect 39282 44718 39284 44770
rect 39228 42980 39284 44718
rect 39788 44770 39956 44772
rect 39788 44718 39902 44770
rect 39954 44718 39956 44770
rect 39788 44716 39956 44718
rect 40684 44772 40740 46732
rect 41132 46004 41188 46014
rect 41132 45910 41188 45948
rect 41356 45892 41412 47518
rect 41244 45890 41412 45892
rect 41244 45838 41358 45890
rect 41410 45838 41412 45890
rect 41244 45836 41412 45838
rect 40796 44772 40852 44782
rect 40684 44770 40964 44772
rect 40684 44718 40798 44770
rect 40850 44718 40964 44770
rect 40684 44716 40964 44718
rect 39452 43876 39508 43886
rect 39452 43782 39508 43820
rect 39228 42914 39284 42924
rect 39564 43764 39620 43774
rect 38668 42814 38670 42866
rect 38722 42814 38724 42866
rect 38444 40852 38500 40862
rect 38668 40852 38724 42814
rect 39452 42868 39508 42878
rect 39564 42868 39620 43708
rect 39788 42978 39844 44716
rect 39900 44706 39956 44716
rect 40796 44706 40852 44716
rect 40236 44658 40292 44670
rect 40236 44606 40238 44658
rect 40290 44606 40292 44658
rect 39900 43762 39956 43774
rect 39900 43710 39902 43762
rect 39954 43710 39956 43762
rect 39900 43650 39956 43710
rect 39900 43598 39902 43650
rect 39954 43598 39956 43650
rect 39900 43586 39956 43598
rect 39788 42926 39790 42978
rect 39842 42926 39844 42978
rect 39788 42914 39844 42926
rect 40124 43540 40180 43550
rect 39676 42868 39732 42878
rect 39452 42866 39676 42868
rect 39452 42814 39454 42866
rect 39506 42814 39676 42866
rect 39452 42812 39676 42814
rect 39452 42802 39508 42812
rect 39676 42802 39732 42812
rect 39228 42756 39284 42766
rect 38892 41972 38948 41982
rect 38780 40852 38836 40862
rect 38500 40796 38780 40852
rect 38444 40758 38500 40796
rect 37996 40450 38052 40460
rect 38444 40068 38500 40078
rect 38444 39954 38500 40012
rect 38444 39902 38446 39954
rect 38498 39902 38500 39954
rect 37996 39844 38052 39854
rect 37884 39788 37996 39844
rect 37996 39750 38052 39788
rect 37660 38782 37662 38834
rect 37714 38782 37716 38834
rect 37660 38770 37716 38782
rect 37996 38610 38052 38622
rect 37996 38558 37998 38610
rect 38050 38558 38052 38610
rect 36652 37714 37156 37716
rect 36652 37662 36654 37714
rect 36706 37662 37102 37714
rect 37154 37662 37156 37714
rect 36652 37660 37156 37662
rect 36652 37650 36708 37660
rect 37100 37604 37156 37660
rect 37660 37716 37716 37726
rect 37660 37622 37716 37660
rect 37100 37538 37156 37548
rect 36428 36932 36484 36942
rect 37996 36932 38052 38558
rect 38220 37826 38276 37838
rect 38220 37774 38222 37826
rect 38274 37774 38276 37826
rect 38220 37716 38276 37774
rect 38276 37660 38388 37716
rect 38220 37650 38276 37660
rect 36316 36930 36484 36932
rect 36316 36878 36430 36930
rect 36482 36878 36484 36930
rect 36316 36876 36484 36878
rect 36428 36866 36484 36876
rect 36988 36876 38052 36932
rect 36652 36146 36708 36158
rect 36652 36094 36654 36146
rect 36706 36094 36708 36146
rect 36204 36036 36260 36046
rect 36204 35942 36260 35980
rect 36652 36034 36708 36094
rect 36652 35982 36654 36034
rect 36706 35982 36708 36034
rect 36652 35970 36708 35982
rect 34748 35298 34804 35308
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35308 35140 35364 35150
rect 35308 35046 35364 35084
rect 35644 35140 35700 35150
rect 35196 34804 35252 34814
rect 35196 34710 35252 34748
rect 33964 34690 34132 34692
rect 33964 34638 33966 34690
rect 34018 34638 34132 34690
rect 33964 34636 34132 34638
rect 33964 34626 34020 34636
rect 33628 33854 33630 33906
rect 33682 33854 33684 33906
rect 33628 33842 33684 33854
rect 33516 32786 33572 32798
rect 33516 32734 33518 32786
rect 33570 32734 33572 32786
rect 33516 31780 33572 32734
rect 34076 32786 34132 34636
rect 34860 34692 34916 34702
rect 34860 34598 34916 34636
rect 35532 34692 35588 34702
rect 34188 33908 34244 33918
rect 34188 33906 34468 33908
rect 34188 33854 34190 33906
rect 34242 33854 34468 33906
rect 34188 33852 34468 33854
rect 34188 33842 34244 33852
rect 34412 33796 34468 33852
rect 35532 33906 35588 34636
rect 35532 33854 35534 33906
rect 35586 33854 35588 33906
rect 35532 33842 35588 33854
rect 35084 33796 35140 33806
rect 34412 33740 34804 33796
rect 34300 33684 34356 33694
rect 34300 33590 34356 33628
rect 34636 33460 34692 33470
rect 34076 32734 34078 32786
rect 34130 32734 34132 32786
rect 34076 32676 34132 32734
rect 34076 32610 34132 32620
rect 34300 33458 34692 33460
rect 34300 33406 34638 33458
rect 34690 33406 34692 33458
rect 34300 33404 34692 33406
rect 33516 31714 33572 31724
rect 33628 31892 34132 31948
rect 33404 30718 33406 30770
rect 33458 30718 33460 30770
rect 33404 30706 33460 30718
rect 32844 30658 32900 30670
rect 32844 30606 32846 30658
rect 32898 30606 32900 30658
rect 32844 30548 32900 30606
rect 33516 30660 33572 30670
rect 32732 28532 32788 28542
rect 32620 28530 32788 28532
rect 32620 28478 32734 28530
rect 32786 28478 32788 28530
rect 32620 28476 32788 28478
rect 32508 27634 32564 28476
rect 32508 27582 32510 27634
rect 32562 27582 32564 27634
rect 32508 26964 32564 27582
rect 32732 27300 32788 28476
rect 32732 27234 32788 27244
rect 32508 26898 32564 26908
rect 32508 26516 32564 26526
rect 32508 25842 32564 26460
rect 32508 25790 32510 25842
rect 32562 25790 32564 25842
rect 32508 25778 32564 25790
rect 32284 25730 32452 25732
rect 32284 25678 32286 25730
rect 32338 25678 32452 25730
rect 32284 25676 32452 25678
rect 32284 25666 32340 25676
rect 31612 24782 31614 24834
rect 31666 24782 31668 24834
rect 31612 23828 31668 24782
rect 31612 23762 31668 23772
rect 31836 25508 31892 25518
rect 29372 21410 29428 21420
rect 29596 21698 29652 21710
rect 29596 21646 29598 21698
rect 29650 21646 29652 21698
rect 29596 21028 29652 21646
rect 30380 21588 30436 21598
rect 30380 21494 30436 21532
rect 29708 21028 29764 21038
rect 29596 21026 29764 21028
rect 29596 20974 29710 21026
rect 29762 20974 29764 21026
rect 29596 20972 29764 20974
rect 29708 20962 29764 20972
rect 30156 20356 30212 20366
rect 29708 20244 29764 20254
rect 29260 20132 29540 20188
rect 28364 19682 28532 19684
rect 28364 19630 28366 19682
rect 28418 19630 28532 19682
rect 28364 19628 28532 19630
rect 28364 19618 28420 19628
rect 29484 19570 29540 20132
rect 29484 19518 29486 19570
rect 29538 19518 29540 19570
rect 29484 19506 29540 19518
rect 28588 18564 28644 18574
rect 28588 18470 28644 18508
rect 28364 17892 28420 17902
rect 28364 17778 28420 17836
rect 28364 17726 28366 17778
rect 28418 17726 28420 17778
rect 28364 17714 28420 17726
rect 28476 17780 28532 17790
rect 28476 16770 28532 17724
rect 29596 17780 29652 17790
rect 29596 17686 29652 17724
rect 28476 16718 28478 16770
rect 28530 16718 28532 16770
rect 28476 16706 28532 16718
rect 28924 17666 28980 17678
rect 28924 17614 28926 17666
rect 28978 17614 28980 17666
rect 28252 15698 28308 15708
rect 28924 16324 28980 17614
rect 28924 15538 28980 16268
rect 29260 16658 29316 16670
rect 29260 16606 29262 16658
rect 29314 16606 29316 16658
rect 29260 16548 29316 16606
rect 28924 15486 28926 15538
rect 28978 15486 28980 15538
rect 28364 15092 28420 15102
rect 28252 15036 28364 15092
rect 27580 14756 27636 14766
rect 27580 14642 27636 14700
rect 27580 14590 27582 14642
rect 27634 14590 27636 14642
rect 27580 14578 27636 14590
rect 28252 14532 28308 15036
rect 28364 15026 28420 15036
rect 28252 14438 28308 14476
rect 28700 14420 28756 14430
rect 28924 14420 28980 15486
rect 28700 14418 28980 14420
rect 28700 14366 28702 14418
rect 28754 14366 28980 14418
rect 28700 14364 28980 14366
rect 29148 15876 29204 15886
rect 28700 14354 28756 14364
rect 29148 13858 29204 15820
rect 29260 14866 29316 16492
rect 29708 15876 29764 20188
rect 30156 20188 30212 20300
rect 31276 20188 31332 22428
rect 30156 20132 30324 20188
rect 30268 20066 30324 20076
rect 30940 20132 31332 20188
rect 31388 21588 31444 21598
rect 30156 18788 30212 18798
rect 30940 18788 30996 20132
rect 31388 20018 31444 21532
rect 31724 20132 31780 20142
rect 31388 19966 31390 20018
rect 31442 19966 31444 20018
rect 31388 19954 31444 19966
rect 31612 20076 31724 20132
rect 30156 18694 30212 18732
rect 30492 18786 30996 18788
rect 30492 18734 30942 18786
rect 30994 18734 30996 18786
rect 30492 18732 30996 18734
rect 30492 18674 30548 18732
rect 30940 18722 30996 18732
rect 31612 19010 31668 20076
rect 31724 20066 31780 20076
rect 31724 19684 31780 19694
rect 31724 19590 31780 19628
rect 31612 18958 31614 19010
rect 31666 18958 31668 19010
rect 31612 18788 31668 18958
rect 31724 18788 31780 18798
rect 31612 18786 31780 18788
rect 31612 18734 31726 18786
rect 31778 18734 31780 18786
rect 31612 18732 31780 18734
rect 30492 18622 30494 18674
rect 30546 18622 30548 18674
rect 30492 18610 30548 18622
rect 31052 18676 31108 18686
rect 30044 18564 30100 18574
rect 30044 16658 30100 18508
rect 30044 16606 30046 16658
rect 30098 16606 30100 16658
rect 30044 16594 30100 16606
rect 30604 18002 30660 18014
rect 30604 17950 30606 18002
rect 30658 17950 30660 18002
rect 30604 17890 30660 17950
rect 30604 17838 30606 17890
rect 30658 17838 30660 17890
rect 30380 16324 30436 16334
rect 30380 16230 30436 16268
rect 29708 15762 29764 15820
rect 29708 15710 29710 15762
rect 29762 15710 29764 15762
rect 29708 15698 29764 15710
rect 30492 15650 30548 15662
rect 30492 15598 30494 15650
rect 30546 15598 30548 15650
rect 29260 14814 29262 14866
rect 29314 14814 29316 14866
rect 29260 14754 29316 14814
rect 29260 14702 29262 14754
rect 29314 14702 29316 14754
rect 29260 14690 29316 14702
rect 29820 14866 29876 14878
rect 29820 14814 29822 14866
rect 29874 14814 29876 14866
rect 29148 13806 29150 13858
rect 29202 13806 29204 13858
rect 29148 13794 29204 13806
rect 29708 14420 29764 14430
rect 28588 13748 28644 13758
rect 28588 13654 28644 13692
rect 29708 13748 29764 14364
rect 29708 13682 29764 13692
rect 27244 13346 27300 13356
rect 27020 12646 27076 12684
rect 25900 11638 25956 11676
rect 26124 12402 26180 12414
rect 26124 12350 26126 12402
rect 26178 12350 26180 12402
rect 25452 11620 25508 11630
rect 25452 11526 25508 11564
rect 25788 10386 25844 10398
rect 25788 10334 25790 10386
rect 25842 10334 25844 10386
rect 25788 10052 25844 10334
rect 26012 10052 26068 10062
rect 25676 9996 26012 10052
rect 25676 9828 25732 9996
rect 25676 9734 25732 9772
rect 25228 9650 25284 9660
rect 26012 9602 26068 9996
rect 26012 9550 26014 9602
rect 26066 9550 26068 9602
rect 26012 9538 26068 9550
rect 26124 8932 26180 12350
rect 27132 11732 27188 11742
rect 26348 11620 26404 11630
rect 26796 11620 26852 11630
rect 26348 11618 26852 11620
rect 26348 11566 26350 11618
rect 26402 11566 26798 11618
rect 26850 11566 26852 11618
rect 26348 11564 26852 11566
rect 26348 11554 26404 11564
rect 26796 10052 26852 11564
rect 27132 11618 27188 11676
rect 29484 11730 29540 11742
rect 29484 11678 29486 11730
rect 29538 11678 29540 11730
rect 27132 11566 27134 11618
rect 27186 11566 27188 11618
rect 27132 11554 27188 11566
rect 28812 11620 28868 11630
rect 26796 9986 26852 9996
rect 26572 9716 26628 9726
rect 26572 9602 26628 9660
rect 26572 9550 26574 9602
rect 26626 9550 26628 9602
rect 26572 9538 26628 9550
rect 28140 9716 28196 9726
rect 26236 8932 26292 8942
rect 26124 8930 26292 8932
rect 26124 8878 26238 8930
rect 26290 8878 26292 8930
rect 26124 8876 26292 8878
rect 26236 8866 26292 8876
rect 28140 8708 28196 9660
rect 28140 8614 28196 8652
rect 28812 9602 28868 11564
rect 29484 11396 29540 11678
rect 29820 11620 29876 14814
rect 30156 14866 30212 14878
rect 30156 14814 30158 14866
rect 30210 14814 30212 14866
rect 30156 14754 30212 14814
rect 30156 14702 30158 14754
rect 30210 14702 30212 14754
rect 30156 14690 30212 14702
rect 30492 14420 30548 15598
rect 30604 15428 30660 17838
rect 31052 17892 31108 18620
rect 31500 18564 31556 18574
rect 31052 17890 31444 17892
rect 31052 17838 31054 17890
rect 31106 17838 31444 17890
rect 31052 17836 31444 17838
rect 31052 17826 31108 17836
rect 30828 16548 30884 16558
rect 31052 16548 31108 16558
rect 30828 16454 30884 16492
rect 30940 16546 31108 16548
rect 30940 16494 31054 16546
rect 31106 16494 31108 16546
rect 30940 16492 31108 16494
rect 31388 16548 31444 17836
rect 31500 17890 31556 18508
rect 31612 18002 31668 18732
rect 31724 18722 31780 18732
rect 31612 17950 31614 18002
rect 31666 17950 31668 18002
rect 31612 17938 31668 17950
rect 31500 17838 31502 17890
rect 31554 17838 31556 17890
rect 31500 16772 31556 17838
rect 31500 16706 31556 16716
rect 31500 16548 31556 16558
rect 31388 16546 31556 16548
rect 31388 16494 31502 16546
rect 31554 16494 31556 16546
rect 31388 16492 31556 16494
rect 30604 15362 30660 15372
rect 30940 15540 30996 16492
rect 31052 16482 31108 16492
rect 31276 15988 31332 15998
rect 31276 15894 31332 15932
rect 30492 14354 30548 14364
rect 30940 14420 30996 15484
rect 31276 15428 31332 15438
rect 31276 14532 31332 15372
rect 31500 15092 31556 16492
rect 31500 15026 31556 15036
rect 31724 15650 31780 15662
rect 31724 15598 31726 15650
rect 31778 15598 31780 15650
rect 30940 14326 30996 14364
rect 31164 14530 31332 14532
rect 31164 14478 31278 14530
rect 31330 14478 31332 14530
rect 31164 14476 31332 14478
rect 30940 13860 30996 13870
rect 31164 13860 31220 14476
rect 31276 14466 31332 14476
rect 30940 13858 31220 13860
rect 30940 13806 30942 13858
rect 30994 13806 31220 13858
rect 30940 13804 31220 13806
rect 30940 13794 30996 13804
rect 30380 13412 30436 13422
rect 30380 12626 30436 13356
rect 30380 12574 30382 12626
rect 30434 12574 30436 12626
rect 30380 12562 30436 12574
rect 30044 12516 30100 12526
rect 30044 12514 30212 12516
rect 30044 12462 30046 12514
rect 30098 12462 30212 12514
rect 30044 12460 30212 12462
rect 30044 12450 30100 12460
rect 29820 11526 29876 11564
rect 29484 11330 29540 11340
rect 28812 9550 28814 9602
rect 28866 9550 28868 9602
rect 24892 8542 24894 8594
rect 24946 8542 24948 8594
rect 21308 7746 21364 7756
rect 22316 7812 22372 7822
rect 22316 7718 22372 7756
rect 22764 7810 22820 8372
rect 22764 7758 22766 7810
rect 22818 7758 22820 7810
rect 22764 7746 22820 7758
rect 24892 7812 24948 8542
rect 28588 8596 28644 8606
rect 27692 8484 27748 8522
rect 28588 8502 28644 8540
rect 27692 8418 27748 8428
rect 28700 8484 28756 8494
rect 28812 8428 28868 9550
rect 29708 10052 29764 10062
rect 28700 8372 28868 8428
rect 29148 8708 29204 8718
rect 24892 7746 24948 7756
rect 28252 7812 28308 7822
rect 28252 7718 28308 7756
rect 28700 7810 28756 8372
rect 28700 7758 28702 7810
rect 28754 7758 28756 7810
rect 28700 7746 28756 7758
rect 29148 7700 29204 8652
rect 29596 8708 29652 8718
rect 29260 8596 29316 8606
rect 29260 8428 29316 8540
rect 29596 8594 29652 8652
rect 29596 8542 29598 8594
rect 29650 8542 29652 8594
rect 29596 8530 29652 8542
rect 29708 8428 29764 9996
rect 30156 9938 30212 12460
rect 30716 12514 30772 12526
rect 30716 12462 30718 12514
rect 30770 12462 30772 12514
rect 30604 11844 30660 11854
rect 30716 11844 30772 12462
rect 31052 12402 31108 12414
rect 31052 12350 31054 12402
rect 31106 12350 31108 12402
rect 31052 11954 31108 12350
rect 31052 11902 31054 11954
rect 31106 11902 31108 11954
rect 31052 11890 31108 11902
rect 30604 11842 30772 11844
rect 30604 11790 30606 11842
rect 30658 11790 30772 11842
rect 30604 11788 30772 11790
rect 30604 11778 30660 11788
rect 30828 11732 30884 11742
rect 30380 11620 30436 11630
rect 30380 10724 30436 11564
rect 30380 10630 30436 10668
rect 30828 10722 30884 11676
rect 30828 10670 30830 10722
rect 30882 10670 30884 10722
rect 30828 10658 30884 10670
rect 31164 11730 31220 13804
rect 31612 12740 31668 12750
rect 31612 12626 31668 12684
rect 31612 12574 31614 12626
rect 31666 12574 31668 12626
rect 31612 12562 31668 12574
rect 31724 11954 31780 15598
rect 31836 15652 31892 25452
rect 32508 25060 32564 25070
rect 32508 24966 32564 25004
rect 31948 24836 32004 24846
rect 31948 24500 32004 24780
rect 32396 24724 32452 24734
rect 32172 24722 32452 24724
rect 32172 24670 32398 24722
rect 32450 24670 32452 24722
rect 32172 24668 32452 24670
rect 32060 24500 32116 24510
rect 31948 24498 32116 24500
rect 31948 24446 32062 24498
rect 32114 24446 32116 24498
rect 31948 24444 32116 24446
rect 31948 23604 32004 24444
rect 32060 24434 32116 24444
rect 32060 24052 32116 24062
rect 32172 24052 32228 24668
rect 32396 24658 32452 24668
rect 32620 24724 32676 24734
rect 32620 24630 32676 24668
rect 32060 24050 32228 24052
rect 32060 23998 32062 24050
rect 32114 23998 32228 24050
rect 32060 23996 32228 23998
rect 32844 24498 32900 30492
rect 32956 30546 33012 30558
rect 32956 30494 32958 30546
rect 33010 30494 33012 30546
rect 32956 28756 33012 30494
rect 33516 29874 33572 30604
rect 33628 30658 33684 31892
rect 34076 31890 34132 31892
rect 34076 31838 34078 31890
rect 34130 31838 34132 31890
rect 34076 31826 34132 31838
rect 33852 31778 33908 31790
rect 33852 31726 33854 31778
rect 33906 31726 33908 31778
rect 33852 31220 33908 31726
rect 34300 31778 34356 33404
rect 34636 33394 34692 33404
rect 34412 33010 34468 33022
rect 34412 32958 34414 33010
rect 34466 32958 34468 33010
rect 34412 32788 34468 32958
rect 34748 33010 34804 33740
rect 34748 32958 34750 33010
rect 34802 32958 34804 33010
rect 34748 32946 34804 32958
rect 34860 33794 35140 33796
rect 34860 33742 35086 33794
rect 35138 33742 35140 33794
rect 34860 33740 35140 33742
rect 34860 32788 34916 33740
rect 35084 33730 35140 33740
rect 35308 33794 35364 33806
rect 35308 33742 35310 33794
rect 35362 33742 35364 33794
rect 35308 33684 35364 33742
rect 35308 33618 35364 33628
rect 35196 33292 35460 33302
rect 35252 33236 35300 33292
rect 35356 33236 35404 33292
rect 35196 33226 35460 33236
rect 34412 32732 34916 32788
rect 35084 32676 35140 32686
rect 35532 32676 35588 32686
rect 35084 32674 35532 32676
rect 35084 32622 35086 32674
rect 35138 32622 35532 32674
rect 35084 32620 35532 32622
rect 34300 31726 34302 31778
rect 34354 31726 34356 31778
rect 34300 31714 34356 31726
rect 34636 31892 34692 31902
rect 33740 30884 33796 30894
rect 33740 30790 33796 30828
rect 33852 30770 33908 31164
rect 33852 30718 33854 30770
rect 33906 30718 33908 30770
rect 33852 30706 33908 30718
rect 33964 31442 34020 31454
rect 33964 31390 33966 31442
rect 34018 31390 34020 31442
rect 33628 30606 33630 30658
rect 33682 30606 33684 30658
rect 33628 30548 33684 30606
rect 33628 30482 33684 30492
rect 33964 30212 34020 31390
rect 34636 30658 34692 31836
rect 34748 31668 34804 31678
rect 35084 31668 35140 32620
rect 35532 32582 35588 32620
rect 35644 31892 35700 35084
rect 36204 34804 36260 34814
rect 36204 33906 36260 34748
rect 36988 34802 37044 36876
rect 38332 36818 38388 37660
rect 38332 36766 38334 36818
rect 38386 36766 38388 36818
rect 37548 36706 37604 36718
rect 37548 36654 37550 36706
rect 37602 36654 37604 36706
rect 37100 36596 37156 36606
rect 37548 36596 37604 36654
rect 37100 36594 37604 36596
rect 37100 36542 37102 36594
rect 37154 36542 37604 36594
rect 37100 36540 37604 36542
rect 37100 36146 37156 36540
rect 37100 36094 37102 36146
rect 37154 36094 37156 36146
rect 37100 36082 37156 36094
rect 37100 35924 37156 35934
rect 37100 35830 37156 35868
rect 37548 35812 37604 36540
rect 37772 36708 37828 36718
rect 37772 36036 37828 36652
rect 37660 35812 37716 35822
rect 37548 35810 37716 35812
rect 37548 35758 37662 35810
rect 37714 35758 37716 35810
rect 37548 35756 37716 35758
rect 37772 35812 37828 35980
rect 38332 35924 38388 36766
rect 37884 35812 37940 35822
rect 37772 35810 37940 35812
rect 37772 35758 37886 35810
rect 37938 35758 37940 35810
rect 37772 35756 37940 35758
rect 36988 34750 36990 34802
rect 37042 34750 37044 34802
rect 36988 34738 37044 34750
rect 37212 34804 37268 34814
rect 36540 34020 36596 34030
rect 36540 34018 36932 34020
rect 36540 33966 36542 34018
rect 36594 33966 36932 34018
rect 36540 33964 36932 33966
rect 36540 33954 36596 33964
rect 36204 33854 36206 33906
rect 36258 33854 36260 33906
rect 36204 33842 36260 33854
rect 36876 33906 36932 33964
rect 36876 33854 36878 33906
rect 36930 33854 36932 33906
rect 35644 31826 35700 31836
rect 35756 33012 35812 33022
rect 34748 31666 35140 31668
rect 34748 31614 34750 31666
rect 34802 31614 35140 31666
rect 34748 31612 35140 31614
rect 34748 31602 34804 31612
rect 34636 30606 34638 30658
rect 34690 30606 34692 30658
rect 34636 30594 34692 30606
rect 33964 30146 34020 30156
rect 34188 30548 34244 30558
rect 33516 29822 33518 29874
rect 33570 29822 33572 29874
rect 33516 29810 33572 29822
rect 33852 29876 33908 29886
rect 33852 29782 33908 29820
rect 33628 29764 33684 29774
rect 33180 29650 33236 29662
rect 33180 29598 33182 29650
rect 33234 29598 33236 29650
rect 33180 29540 33236 29598
rect 33628 29540 33684 29708
rect 34188 29762 34244 30492
rect 34300 30546 34356 30558
rect 34300 30494 34302 30546
rect 34354 30494 34356 30546
rect 34300 30324 34356 30494
rect 34300 30258 34356 30268
rect 34748 30324 34804 30334
rect 34748 29986 34804 30268
rect 34748 29934 34750 29986
rect 34802 29934 34804 29986
rect 34748 29922 34804 29934
rect 34188 29710 34190 29762
rect 34242 29710 34244 29762
rect 34188 29698 34244 29710
rect 34748 29764 34804 29774
rect 34860 29764 34916 31612
rect 35644 31556 35700 31566
rect 35196 31276 35460 31286
rect 35252 31220 35300 31276
rect 35356 31220 35404 31276
rect 35196 31210 35460 31220
rect 34972 30884 35028 30894
rect 34972 30770 35028 30828
rect 34972 30718 34974 30770
rect 35026 30718 35028 30770
rect 34972 30706 35028 30718
rect 35196 30770 35252 30782
rect 35196 30718 35198 30770
rect 35250 30718 35252 30770
rect 35084 30548 35140 30558
rect 35084 30454 35140 30492
rect 34804 29708 34916 29764
rect 34972 30436 35028 30446
rect 34748 29698 34804 29708
rect 33852 29652 33908 29662
rect 34972 29652 35028 30380
rect 35084 30324 35140 30334
rect 35084 29986 35140 30268
rect 35084 29934 35086 29986
rect 35138 29934 35140 29986
rect 35084 29922 35140 29934
rect 34972 29596 35140 29652
rect 33852 29558 33908 29596
rect 33236 29484 33684 29540
rect 33180 29446 33236 29484
rect 32956 28690 33012 28700
rect 33292 28754 33348 28766
rect 33292 28702 33294 28754
rect 33346 28702 33348 28754
rect 33068 28530 33124 28542
rect 33068 28478 33070 28530
rect 33122 28478 33124 28530
rect 33068 27858 33124 28478
rect 33292 28532 33348 28702
rect 33628 28756 33684 29484
rect 34972 29428 35028 29438
rect 33852 29426 35028 29428
rect 33852 29374 34974 29426
rect 35026 29374 35028 29426
rect 33852 29372 35028 29374
rect 33740 28756 33796 28766
rect 33628 28754 33796 28756
rect 33628 28702 33742 28754
rect 33794 28702 33796 28754
rect 33628 28700 33796 28702
rect 33292 28466 33348 28476
rect 33516 28644 33572 28654
rect 33516 28082 33572 28588
rect 33516 28030 33518 28082
rect 33570 28030 33572 28082
rect 33516 28018 33572 28030
rect 33068 27806 33070 27858
rect 33122 27806 33124 27858
rect 33068 27794 33124 27806
rect 33404 27860 33460 27870
rect 33404 27766 33460 27804
rect 33516 27858 33572 27870
rect 33516 27806 33518 27858
rect 33570 27806 33572 27858
rect 33404 27412 33460 27422
rect 33292 27076 33348 27086
rect 33068 26740 33124 26750
rect 33068 26646 33124 26684
rect 33292 25842 33348 27020
rect 33292 25790 33294 25842
rect 33346 25790 33348 25842
rect 33292 25778 33348 25790
rect 32844 24446 32846 24498
rect 32898 24446 32900 24498
rect 32060 23986 32116 23996
rect 32060 23604 32116 23614
rect 31948 23548 32060 23604
rect 32060 23538 32116 23548
rect 32620 23604 32676 23614
rect 32508 22484 32564 22494
rect 32508 22390 32564 22428
rect 32060 21586 32116 21598
rect 32060 21534 32062 21586
rect 32114 21534 32116 21586
rect 32060 20132 32116 21534
rect 32060 20066 32116 20076
rect 32508 21588 32564 21598
rect 32620 21588 32676 23548
rect 32508 21586 32676 21588
rect 32508 21534 32510 21586
rect 32562 21534 32676 21586
rect 32508 21532 32676 21534
rect 32172 19572 32228 19582
rect 32060 19010 32116 19022
rect 32060 18958 32062 19010
rect 32114 18958 32116 19010
rect 32060 18674 32116 18958
rect 32060 18622 32062 18674
rect 32114 18622 32116 18674
rect 31948 16772 32004 16782
rect 31948 16436 32004 16716
rect 32060 16658 32116 18622
rect 32172 17892 32228 19516
rect 32508 18676 32564 21532
rect 32844 20468 32900 24446
rect 33292 24498 33348 24510
rect 33292 24446 33294 24498
rect 33346 24446 33348 24498
rect 33180 23940 33236 23950
rect 33292 23940 33348 24446
rect 33180 23938 33348 23940
rect 33180 23886 33182 23938
rect 33234 23886 33348 23938
rect 33180 23884 33348 23886
rect 33180 23874 33236 23884
rect 32956 23828 33012 23838
rect 32956 22818 33012 23772
rect 33292 23716 33348 23884
rect 33292 23650 33348 23660
rect 32956 22766 32958 22818
rect 33010 22766 33012 22818
rect 32956 22754 33012 22766
rect 33292 22594 33348 22606
rect 33292 22542 33294 22594
rect 33346 22542 33348 22594
rect 33292 22484 33348 22542
rect 33292 22418 33348 22428
rect 33404 22260 33460 27356
rect 33516 26850 33572 27806
rect 33740 27636 33796 28700
rect 33740 27570 33796 27580
rect 33852 27858 33908 29372
rect 34972 29362 35028 29372
rect 35084 29204 35140 29596
rect 35196 29428 35252 30718
rect 35420 30772 35476 30782
rect 35420 30770 35588 30772
rect 35420 30718 35422 30770
rect 35474 30718 35588 30770
rect 35420 30716 35588 30718
rect 35420 30706 35476 30716
rect 35532 30324 35588 30716
rect 35644 30770 35700 31500
rect 35756 31108 35812 32956
rect 36876 32228 36932 33854
rect 37212 34018 37268 34748
rect 37660 34580 37716 35756
rect 37884 35700 37940 35756
rect 38332 35810 38388 35868
rect 38332 35758 38334 35810
rect 38386 35758 38388 35810
rect 38332 35746 38388 35758
rect 37884 35644 38276 35700
rect 38108 34804 38164 34814
rect 38108 34710 38164 34748
rect 37660 34514 37716 34524
rect 37324 34468 37380 34478
rect 37996 34468 38052 34478
rect 37324 34466 37492 34468
rect 37324 34414 37326 34466
rect 37378 34414 37492 34466
rect 37324 34412 37492 34414
rect 37324 34402 37380 34412
rect 37212 33966 37214 34018
rect 37266 33966 37268 34018
rect 37212 33908 37268 33966
rect 37212 33842 37268 33852
rect 37100 32676 37156 32686
rect 37100 32582 37156 32620
rect 37324 32564 37380 32574
rect 36876 32172 37156 32228
rect 36652 31780 36708 31790
rect 35756 31042 35812 31052
rect 35980 31666 36036 31678
rect 35980 31614 35982 31666
rect 36034 31614 36036 31666
rect 35644 30718 35646 30770
rect 35698 30718 35700 30770
rect 35644 30706 35700 30718
rect 35980 30324 36036 31614
rect 36652 30996 36708 31724
rect 37100 31780 37156 32172
rect 37324 31890 37380 32508
rect 37324 31838 37326 31890
rect 37378 31838 37380 31890
rect 37324 31826 37380 31838
rect 37100 31778 37268 31780
rect 37100 31726 37102 31778
rect 37154 31726 37268 31778
rect 37100 31724 37268 31726
rect 37100 31714 37156 31724
rect 37212 31668 37268 31724
rect 37324 31668 37380 31678
rect 37212 31666 37380 31668
rect 37212 31614 37326 31666
rect 37378 31614 37380 31666
rect 37212 31612 37380 31614
rect 37324 31602 37380 31612
rect 36988 31556 37044 31566
rect 36988 31462 37044 31500
rect 36428 30772 36484 30782
rect 36428 30658 36484 30716
rect 36428 30606 36430 30658
rect 36482 30606 36484 30658
rect 36428 30594 36484 30606
rect 35532 30268 36036 30324
rect 36092 30546 36148 30558
rect 36092 30494 36094 30546
rect 36146 30494 36148 30546
rect 35420 30212 35476 30222
rect 35420 29762 35476 30156
rect 35420 29710 35422 29762
rect 35474 29710 35476 29762
rect 35420 29698 35476 29710
rect 35644 29764 35700 29774
rect 35868 29768 35924 30268
rect 36092 29988 36148 30494
rect 36092 29922 36148 29932
rect 36204 30436 36260 30446
rect 35644 29762 35812 29764
rect 35644 29710 35646 29762
rect 35698 29710 35812 29762
rect 35644 29708 35812 29710
rect 35644 29698 35700 29708
rect 35196 29372 35588 29428
rect 34972 29148 35140 29204
rect 35196 29260 35460 29270
rect 35252 29204 35300 29260
rect 35356 29204 35404 29260
rect 35196 29194 35460 29204
rect 34748 28980 34804 28990
rect 34300 28756 34356 28766
rect 34300 28662 34356 28700
rect 34524 28754 34580 28766
rect 34524 28702 34526 28754
rect 34578 28702 34580 28754
rect 34524 28644 34580 28702
rect 34748 28754 34804 28924
rect 34748 28702 34750 28754
rect 34802 28702 34804 28754
rect 34748 28690 34804 28702
rect 34972 28754 35028 29148
rect 35532 29092 35588 29372
rect 35420 29036 35588 29092
rect 34972 28702 34974 28754
rect 35026 28702 35028 28754
rect 34972 28690 35028 28702
rect 35084 28978 35140 28990
rect 35084 28926 35086 28978
rect 35138 28926 35140 28978
rect 35084 28756 35140 28926
rect 35308 28756 35364 28766
rect 35084 28754 35364 28756
rect 35084 28702 35310 28754
rect 35362 28702 35364 28754
rect 35084 28700 35364 28702
rect 35308 28690 35364 28700
rect 34524 28578 34580 28588
rect 33852 27806 33854 27858
rect 33906 27806 33908 27858
rect 33516 26798 33518 26850
rect 33570 26798 33572 26850
rect 33516 26786 33572 26798
rect 33740 26740 33796 26750
rect 33740 26646 33796 26684
rect 33628 25508 33684 25518
rect 33628 25414 33684 25452
rect 33852 25396 33908 27806
rect 34412 27970 34468 27982
rect 34412 27918 34414 27970
rect 34466 27918 34468 27970
rect 34188 27746 34244 27758
rect 34188 27694 34190 27746
rect 34242 27694 34244 27746
rect 34188 26908 34244 27694
rect 33852 25330 33908 25340
rect 33964 26852 34244 26908
rect 34412 27636 34468 27918
rect 35420 27636 35476 29036
rect 35644 28754 35700 28766
rect 35644 28702 35646 28754
rect 35698 28702 35700 28754
rect 35532 28642 35588 28654
rect 35532 28590 35534 28642
rect 35586 28590 35588 28642
rect 35532 28196 35588 28590
rect 35532 28130 35588 28140
rect 35644 28084 35700 28702
rect 35756 28084 35812 29708
rect 35868 29716 35870 29768
rect 35922 29764 35924 29768
rect 35980 29764 36036 29774
rect 35922 29716 35980 29764
rect 35868 29708 35980 29716
rect 35868 29704 35924 29708
rect 35980 29698 36036 29708
rect 36092 29764 36148 29774
rect 36204 29764 36260 30380
rect 36652 30324 36708 30940
rect 37324 30996 37380 31006
rect 36988 30884 37044 30894
rect 36988 30790 37044 30828
rect 37324 30770 37380 30940
rect 37324 30718 37326 30770
rect 37378 30718 37380 30770
rect 37324 30706 37380 30718
rect 36652 30258 36708 30268
rect 37324 30324 37380 30334
rect 37100 29988 37156 29998
rect 36652 29764 36708 29774
rect 36092 29762 36260 29764
rect 36092 29710 36094 29762
rect 36146 29710 36260 29762
rect 36092 29708 36260 29710
rect 36428 29762 36708 29764
rect 36428 29710 36654 29762
rect 36706 29710 36708 29762
rect 36428 29708 36708 29710
rect 36092 29698 36148 29708
rect 35980 29428 36036 29438
rect 35980 28644 36036 29372
rect 36204 29426 36260 29438
rect 36204 29374 36206 29426
rect 36258 29374 36260 29426
rect 36204 29316 36260 29374
rect 36204 29250 36260 29260
rect 36428 29204 36484 29708
rect 36652 29698 36708 29708
rect 36876 29762 36932 29774
rect 36876 29710 36878 29762
rect 36930 29710 36932 29762
rect 36764 29652 36820 29662
rect 36764 29558 36820 29596
rect 36876 29540 36932 29710
rect 37100 29762 37156 29932
rect 37100 29710 37102 29762
rect 37154 29710 37156 29762
rect 37100 29698 37156 29710
rect 37324 29762 37380 30268
rect 37324 29710 37326 29762
rect 37378 29710 37380 29762
rect 37324 29698 37380 29710
rect 37436 29540 37492 34412
rect 37884 34466 38052 34468
rect 37884 34414 37998 34466
rect 38050 34414 38052 34466
rect 37884 34412 38052 34414
rect 37548 32562 37604 32574
rect 37548 32510 37550 32562
rect 37602 32510 37604 32562
rect 37548 31668 37604 32510
rect 37772 31668 37828 31678
rect 37548 31612 37772 31668
rect 37772 31574 37828 31612
rect 37660 31442 37716 31454
rect 37660 31390 37662 31442
rect 37714 31390 37716 31442
rect 37660 30882 37716 31390
rect 37884 30884 37940 34412
rect 37996 34402 38052 34412
rect 37996 33684 38052 33694
rect 38220 33684 38276 35644
rect 38332 35588 38388 35598
rect 38332 34802 38388 35532
rect 38332 34750 38334 34802
rect 38386 34750 38388 34802
rect 38332 34738 38388 34750
rect 38332 34020 38388 34030
rect 38332 33684 38388 33964
rect 37996 33682 38388 33684
rect 37996 33630 37998 33682
rect 38050 33630 38388 33682
rect 37996 33628 38388 33630
rect 37996 33618 38052 33628
rect 38220 32786 38276 32798
rect 38220 32734 38222 32786
rect 38274 32734 38276 32786
rect 38220 31668 38276 32734
rect 38332 32786 38388 33628
rect 38332 32734 38334 32786
rect 38386 32734 38388 32786
rect 38332 32722 38388 32734
rect 38444 31948 38500 39902
rect 38780 39842 38836 40796
rect 38892 40850 38948 41916
rect 38892 40798 38894 40850
rect 38946 40798 38948 40850
rect 38892 40786 38948 40798
rect 39228 40068 39284 42700
rect 39564 41970 39620 41982
rect 39564 41918 39566 41970
rect 39618 41918 39620 41970
rect 39564 40852 39620 41918
rect 39788 41972 39844 41982
rect 39844 41916 39956 41972
rect 39788 41906 39844 41916
rect 39900 41858 39956 41916
rect 39900 41806 39902 41858
rect 39954 41806 39956 41858
rect 39900 41794 39956 41806
rect 39564 40786 39620 40796
rect 39676 40738 39732 40750
rect 39676 40686 39678 40738
rect 39730 40686 39732 40738
rect 39228 40002 39284 40012
rect 39564 40626 39620 40638
rect 39564 40574 39566 40626
rect 39618 40574 39620 40626
rect 38780 39790 38782 39842
rect 38834 39790 38836 39842
rect 38780 39620 38836 39790
rect 38780 39554 38836 39564
rect 39564 39508 39620 40574
rect 39676 40516 39732 40686
rect 39676 40450 39732 40460
rect 39788 39956 39844 39966
rect 39788 39732 39844 39900
rect 39788 39638 39844 39676
rect 39564 39452 39844 39508
rect 39452 39060 39508 39070
rect 38556 38948 38612 38958
rect 38556 38834 38612 38892
rect 38556 38782 38558 38834
rect 38610 38782 38612 38834
rect 38556 38770 38612 38782
rect 39116 38836 39172 38846
rect 39116 38742 39172 38780
rect 39452 38836 39508 39004
rect 38556 37940 38612 37950
rect 38556 37604 38612 37884
rect 38892 37940 38948 37950
rect 38892 37846 38948 37884
rect 38556 36708 38612 37548
rect 39452 36820 39508 38780
rect 39788 38722 39844 39452
rect 39788 38670 39790 38722
rect 39842 38670 39844 38722
rect 39788 38658 39844 38670
rect 40124 37828 40180 43484
rect 40236 42756 40292 44606
rect 40796 44212 40852 44222
rect 40460 44210 40852 44212
rect 40460 44158 40798 44210
rect 40850 44158 40852 44210
rect 40460 44156 40852 44158
rect 40348 43764 40404 43774
rect 40348 43650 40404 43708
rect 40348 43598 40350 43650
rect 40402 43598 40404 43650
rect 40348 43586 40404 43598
rect 40460 43204 40516 44156
rect 40796 44146 40852 44156
rect 40796 43540 40852 43550
rect 40908 43540 40964 44716
rect 41020 43764 41076 43774
rect 41244 43764 41300 45836
rect 41356 45826 41412 45836
rect 41580 45890 41636 47630
rect 41580 45838 41582 45890
rect 41634 45838 41636 45890
rect 41580 45826 41636 45838
rect 41804 45890 41860 48076
rect 41916 47794 41972 47806
rect 41916 47742 41918 47794
rect 41970 47742 41972 47794
rect 41916 47570 41972 47742
rect 42364 47794 42420 47806
rect 42364 47742 42366 47794
rect 42418 47742 42420 47794
rect 42364 47682 42420 47742
rect 42364 47630 42366 47682
rect 42418 47630 42420 47682
rect 42364 47618 42420 47630
rect 42812 47794 42868 47806
rect 42812 47742 42814 47794
rect 42866 47742 42868 47794
rect 41916 47518 41918 47570
rect 41970 47518 41972 47570
rect 41916 47506 41972 47518
rect 42812 47570 42868 47742
rect 43260 47794 43316 47806
rect 43260 47742 43262 47794
rect 43314 47742 43316 47794
rect 42812 47518 42814 47570
rect 42866 47518 42868 47570
rect 42812 47506 42868 47518
rect 43148 47684 43204 47694
rect 43260 47684 43316 47742
rect 43148 47682 43316 47684
rect 43148 47630 43150 47682
rect 43202 47630 43316 47682
rect 43148 47628 43316 47630
rect 43148 47010 43204 47628
rect 43148 46958 43150 47010
rect 43202 46958 43204 47010
rect 41916 46674 41972 46686
rect 41916 46622 41918 46674
rect 41970 46622 41972 46674
rect 41916 46226 41972 46622
rect 42700 46676 42756 46686
rect 42700 46674 42868 46676
rect 42700 46622 42702 46674
rect 42754 46622 42868 46674
rect 42700 46620 42868 46622
rect 42700 46610 42756 46620
rect 41916 46174 41918 46226
rect 41970 46174 41972 46226
rect 41916 46162 41972 46174
rect 41804 45838 41806 45890
rect 41858 45838 41860 45890
rect 41804 45826 41860 45838
rect 42812 46004 42868 46620
rect 43148 46562 43204 46958
rect 43148 46510 43150 46562
rect 43202 46510 43204 46562
rect 43148 46498 43204 46510
rect 43372 46676 43428 48076
rect 43596 47012 43652 47022
rect 43708 47012 43764 48748
rect 50556 48412 50820 48422
rect 50612 48356 50660 48412
rect 50716 48356 50764 48412
rect 50556 48346 50820 48356
rect 43596 47010 43764 47012
rect 43596 46958 43598 47010
rect 43650 46958 43764 47010
rect 43596 46956 43764 46958
rect 43596 46946 43652 46956
rect 42812 45890 42868 45948
rect 42812 45838 42814 45890
rect 42866 45838 42868 45890
rect 42140 45444 42196 45454
rect 41356 44770 41412 44782
rect 41356 44718 41358 44770
rect 41410 44718 41412 44770
rect 41356 44210 41412 44718
rect 41356 44158 41358 44210
rect 41410 44158 41412 44210
rect 41356 44146 41412 44158
rect 42028 44658 42084 44670
rect 42028 44606 42030 44658
rect 42082 44606 42084 44658
rect 41468 43764 41524 43774
rect 41076 43708 41300 43764
rect 41356 43708 41468 43764
rect 41020 43670 41076 43708
rect 40852 43484 40964 43540
rect 40796 43474 40852 43484
rect 41356 43204 41412 43708
rect 41468 43670 41524 43708
rect 41692 43540 41748 43550
rect 41692 43538 41860 43540
rect 41692 43486 41694 43538
rect 41746 43486 41860 43538
rect 41692 43484 41860 43486
rect 41692 43474 41748 43484
rect 40236 42690 40292 42700
rect 40348 43148 40516 43204
rect 41020 43148 41412 43204
rect 40348 41746 40404 43148
rect 41020 42868 41076 43148
rect 40348 41694 40350 41746
rect 40402 41694 40404 41746
rect 40348 41682 40404 41694
rect 40460 42754 40516 42766
rect 40460 42702 40462 42754
rect 40514 42702 40516 42754
rect 40348 40740 40404 40750
rect 40236 40068 40292 40078
rect 40236 39730 40292 40012
rect 40236 39678 40238 39730
rect 40290 39678 40292 39730
rect 40236 39060 40292 39678
rect 40236 38994 40292 39004
rect 40236 38724 40292 38734
rect 40236 38162 40292 38668
rect 40236 38110 40238 38162
rect 40290 38110 40292 38162
rect 40236 38098 40292 38110
rect 40124 37772 40292 37828
rect 39452 36818 39620 36820
rect 39452 36766 39454 36818
rect 39506 36766 39620 36818
rect 39452 36764 39620 36766
rect 39452 36754 39508 36764
rect 38556 36642 38612 36652
rect 38668 36708 38724 36718
rect 39116 36708 39172 36718
rect 38668 36706 39172 36708
rect 38668 36654 38670 36706
rect 38722 36654 39118 36706
rect 39170 36654 39172 36706
rect 38668 36652 39172 36654
rect 38668 36642 38724 36652
rect 39116 36642 39172 36652
rect 38892 36484 38948 36494
rect 38668 34804 38724 34842
rect 38668 34738 38724 34748
rect 38892 34802 38948 36428
rect 39564 35028 39620 36764
rect 39788 36706 39844 36718
rect 39788 36654 39790 36706
rect 39842 36654 39844 36706
rect 39676 36036 39732 36046
rect 39788 36036 39844 36654
rect 39676 36034 39844 36036
rect 39676 35982 39678 36034
rect 39730 35982 39844 36034
rect 39676 35980 39844 35982
rect 40124 36594 40180 36606
rect 40124 36542 40126 36594
rect 40178 36542 40180 36594
rect 39676 35970 39732 35980
rect 40012 35586 40068 35598
rect 40012 35534 40014 35586
rect 40066 35534 40068 35586
rect 39676 35028 39732 35038
rect 39564 35026 39732 35028
rect 39564 34974 39678 35026
rect 39730 34974 39732 35026
rect 39564 34972 39732 34974
rect 39676 34962 39732 34972
rect 38892 34750 38894 34802
rect 38946 34750 38948 34802
rect 38892 34738 38948 34750
rect 40012 34690 40068 35534
rect 40124 35588 40180 36542
rect 40124 35522 40180 35532
rect 40012 34638 40014 34690
rect 40066 34638 40068 34690
rect 38668 34578 38724 34590
rect 38668 34526 38670 34578
rect 38722 34526 38724 34578
rect 38668 33684 38724 34526
rect 38668 33628 38836 33684
rect 38780 31948 38836 33628
rect 39788 32788 39844 32798
rect 39788 32694 39844 32732
rect 38220 31602 38276 31612
rect 38332 31892 38500 31948
rect 38668 31892 38836 31948
rect 38892 32676 38948 32686
rect 37660 30830 37662 30882
rect 37714 30830 37716 30882
rect 37660 30818 37716 30830
rect 37772 30828 37940 30884
rect 38108 31442 38164 31454
rect 38108 31390 38110 31442
rect 38162 31390 38164 31442
rect 38108 30884 38164 31390
rect 38220 30884 38276 30894
rect 38108 30882 38276 30884
rect 38108 30830 38222 30882
rect 38274 30830 38276 30882
rect 38108 30828 38276 30830
rect 37548 30548 37604 30558
rect 37548 30454 37604 30492
rect 37772 30324 37828 30828
rect 38220 30818 38276 30828
rect 37996 30772 38052 30782
rect 37772 30258 37828 30268
rect 37884 30658 37940 30670
rect 37884 30606 37886 30658
rect 37938 30606 37940 30658
rect 36876 29484 37044 29540
rect 36652 29316 36708 29326
rect 36708 29260 36932 29316
rect 36652 29250 36708 29260
rect 36428 29148 36596 29204
rect 36428 28980 36484 28990
rect 36428 28866 36484 28924
rect 36428 28814 36430 28866
rect 36482 28814 36484 28866
rect 36428 28802 36484 28814
rect 35980 28550 36036 28588
rect 36540 28420 36596 29148
rect 36876 28754 36932 29260
rect 36876 28702 36878 28754
rect 36930 28702 36932 28754
rect 36876 28690 36932 28702
rect 36988 28532 37044 29484
rect 37324 29484 37492 29540
rect 37548 29988 37604 29998
rect 37100 28868 37156 28878
rect 37100 28774 37156 28812
rect 36540 28354 36596 28364
rect 36652 28476 37044 28532
rect 37212 28754 37268 28766
rect 37212 28702 37214 28754
rect 37266 28702 37268 28754
rect 36204 28084 36260 28094
rect 35756 28082 36260 28084
rect 35756 28030 36206 28082
rect 36258 28030 36260 28082
rect 35756 28028 36260 28030
rect 35644 28018 35700 28028
rect 36204 28018 36260 28028
rect 35532 27860 35588 27870
rect 35980 27860 36036 27870
rect 35532 27858 36036 27860
rect 35532 27806 35534 27858
rect 35586 27806 35982 27858
rect 36034 27806 36036 27858
rect 35532 27804 36036 27806
rect 35532 27794 35588 27804
rect 35980 27794 36036 27804
rect 36316 27860 36372 27870
rect 36316 27766 36372 27804
rect 36540 27858 36596 27870
rect 36540 27806 36542 27858
rect 36594 27806 36596 27858
rect 35980 27636 36036 27646
rect 35420 27580 35812 27636
rect 33964 25508 34020 26852
rect 34188 26738 34244 26750
rect 34188 26686 34190 26738
rect 34242 26686 34244 26738
rect 34188 26628 34244 26686
rect 34188 26562 34244 26572
rect 34412 25956 34468 27580
rect 35644 27412 35700 27422
rect 35532 27356 35644 27412
rect 35196 27244 35460 27254
rect 35252 27188 35300 27244
rect 35356 27188 35404 27244
rect 35196 27178 35460 27188
rect 35308 26964 35364 26974
rect 35532 26964 35588 27356
rect 35644 27346 35700 27356
rect 35308 26962 35588 26964
rect 35308 26910 35310 26962
rect 35362 26910 35588 26962
rect 35308 26908 35588 26910
rect 35308 26898 35364 26908
rect 34748 26738 34804 26750
rect 34748 26686 34750 26738
rect 34802 26686 34804 26738
rect 34748 26628 34804 26686
rect 35084 26740 35140 26750
rect 35644 26740 35700 26750
rect 35084 26738 35700 26740
rect 35084 26686 35086 26738
rect 35138 26686 35646 26738
rect 35698 26686 35700 26738
rect 35084 26684 35700 26686
rect 35084 26674 35140 26684
rect 35644 26674 35700 26684
rect 34748 26562 34804 26572
rect 35756 26066 35812 27580
rect 35980 26628 36036 27580
rect 36540 27412 36596 27806
rect 36540 27346 36596 27356
rect 36652 27188 36708 28476
rect 37212 27972 37268 28702
rect 37100 27916 37268 27972
rect 35756 26014 35758 26066
rect 35810 26014 35812 26066
rect 35756 26002 35812 26014
rect 35868 26626 36036 26628
rect 35868 26574 35982 26626
rect 36034 26574 36036 26626
rect 35868 26572 36036 26574
rect 34076 25900 34468 25956
rect 34076 25730 34132 25900
rect 34076 25678 34078 25730
rect 34130 25678 34132 25730
rect 34076 25666 34132 25678
rect 34188 25730 34244 25742
rect 34188 25678 34190 25730
rect 34242 25678 34244 25730
rect 34188 25508 34244 25678
rect 33964 25452 34244 25508
rect 33964 24836 34020 25452
rect 33740 24500 33796 24510
rect 33964 24500 34020 24780
rect 33740 24498 34020 24500
rect 33740 24446 33742 24498
rect 33794 24446 34020 24498
rect 33740 24444 34020 24446
rect 33740 24434 33796 24444
rect 33740 23716 33796 23726
rect 33740 23622 33796 23660
rect 33964 23716 34020 24444
rect 34188 24836 34244 24846
rect 34412 24836 34468 25900
rect 35532 25844 35588 25854
rect 35756 25844 35812 25854
rect 35532 25750 35588 25788
rect 35644 25842 35812 25844
rect 35644 25790 35758 25842
rect 35810 25790 35812 25842
rect 35644 25788 35812 25790
rect 34524 25730 34580 25742
rect 34524 25678 34526 25730
rect 34578 25678 34580 25730
rect 34524 25060 34580 25678
rect 34860 25732 34916 25742
rect 35196 25732 35252 25742
rect 34860 25730 35252 25732
rect 34860 25678 34862 25730
rect 34914 25678 35198 25730
rect 35250 25678 35252 25730
rect 34860 25676 35252 25678
rect 34860 25666 34916 25676
rect 35196 25666 35252 25676
rect 34524 24994 34580 25004
rect 34860 25396 34916 25406
rect 35644 25396 35700 25788
rect 35756 25778 35812 25788
rect 34188 24834 34468 24836
rect 34188 24782 34190 24834
rect 34242 24782 34468 24834
rect 34188 24780 34468 24782
rect 34188 23938 34244 24780
rect 34860 24610 34916 25340
rect 34860 24558 34862 24610
rect 34914 24558 34916 24610
rect 34860 24546 34916 24558
rect 35084 25340 35700 25396
rect 34524 24500 34580 24510
rect 34524 24406 34580 24444
rect 34188 23886 34190 23938
rect 34242 23886 34244 23938
rect 34188 23874 34244 23886
rect 34300 23940 34356 23950
rect 34300 23938 34804 23940
rect 34300 23886 34302 23938
rect 34354 23886 34804 23938
rect 34300 23884 34804 23886
rect 34300 23874 34356 23884
rect 33964 23714 34132 23716
rect 33964 23662 33966 23714
rect 34018 23662 34132 23714
rect 33964 23660 34132 23662
rect 33964 23650 34020 23660
rect 34076 23604 34132 23660
rect 33628 23042 33684 23054
rect 33628 22990 33630 23042
rect 33682 22990 33684 23042
rect 33628 22482 33684 22990
rect 34076 22818 34132 23548
rect 34076 22766 34078 22818
rect 34130 22766 34132 22818
rect 34076 22754 34132 22766
rect 34412 23714 34468 23726
rect 34412 23662 34414 23714
rect 34466 23662 34468 23714
rect 34412 23042 34468 23662
rect 34748 23714 34804 23884
rect 35084 23938 35140 25340
rect 35196 25228 35460 25238
rect 35252 25172 35300 25228
rect 35356 25172 35404 25228
rect 35196 25162 35460 25172
rect 35084 23886 35086 23938
rect 35138 23886 35140 23938
rect 35084 23874 35140 23886
rect 35196 25060 35252 25070
rect 35196 24722 35252 25004
rect 35196 24670 35198 24722
rect 35250 24670 35252 24722
rect 34748 23662 34750 23714
rect 34802 23662 34804 23714
rect 34748 23650 34804 23662
rect 35196 23716 35252 24670
rect 35644 24836 35700 24846
rect 35644 24722 35700 24780
rect 35868 24724 35924 26572
rect 35980 26562 36036 26572
rect 36092 27132 36708 27188
rect 36764 27858 36820 27870
rect 36764 27806 36766 27858
rect 36818 27806 36820 27858
rect 35980 26068 36036 26078
rect 35980 25842 36036 26012
rect 35980 25790 35982 25842
rect 36034 25790 36036 25842
rect 35980 25778 36036 25790
rect 35644 24670 35646 24722
rect 35698 24670 35700 24722
rect 35644 24658 35700 24670
rect 35756 24722 35924 24724
rect 35756 24670 35870 24722
rect 35922 24670 35924 24722
rect 35756 24668 35924 24670
rect 35420 24500 35476 24510
rect 35420 23826 35476 24444
rect 35756 24052 35812 24668
rect 35868 24658 35924 24668
rect 35420 23774 35422 23826
rect 35474 23774 35476 23826
rect 35420 23762 35476 23774
rect 35644 23996 35812 24052
rect 35868 24164 35924 24174
rect 35196 23492 35252 23660
rect 35196 23436 35588 23492
rect 35196 23212 35460 23222
rect 35252 23156 35300 23212
rect 35356 23156 35404 23212
rect 35196 23146 35460 23156
rect 34412 22990 34414 23042
rect 34466 22990 34468 23042
rect 34412 22820 34468 22990
rect 34412 22754 34468 22764
rect 35420 22708 35476 22718
rect 35532 22708 35588 23436
rect 35644 23042 35700 23996
rect 35868 23938 35924 24108
rect 36092 24050 36148 27132
rect 36316 26852 36372 26862
rect 36316 26850 36596 26852
rect 36316 26798 36318 26850
rect 36370 26798 36596 26850
rect 36316 26796 36596 26798
rect 36316 26786 36372 26796
rect 36540 26404 36596 26796
rect 36540 25730 36596 26348
rect 36764 26068 36820 27806
rect 36988 27636 37044 27646
rect 36988 26908 37044 27580
rect 37100 27076 37156 27916
rect 37324 27746 37380 29484
rect 37436 28644 37492 28654
rect 37436 28550 37492 28588
rect 37324 27694 37326 27746
rect 37378 27694 37380 27746
rect 37324 27682 37380 27694
rect 37548 27746 37604 29932
rect 37884 29988 37940 30606
rect 37996 30212 38052 30716
rect 38332 30548 38388 31892
rect 38444 31780 38500 31790
rect 38444 30770 38500 31724
rect 38556 31668 38612 31678
rect 38556 31574 38612 31612
rect 38444 30718 38446 30770
rect 38498 30718 38500 30770
rect 38444 30706 38500 30718
rect 38556 30996 38612 31006
rect 38556 30548 38612 30940
rect 38332 30492 38500 30548
rect 38108 30436 38164 30446
rect 38108 30342 38164 30380
rect 37996 30156 38276 30212
rect 37884 29922 37940 29932
rect 38220 29986 38276 30156
rect 38220 29934 38222 29986
rect 38274 29934 38276 29986
rect 38220 29922 38276 29934
rect 38332 29876 38388 29886
rect 38332 29782 38388 29820
rect 37884 29764 37940 29774
rect 37884 29670 37940 29708
rect 38444 28978 38500 30492
rect 38556 30482 38612 30492
rect 38444 28926 38446 28978
rect 38498 28926 38500 28978
rect 38444 28866 38500 28926
rect 38444 28814 38446 28866
rect 38498 28814 38500 28866
rect 38444 28802 38500 28814
rect 38668 28756 38724 31892
rect 38780 30996 38836 31006
rect 38892 30996 38948 32620
rect 39116 32676 39172 32686
rect 39452 32676 39508 32686
rect 39116 32674 39508 32676
rect 39116 32622 39118 32674
rect 39170 32622 39454 32674
rect 39506 32622 39508 32674
rect 39116 32620 39508 32622
rect 39116 32610 39172 32620
rect 39452 32610 39508 32620
rect 39004 31892 39060 31902
rect 39004 31778 39060 31836
rect 39004 31726 39006 31778
rect 39058 31726 39060 31778
rect 39004 31714 39060 31726
rect 38780 30994 38948 30996
rect 38780 30942 38782 30994
rect 38834 30942 38948 30994
rect 38780 30940 38948 30942
rect 39900 31668 39956 31678
rect 38780 30930 38836 30940
rect 38556 28700 38724 28756
rect 39004 30884 39060 30894
rect 39004 30660 39060 30828
rect 39116 30660 39172 30670
rect 39452 30660 39508 30670
rect 39004 30658 39172 30660
rect 39004 30606 39118 30658
rect 39170 30606 39172 30658
rect 39004 30604 39172 30606
rect 37996 28532 38052 28542
rect 37996 28438 38052 28476
rect 37884 28084 37940 28094
rect 37884 27970 37940 28028
rect 37884 27918 37886 27970
rect 37938 27918 37940 27970
rect 37884 27906 37940 27918
rect 37772 27748 37828 27758
rect 37548 27694 37550 27746
rect 37602 27694 37604 27746
rect 37436 27076 37492 27086
rect 37100 27074 37492 27076
rect 37100 27022 37438 27074
rect 37490 27022 37492 27074
rect 37100 27020 37492 27022
rect 37436 27010 37492 27020
rect 36764 26002 36820 26012
rect 36876 26852 37044 26908
rect 37212 26852 37268 26862
rect 36764 25844 36820 25854
rect 36876 25844 36932 26852
rect 37100 26740 37156 26750
rect 37100 26646 37156 26684
rect 36764 25842 36932 25844
rect 36764 25790 36766 25842
rect 36818 25790 36932 25842
rect 36764 25788 36932 25790
rect 36764 25778 36820 25788
rect 36540 25678 36542 25730
rect 36594 25678 36596 25730
rect 36204 24948 36260 24958
rect 36204 24498 36260 24892
rect 36540 24836 36596 25678
rect 36540 24770 36596 24780
rect 36652 25730 36708 25742
rect 36652 25678 36654 25730
rect 36706 25678 36708 25730
rect 36204 24446 36206 24498
rect 36258 24446 36260 24498
rect 36204 24434 36260 24446
rect 36092 23998 36094 24050
rect 36146 23998 36148 24050
rect 36092 23986 36148 23998
rect 35868 23886 35870 23938
rect 35922 23886 35924 23938
rect 35868 23874 35924 23886
rect 35644 22990 35646 23042
rect 35698 22990 35700 23042
rect 35644 22978 35700 22990
rect 35756 23826 35812 23838
rect 35756 23774 35758 23826
rect 35810 23774 35812 23826
rect 35756 22932 35812 23774
rect 36540 23828 36596 23838
rect 36652 23828 36708 25678
rect 36988 25730 37044 25742
rect 36988 25678 36990 25730
rect 37042 25678 37044 25730
rect 36988 25284 37044 25678
rect 37212 25730 37268 26796
rect 37212 25678 37214 25730
rect 37266 25678 37268 25730
rect 37212 25666 37268 25678
rect 37324 26738 37380 26750
rect 37324 26686 37326 26738
rect 37378 26686 37380 26738
rect 36988 25218 37044 25228
rect 36764 24948 36820 24958
rect 36820 24892 36932 24948
rect 36764 24882 36820 24892
rect 36876 24722 36932 24892
rect 36876 24670 36878 24722
rect 36930 24670 36932 24722
rect 36876 24658 36932 24670
rect 37212 24498 37268 24510
rect 37212 24446 37214 24498
rect 37266 24446 37268 24498
rect 37212 24388 37268 24446
rect 36764 24332 37212 24388
rect 36764 24164 36820 24332
rect 37212 24294 37268 24332
rect 36764 23938 36820 24108
rect 36988 24052 37044 24062
rect 37324 24052 37380 26686
rect 37548 26738 37604 27694
rect 37548 26686 37550 26738
rect 37602 26686 37604 26738
rect 37548 26516 37604 26686
rect 37548 26450 37604 26460
rect 37660 27746 37828 27748
rect 37660 27694 37774 27746
rect 37826 27694 37828 27746
rect 37660 27692 37828 27694
rect 37660 26068 37716 27692
rect 37772 27682 37828 27692
rect 37996 27746 38052 27758
rect 37996 27694 37998 27746
rect 38050 27694 38052 27746
rect 37772 27412 37828 27422
rect 37772 26738 37828 27356
rect 37772 26686 37774 26738
rect 37826 26686 37828 26738
rect 37772 26674 37828 26686
rect 37436 26012 37716 26068
rect 37772 26068 37828 26078
rect 37436 24386 37492 26012
rect 37772 25956 37828 26012
rect 37996 26068 38052 27694
rect 38444 27636 38500 27646
rect 38444 27542 38500 27580
rect 38556 27412 38612 28700
rect 38892 28530 38948 28542
rect 38892 28478 38894 28530
rect 38946 28478 38948 28530
rect 38668 28420 38724 28430
rect 38724 28364 38836 28420
rect 38668 28354 38724 28364
rect 38556 27346 38612 27356
rect 38668 27860 38724 27870
rect 38668 26964 38724 27804
rect 38556 26908 38724 26964
rect 38780 26964 38836 28364
rect 38892 27748 38948 28478
rect 38892 27300 38948 27692
rect 39004 27524 39060 30604
rect 39116 30594 39172 30604
rect 39228 30604 39452 30660
rect 39228 30548 39284 30604
rect 39452 30566 39508 30604
rect 39228 29986 39284 30492
rect 39228 29934 39230 29986
rect 39282 29934 39284 29986
rect 39228 29922 39284 29934
rect 39788 30546 39844 30558
rect 39788 30494 39790 30546
rect 39842 30494 39844 30546
rect 39788 30212 39844 30494
rect 39676 29652 39732 29662
rect 39340 28756 39396 28766
rect 39676 28756 39732 29596
rect 39788 29092 39844 30156
rect 39788 29026 39844 29036
rect 39900 30098 39956 31612
rect 39900 30046 39902 30098
rect 39954 30046 39956 30098
rect 39900 29650 39956 30046
rect 39900 29598 39902 29650
rect 39954 29598 39956 29650
rect 39340 28754 39732 28756
rect 39340 28702 39342 28754
rect 39394 28702 39732 28754
rect 39340 28700 39732 28702
rect 39340 28690 39396 28700
rect 39452 28532 39508 28542
rect 39228 28418 39284 28430
rect 39228 28366 39230 28418
rect 39282 28366 39284 28418
rect 39228 27970 39284 28366
rect 39228 27918 39230 27970
rect 39282 27918 39284 27970
rect 39228 27906 39284 27918
rect 39116 27748 39172 27758
rect 39452 27748 39508 28476
rect 39676 27858 39732 28700
rect 39900 28644 39956 29598
rect 40012 28868 40068 34638
rect 40124 32674 40180 32686
rect 40124 32622 40126 32674
rect 40178 32622 40180 32674
rect 40124 31890 40180 32622
rect 40124 31838 40126 31890
rect 40178 31838 40180 31890
rect 40124 31826 40180 31838
rect 40236 30212 40292 37772
rect 40348 37716 40404 40684
rect 40460 39732 40516 42702
rect 40460 39666 40516 39676
rect 41020 40066 41076 42812
rect 41244 42868 41300 42878
rect 41244 42754 41300 42812
rect 41244 42702 41246 42754
rect 41298 42702 41300 42754
rect 41244 41972 41300 42702
rect 41244 41906 41300 41916
rect 41692 41972 41748 41982
rect 41804 41972 41860 43484
rect 42028 42980 42084 44606
rect 42140 43986 42196 45388
rect 42140 43934 42142 43986
rect 42194 43934 42196 43986
rect 42140 43922 42196 43934
rect 42588 45332 42644 45342
rect 42588 43986 42644 45276
rect 42812 44772 42868 45838
rect 43372 45556 43428 46620
rect 43708 46228 43764 46956
rect 43820 47796 43876 47806
rect 44156 47796 44212 47806
rect 43820 47794 44212 47796
rect 43820 47742 43822 47794
rect 43874 47742 44158 47794
rect 44210 47742 44212 47794
rect 43820 47740 44212 47742
rect 43820 46788 43876 47740
rect 44156 47730 44212 47740
rect 45164 47794 45220 47806
rect 45164 47742 45166 47794
rect 45218 47742 45220 47794
rect 43820 46722 43876 46732
rect 45164 46900 45220 47742
rect 50204 47794 50260 47806
rect 50652 47796 50708 47806
rect 50204 47742 50206 47794
rect 50258 47742 50260 47794
rect 45500 46900 45556 46910
rect 45164 46898 45556 46900
rect 45164 46846 45502 46898
rect 45554 46846 45556 46898
rect 45164 46844 45556 46846
rect 44044 46676 44100 46686
rect 44044 46582 44100 46620
rect 44940 46674 44996 46686
rect 44940 46622 44942 46674
rect 44994 46622 44996 46674
rect 43708 46162 43764 46172
rect 43932 46562 43988 46574
rect 43932 46510 43934 46562
rect 43986 46510 43988 46562
rect 43932 46116 43988 46510
rect 43932 45892 43988 46060
rect 43260 44772 43316 44782
rect 42812 44770 43316 44772
rect 42812 44718 43262 44770
rect 43314 44718 43316 44770
rect 42812 44716 43316 44718
rect 42588 43934 42590 43986
rect 42642 43934 42644 43986
rect 42588 43922 42644 43934
rect 42700 44100 42756 44110
rect 42476 42980 42532 42990
rect 42028 42978 42532 42980
rect 42028 42926 42478 42978
rect 42530 42926 42532 42978
rect 42028 42924 42532 42926
rect 42476 42914 42532 42924
rect 42588 42868 42644 42878
rect 42588 42774 42644 42812
rect 42700 42866 42756 44044
rect 42812 43762 42868 43774
rect 42812 43710 42814 43762
rect 42866 43710 42868 43762
rect 42812 43092 42868 43710
rect 43260 43764 43316 44716
rect 42812 43026 42868 43036
rect 43036 43316 43092 43326
rect 42700 42814 42702 42866
rect 42754 42814 42756 42866
rect 41916 42644 41972 42654
rect 41916 42550 41972 42588
rect 42700 42644 42756 42814
rect 42700 42578 42756 42588
rect 42364 42532 42420 42542
rect 41916 41972 41972 41982
rect 41804 41970 41972 41972
rect 41804 41918 41918 41970
rect 41970 41918 41972 41970
rect 41804 41916 41972 41918
rect 41356 41748 41412 41758
rect 41356 40740 41412 41692
rect 41468 41524 41524 41534
rect 41468 41430 41524 41468
rect 41692 41076 41748 41916
rect 41916 41906 41972 41916
rect 42364 41970 42420 42476
rect 42364 41918 42366 41970
rect 42418 41918 42420 41970
rect 42364 41906 42420 41918
rect 43036 41970 43092 43260
rect 43260 42868 43316 43708
rect 43260 42802 43316 42812
rect 43036 41918 43038 41970
rect 43090 41918 43092 41970
rect 43036 41906 43092 41918
rect 43148 42644 43204 42654
rect 42140 41858 42196 41870
rect 42140 41806 42142 41858
rect 42194 41806 42196 41858
rect 42140 41748 42196 41806
rect 42140 41682 42196 41692
rect 42700 41186 42756 41198
rect 42700 41134 42702 41186
rect 42754 41134 42756 41186
rect 41692 41020 41972 41076
rect 41356 40674 41412 40684
rect 41916 40962 41972 41020
rect 41916 40910 41918 40962
rect 41970 40910 41972 40962
rect 41020 40014 41022 40066
rect 41074 40014 41076 40066
rect 41020 39844 41076 40014
rect 41916 40068 41972 40910
rect 42700 40626 42756 41134
rect 43148 40964 43204 42588
rect 43372 41858 43428 45500
rect 43708 45890 43988 45892
rect 43708 45838 43934 45890
rect 43986 45838 43988 45890
rect 43708 45836 43988 45838
rect 43708 44884 43764 45836
rect 43932 45826 43988 45836
rect 44044 46228 44100 46238
rect 44044 46002 44100 46172
rect 44044 45950 44046 46002
rect 44098 45950 44100 46002
rect 43708 44790 43764 44828
rect 43820 45666 43876 45678
rect 43820 45614 43822 45666
rect 43874 45614 43876 45666
rect 43484 44770 43540 44782
rect 43484 44718 43486 44770
rect 43538 44718 43540 44770
rect 43484 44324 43540 44718
rect 43484 44258 43540 44268
rect 43596 44658 43652 44670
rect 43596 44606 43598 44658
rect 43650 44606 43652 44658
rect 43484 44100 43540 44110
rect 43484 44006 43540 44044
rect 43596 43204 43652 44606
rect 43596 43138 43652 43148
rect 43596 42868 43652 42878
rect 43596 42774 43652 42812
rect 43708 41972 43764 41982
rect 43820 41972 43876 45614
rect 44044 45108 44100 45950
rect 44940 46004 44996 46622
rect 45164 46228 45220 46844
rect 45500 46834 45556 46844
rect 45164 46162 45220 46172
rect 46172 46116 46228 46126
rect 46172 46022 46228 46060
rect 44940 45948 45332 46004
rect 45276 45917 45332 45948
rect 45276 45865 45278 45917
rect 45330 45865 45332 45917
rect 43932 45052 44212 45108
rect 43932 44770 43988 45052
rect 43932 44718 43934 44770
rect 43986 44718 43988 44770
rect 43932 44706 43988 44718
rect 44044 44884 44100 44894
rect 43932 44324 43988 44334
rect 43932 43652 43988 44268
rect 44044 43874 44100 44828
rect 44156 44772 44212 45052
rect 44716 44884 44772 44894
rect 44830 44884 44886 44894
rect 45276 44884 45332 45865
rect 48076 45892 48132 45902
rect 48748 45892 48804 45902
rect 44772 44882 44886 44884
rect 44772 44830 44832 44882
rect 44884 44830 44886 44882
rect 44772 44828 44886 44830
rect 44716 44818 44772 44828
rect 44830 44818 44886 44828
rect 45164 44882 45332 44884
rect 45164 44830 45278 44882
rect 45330 44830 45332 44882
rect 45164 44828 45332 44830
rect 44156 44100 44212 44716
rect 45052 44772 45108 44782
rect 45052 44678 45108 44716
rect 44156 44034 44212 44044
rect 44940 44658 44996 44670
rect 44940 44606 44942 44658
rect 44994 44606 44996 44658
rect 44044 43822 44046 43874
rect 44098 43822 44100 43874
rect 44044 43810 44100 43822
rect 43932 42866 43988 43596
rect 44940 43316 44996 44606
rect 45164 43874 45220 44828
rect 45276 44818 45332 44828
rect 46620 45780 46676 45790
rect 47068 45780 47124 45790
rect 46620 45778 47124 45780
rect 46620 45726 46622 45778
rect 46674 45726 47070 45778
rect 47122 45726 47124 45778
rect 46620 45724 47124 45726
rect 46620 44882 46676 45724
rect 46620 44830 46622 44882
rect 46674 44830 46676 44882
rect 46620 44772 46676 44830
rect 46620 44706 46676 44716
rect 45164 43822 45166 43874
rect 45218 43822 45220 43874
rect 45164 43652 45220 43822
rect 45164 43586 45220 43596
rect 45948 44098 46004 44110
rect 45948 44046 45950 44098
rect 46002 44046 46004 44098
rect 44940 43250 44996 43260
rect 45164 43204 45220 43214
rect 45220 43148 45332 43204
rect 45164 43138 45220 43148
rect 43932 42814 43934 42866
rect 43986 42814 43988 42866
rect 43932 42802 43988 42814
rect 45164 42756 45220 42766
rect 44044 42754 45220 42756
rect 44044 42702 45166 42754
rect 45218 42702 45220 42754
rect 44044 42700 45220 42702
rect 44044 42082 44100 42700
rect 45164 42690 45220 42700
rect 44716 42532 44772 42542
rect 44716 42438 44772 42476
rect 44044 42030 44046 42082
rect 44098 42030 44100 42082
rect 44044 42018 44100 42030
rect 43708 41970 43876 41972
rect 43708 41918 43710 41970
rect 43762 41918 43876 41970
rect 43708 41916 43876 41918
rect 45164 41972 45220 41982
rect 45276 41972 45332 43148
rect 45388 43092 45444 43102
rect 45388 42868 45444 43036
rect 45388 42866 45556 42868
rect 45388 42814 45390 42866
rect 45442 42814 45556 42866
rect 45388 42812 45556 42814
rect 45388 42802 45444 42812
rect 45164 41970 45332 41972
rect 45164 41918 45166 41970
rect 45218 41918 45332 41970
rect 45164 41916 45332 41918
rect 43708 41906 43764 41916
rect 45164 41906 45220 41916
rect 43372 41806 43374 41858
rect 43426 41806 43428 41858
rect 43372 41186 43428 41806
rect 44604 41860 44660 41870
rect 44604 41766 44660 41804
rect 43372 41134 43374 41186
rect 43426 41134 43428 41186
rect 43372 41122 43428 41134
rect 43596 40964 43652 40974
rect 43148 40962 43652 40964
rect 43148 40910 43150 40962
rect 43202 40910 43598 40962
rect 43650 40910 43652 40962
rect 43148 40908 43652 40910
rect 43148 40898 43204 40908
rect 42700 40574 42702 40626
rect 42754 40574 42756 40626
rect 41916 40002 41972 40012
rect 42028 40516 42084 40526
rect 41020 39618 41076 39788
rect 41468 39844 41524 39854
rect 41916 39844 41972 39854
rect 42028 39844 42084 40460
rect 41468 39750 41524 39788
rect 41580 39842 42084 39844
rect 41580 39790 41918 39842
rect 41970 39790 42084 39842
rect 41580 39788 42084 39790
rect 42140 39844 42196 39854
rect 41020 39566 41022 39618
rect 41074 39566 41076 39618
rect 41020 39554 41076 39566
rect 41580 39508 41636 39788
rect 41916 39778 41972 39788
rect 41356 39452 41636 39508
rect 41804 39618 41860 39630
rect 41804 39566 41806 39618
rect 41858 39566 41860 39618
rect 40572 38948 40628 38958
rect 40460 38722 40516 38734
rect 40460 38670 40462 38722
rect 40514 38670 40516 38722
rect 40460 37940 40516 38670
rect 40460 37874 40516 37884
rect 40348 37660 40516 37716
rect 40348 35812 40404 35822
rect 40348 35718 40404 35756
rect 40348 34020 40404 34030
rect 40348 33926 40404 33964
rect 40460 33460 40516 37660
rect 40348 33404 40516 33460
rect 40572 36706 40628 38892
rect 40796 38836 40852 38846
rect 40796 38722 40852 38780
rect 40796 38670 40798 38722
rect 40850 38670 40852 38722
rect 40796 38658 40852 38670
rect 41132 38724 41188 38762
rect 41132 38658 41188 38668
rect 41356 37828 41412 39452
rect 41244 37826 41412 37828
rect 41244 37774 41358 37826
rect 41410 37774 41412 37826
rect 41244 37772 41412 37774
rect 41244 37044 41300 37772
rect 41356 37762 41412 37772
rect 41468 38610 41524 38622
rect 41468 38558 41470 38610
rect 41522 38558 41524 38610
rect 41244 36978 41300 36988
rect 41356 37604 41412 37614
rect 40572 36654 40574 36706
rect 40626 36654 40628 36706
rect 40348 31948 40404 33404
rect 40572 32676 40628 36654
rect 41244 36708 41300 36718
rect 41244 36614 41300 36652
rect 41244 35812 41300 35822
rect 41244 35718 41300 35756
rect 40908 35586 40964 35598
rect 40908 35534 40910 35586
rect 40962 35534 40964 35586
rect 40908 35476 40964 35534
rect 41356 35476 41412 37548
rect 41468 36484 41524 38558
rect 41580 38052 41636 38062
rect 41580 37826 41636 37996
rect 41580 37774 41582 37826
rect 41634 37774 41636 37826
rect 41580 37762 41636 37774
rect 41804 37826 41860 39566
rect 42140 39620 42196 39788
rect 41916 38948 41972 38958
rect 41916 38836 41972 38892
rect 42028 38836 42084 38846
rect 41916 38834 42084 38836
rect 41916 38782 42030 38834
rect 42082 38782 42084 38834
rect 41916 38780 42084 38782
rect 42028 38770 42084 38780
rect 42028 37940 42084 37950
rect 42140 37940 42196 39564
rect 42476 39732 42532 39742
rect 42028 37938 42196 37940
rect 42028 37886 42030 37938
rect 42082 37886 42196 37938
rect 42028 37884 42196 37886
rect 42364 38948 42420 38958
rect 42028 37874 42084 37884
rect 41804 37774 41806 37826
rect 41858 37774 41860 37826
rect 41468 36418 41524 36428
rect 41692 35700 41748 35710
rect 41692 35606 41748 35644
rect 40908 35420 41524 35476
rect 40684 34578 40740 34590
rect 40684 34526 40686 34578
rect 40738 34526 40740 34578
rect 40684 33684 40740 34526
rect 41356 34578 41412 34590
rect 41356 34526 41358 34578
rect 41410 34526 41412 34578
rect 41020 33908 41076 33918
rect 41020 33684 41076 33852
rect 40684 33682 41076 33684
rect 40684 33630 41022 33682
rect 41074 33630 41076 33682
rect 40684 33628 41076 33630
rect 40572 32610 40628 32620
rect 40460 32564 40516 32574
rect 40460 32470 40516 32508
rect 40908 31948 40964 33628
rect 41020 33618 41076 33628
rect 41356 33684 41412 34526
rect 41356 33618 41412 33628
rect 41020 32676 41076 32686
rect 41020 32582 41076 32620
rect 40348 31892 40628 31948
rect 40908 31892 41076 31948
rect 41244 31892 41300 31902
rect 40572 30772 40628 31892
rect 40908 31668 40964 31678
rect 41020 31668 41076 31892
rect 41132 31836 41244 31892
rect 41132 31778 41188 31836
rect 41244 31826 41300 31836
rect 41132 31726 41134 31778
rect 41186 31726 41188 31778
rect 41132 31714 41188 31726
rect 41356 31778 41412 31790
rect 41356 31726 41358 31778
rect 41410 31726 41412 31778
rect 40964 31612 41076 31668
rect 40908 31602 40964 31612
rect 41020 31556 41076 31612
rect 41356 31556 41412 31726
rect 41020 31500 41412 31556
rect 40572 30706 40628 30716
rect 41132 30772 41188 30782
rect 40796 30660 40852 30670
rect 40796 30658 40964 30660
rect 40796 30606 40798 30658
rect 40850 30606 40964 30658
rect 40796 30604 40964 30606
rect 40796 30594 40852 30604
rect 40236 30146 40292 30156
rect 40460 30546 40516 30558
rect 40460 30494 40462 30546
rect 40514 30494 40516 30546
rect 40460 30098 40516 30494
rect 40460 30046 40462 30098
rect 40514 30046 40516 30098
rect 40460 30034 40516 30046
rect 40908 29876 40964 30604
rect 41132 30546 41188 30716
rect 41132 30494 41134 30546
rect 41186 30494 41188 30546
rect 41132 30482 41188 30494
rect 41244 29988 41300 29998
rect 40908 29782 40964 29820
rect 41132 29986 41300 29988
rect 41132 29934 41246 29986
rect 41298 29934 41300 29986
rect 41132 29932 41300 29934
rect 40348 29652 40404 29662
rect 40348 29558 40404 29596
rect 41132 29540 41188 29932
rect 41244 29922 41300 29932
rect 41468 29652 41524 35420
rect 41804 35252 41860 37774
rect 42364 37826 42420 38892
rect 42364 37774 42366 37826
rect 42418 37774 42420 37826
rect 41916 37602 41972 37614
rect 41916 37550 41918 37602
rect 41970 37550 41972 37602
rect 41916 36706 41972 37550
rect 41916 36654 41918 36706
rect 41970 36654 41972 36706
rect 41916 36642 41972 36654
rect 42364 35700 42420 37774
rect 42364 35634 42420 35644
rect 42476 37828 42532 39676
rect 42588 38724 42644 38762
rect 42588 38658 42644 38668
rect 42588 37828 42644 37838
rect 42476 37826 42644 37828
rect 42476 37774 42590 37826
rect 42642 37774 42644 37826
rect 42476 37772 42644 37774
rect 41804 35186 41860 35196
rect 41804 34580 41860 34590
rect 41804 34486 41860 34524
rect 42252 34578 42308 34590
rect 42252 34526 42254 34578
rect 42306 34526 42308 34578
rect 42140 34018 42196 34030
rect 42140 33966 42142 34018
rect 42194 33966 42196 34018
rect 41580 32676 41636 32686
rect 42140 32676 42196 33966
rect 42252 33908 42308 34526
rect 42252 33794 42308 33852
rect 42252 33742 42254 33794
rect 42306 33742 42308 33794
rect 42252 33730 42308 33742
rect 42364 33906 42420 33918
rect 42364 33854 42366 33906
rect 42418 33854 42420 33906
rect 42364 33796 42420 33854
rect 42364 33730 42420 33740
rect 42252 32676 42308 32686
rect 41580 32674 41748 32676
rect 41580 32622 41582 32674
rect 41634 32622 41748 32674
rect 41580 32620 41748 32622
rect 42140 32674 42308 32676
rect 42140 32622 42254 32674
rect 42306 32622 42308 32674
rect 42140 32620 42308 32622
rect 41580 32610 41636 32620
rect 41692 32114 41748 32620
rect 42252 32610 42308 32620
rect 41692 32062 41694 32114
rect 41746 32062 41748 32114
rect 41692 32050 41748 32062
rect 42028 32564 42084 32574
rect 42476 32564 42532 37772
rect 42588 37762 42644 37772
rect 42700 37604 42756 40574
rect 43596 40516 43652 40908
rect 43596 40180 43652 40460
rect 45388 40626 45444 40638
rect 45388 40574 45390 40626
rect 45442 40574 45444 40626
rect 43596 40114 43652 40124
rect 43932 40292 43988 40302
rect 45388 40292 45444 40574
rect 43260 38722 43316 38734
rect 43260 38670 43262 38722
rect 43314 38670 43316 38722
rect 43260 38668 43316 38670
rect 43260 38612 43428 38668
rect 42700 37538 42756 37548
rect 43036 38052 43092 38062
rect 42588 36932 42644 36942
rect 42588 36820 42644 36876
rect 43036 36932 43092 37996
rect 43260 37940 43316 37950
rect 43260 37846 43316 37884
rect 43148 36932 43204 36942
rect 43036 36930 43204 36932
rect 43036 36878 43150 36930
rect 43202 36878 43204 36930
rect 43036 36876 43204 36878
rect 42700 36820 42756 36830
rect 42588 36818 42756 36820
rect 42588 36766 42702 36818
rect 42754 36766 42756 36818
rect 42588 36764 42756 36766
rect 42700 36484 42756 36764
rect 42700 36482 42868 36484
rect 42700 36430 42702 36482
rect 42754 36430 42868 36482
rect 42700 36428 42868 36430
rect 42700 36418 42756 36428
rect 42700 35812 42756 35822
rect 42700 34692 42756 35756
rect 42812 35810 42868 36428
rect 43036 35922 43092 36876
rect 43148 36866 43204 36876
rect 43036 35870 43038 35922
rect 43090 35870 43092 35922
rect 43036 35858 43092 35870
rect 42812 35758 42814 35810
rect 42866 35758 42868 35810
rect 42812 35746 42868 35758
rect 43372 35586 43428 38612
rect 43932 37042 43988 40236
rect 45276 40236 45444 40292
rect 45500 40292 45556 42812
rect 45612 42756 45668 42766
rect 45612 42662 45668 42700
rect 45836 41972 45892 41982
rect 45948 41972 46004 44046
rect 46956 43874 47012 45724
rect 47068 45714 47124 45724
rect 48076 44098 48132 45836
rect 48636 45890 48804 45892
rect 48636 45838 48750 45890
rect 48802 45838 48804 45890
rect 48636 45836 48804 45838
rect 48076 44046 48078 44098
rect 48130 44046 48132 44098
rect 48076 44034 48132 44046
rect 48188 45778 48244 45790
rect 48188 45726 48190 45778
rect 48242 45726 48244 45778
rect 46956 43822 46958 43874
rect 47010 43822 47012 43874
rect 46956 43810 47012 43822
rect 47292 43874 47348 43886
rect 47292 43822 47294 43874
rect 47346 43822 47348 43874
rect 47292 43202 47348 43822
rect 47292 43150 47294 43202
rect 47346 43150 47348 43202
rect 47292 42978 47348 43150
rect 47292 42926 47294 42978
rect 47346 42926 47348 42978
rect 47292 42914 47348 42926
rect 47404 43874 47460 43886
rect 47404 43822 47406 43874
rect 47458 43822 47460 43874
rect 47404 43652 47460 43822
rect 46396 42868 46452 42878
rect 46396 42774 46452 42812
rect 46844 42644 46900 42654
rect 46844 42550 46900 42588
rect 47404 42644 47460 43596
rect 47628 43874 47684 43886
rect 47628 43822 47630 43874
rect 47682 43822 47684 43874
rect 47628 42868 47684 43822
rect 47740 43090 47796 43102
rect 47740 43038 47742 43090
rect 47794 43038 47796 43090
rect 47740 42978 47796 43038
rect 47740 42926 47742 42978
rect 47794 42926 47796 42978
rect 47740 42914 47796 42926
rect 47628 42802 47684 42812
rect 47404 42578 47460 42588
rect 48188 42644 48244 45726
rect 48524 45220 48580 45230
rect 48636 45220 48692 45836
rect 48748 45826 48804 45836
rect 49084 45890 49140 45902
rect 49084 45838 49086 45890
rect 49138 45838 49140 45890
rect 49084 45332 49140 45838
rect 49420 45892 49476 45902
rect 49420 45798 49476 45836
rect 49756 45890 49812 45902
rect 49756 45838 49758 45890
rect 49810 45838 49812 45890
rect 49756 45444 49812 45838
rect 49756 45378 49812 45388
rect 50092 45444 50148 45454
rect 49084 45266 49140 45276
rect 48524 45218 48692 45220
rect 48524 45166 48526 45218
rect 48578 45166 48692 45218
rect 48524 45164 48692 45166
rect 48524 45154 48580 45164
rect 49644 44660 49700 44670
rect 49644 43988 49700 44604
rect 49084 43986 49700 43988
rect 49084 43934 49646 43986
rect 49698 43934 49700 43986
rect 49084 43932 49700 43934
rect 48636 43764 48692 43774
rect 48636 43202 48692 43708
rect 48636 43150 48638 43202
rect 48690 43150 48692 43202
rect 48636 42978 48692 43150
rect 48636 42926 48638 42978
rect 48690 42926 48692 42978
rect 48636 42914 48692 42926
rect 49084 43090 49140 43932
rect 49644 43922 49700 43932
rect 49532 43764 49588 43774
rect 49532 43670 49588 43708
rect 49084 43038 49086 43090
rect 49138 43038 49140 43090
rect 49084 42978 49140 43038
rect 49084 42926 49086 42978
rect 49138 42926 49140 42978
rect 48188 42550 48244 42588
rect 48972 42084 49028 42094
rect 49084 42084 49140 42926
rect 49756 42868 49812 42878
rect 48972 42082 49084 42084
rect 48972 42030 48974 42082
rect 49026 42030 49084 42082
rect 48972 42028 49084 42030
rect 48972 42018 49028 42028
rect 49084 42018 49140 42028
rect 49420 42644 49476 42654
rect 45836 41970 46004 41972
rect 45836 41918 45838 41970
rect 45890 41918 46004 41970
rect 45836 41916 46004 41918
rect 45836 41906 45892 41916
rect 46620 41860 46676 41870
rect 46620 41766 46676 41804
rect 49420 41746 49476 42588
rect 49420 41694 49422 41746
rect 49474 41694 49476 41746
rect 49420 41634 49476 41694
rect 49420 41582 49422 41634
rect 49474 41582 49476 41634
rect 49420 41570 49476 41582
rect 49756 42642 49812 42812
rect 49756 42590 49758 42642
rect 49810 42590 49812 42642
rect 47964 40852 48020 40862
rect 49420 40852 49476 40862
rect 47964 40758 48020 40796
rect 49308 40796 49420 40852
rect 47068 40740 47124 40750
rect 47068 40646 47124 40684
rect 47740 40740 47796 40750
rect 47740 40646 47796 40684
rect 48300 40738 48356 40750
rect 48300 40686 48302 40738
rect 48354 40686 48356 40738
rect 44940 40180 44996 40190
rect 44492 40068 44548 40078
rect 44268 40012 44492 40068
rect 44044 39732 44100 39742
rect 44044 39638 44100 39676
rect 44268 38946 44324 40012
rect 44492 39974 44548 40012
rect 44940 40066 44996 40124
rect 44940 40014 44942 40066
rect 44994 40014 44996 40066
rect 44940 40002 44996 40014
rect 45276 40180 45332 40236
rect 45500 40226 45556 40236
rect 47292 40514 47348 40526
rect 47292 40462 47294 40514
rect 47346 40462 47348 40514
rect 44268 38894 44270 38946
rect 44322 38894 44324 38946
rect 44268 38882 44324 38894
rect 44604 38836 44660 38846
rect 45276 38836 45332 40124
rect 46396 40180 46452 40190
rect 45388 40068 45444 40078
rect 45444 40012 45780 40068
rect 45388 39974 45444 40012
rect 45724 39954 45780 40012
rect 45724 39902 45726 39954
rect 45778 39902 45780 39954
rect 45724 39890 45780 39902
rect 46396 40066 46452 40124
rect 46396 40014 46398 40066
rect 46450 40014 46452 40066
rect 45388 38836 45444 38846
rect 45276 38834 45444 38836
rect 45276 38782 45390 38834
rect 45442 38782 45444 38834
rect 45276 38780 45444 38782
rect 44604 37938 44660 38780
rect 45388 38770 45444 38780
rect 44940 38724 44996 38762
rect 44940 38658 44996 38668
rect 46396 38052 46452 40014
rect 44604 37886 44606 37938
rect 44658 37886 44660 37938
rect 44604 37874 44660 37886
rect 46284 37996 46396 38052
rect 46284 37828 46340 37996
rect 46396 37986 46452 37996
rect 46508 40068 46564 40078
rect 46508 38724 46564 40012
rect 46508 37938 46564 38668
rect 46508 37886 46510 37938
rect 46562 37886 46564 37938
rect 46508 37874 46564 37886
rect 46732 39732 46788 39742
rect 46732 38722 46788 39676
rect 46732 38670 46734 38722
rect 46786 38670 46788 38722
rect 43932 36990 43934 37042
rect 43986 36990 43988 37042
rect 43932 36978 43988 36990
rect 45948 37826 46340 37828
rect 45948 37774 46286 37826
rect 46338 37774 46340 37826
rect 45948 37772 46340 37774
rect 45948 36818 46004 37772
rect 46284 37762 46340 37772
rect 45948 36766 45950 36818
rect 46002 36766 46004 36818
rect 45948 36754 46004 36766
rect 44268 36708 44324 36718
rect 44156 36706 44324 36708
rect 44156 36654 44270 36706
rect 44322 36654 44324 36706
rect 44156 36652 44324 36654
rect 43596 36594 43652 36606
rect 43596 36542 43598 36594
rect 43650 36542 43652 36594
rect 43596 36482 43652 36542
rect 43596 36430 43598 36482
rect 43650 36430 43652 36482
rect 43596 36418 43652 36430
rect 43372 35534 43374 35586
rect 43426 35534 43428 35586
rect 43372 35522 43428 35534
rect 44044 35810 44100 35822
rect 44044 35758 44046 35810
rect 44098 35758 44100 35810
rect 43708 35364 43764 35374
rect 42812 34692 42868 34702
rect 42700 34690 42868 34692
rect 42700 34638 42814 34690
rect 42866 34638 42868 34690
rect 42700 34636 42868 34638
rect 42812 34626 42868 34636
rect 42924 34580 42980 34590
rect 42588 32564 42644 32574
rect 42476 32508 42588 32564
rect 41692 30098 41748 30110
rect 41692 30046 41694 30098
rect 41746 30046 41748 30098
rect 41692 29986 41748 30046
rect 41692 29934 41694 29986
rect 41746 29934 41748 29986
rect 41692 29922 41748 29934
rect 41132 28868 41188 29484
rect 40012 28812 40292 28868
rect 40236 28754 40292 28812
rect 41132 28802 41188 28812
rect 41244 29596 41524 29652
rect 41244 29090 41300 29596
rect 41244 29038 41246 29090
rect 41298 29038 41300 29090
rect 40236 28702 40238 28754
rect 40290 28702 40292 28754
rect 39900 28588 40068 28644
rect 39676 27806 39678 27858
rect 39730 27806 39732 27858
rect 39676 27794 39732 27806
rect 39900 28418 39956 28430
rect 39900 28366 39902 28418
rect 39954 28366 39956 28418
rect 39116 27746 39508 27748
rect 39116 27694 39118 27746
rect 39170 27694 39508 27746
rect 39116 27692 39508 27694
rect 39788 27748 39844 27758
rect 39116 27682 39172 27692
rect 39788 27654 39844 27692
rect 39004 27468 39284 27524
rect 38892 27244 39172 27300
rect 38780 26908 39060 26964
rect 38556 26740 38612 26908
rect 39004 26850 39060 26908
rect 39004 26798 39006 26850
rect 39058 26798 39060 26850
rect 39004 26786 39060 26798
rect 39116 26852 39172 27244
rect 39116 26786 39172 26796
rect 38332 26684 38612 26740
rect 38780 26740 38836 26750
rect 38332 26514 38388 26684
rect 38332 26462 38334 26514
rect 38386 26462 38388 26514
rect 38332 26404 38388 26462
rect 38332 26338 38388 26348
rect 38444 26516 38500 26526
rect 37996 26002 38052 26012
rect 37884 25956 37940 25966
rect 37772 25954 37940 25956
rect 37772 25902 37886 25954
rect 37938 25902 37940 25954
rect 37772 25900 37940 25902
rect 37548 25842 37604 25854
rect 37548 25790 37550 25842
rect 37602 25790 37604 25842
rect 37548 25396 37604 25790
rect 37548 25330 37604 25340
rect 37436 24334 37438 24386
rect 37490 24334 37492 24386
rect 37436 24322 37492 24334
rect 37548 24610 37604 24622
rect 37548 24558 37550 24610
rect 37602 24558 37604 24610
rect 36988 24050 37380 24052
rect 36988 23998 36990 24050
rect 37042 23998 37380 24050
rect 36988 23996 37380 23998
rect 36988 23986 37044 23996
rect 36764 23886 36766 23938
rect 36818 23886 36820 23938
rect 36764 23874 36820 23886
rect 37548 23940 37604 24558
rect 37772 24610 37828 25900
rect 37884 25890 37940 25900
rect 37772 24558 37774 24610
rect 37826 24558 37828 24610
rect 37660 23940 37716 23950
rect 37548 23938 37716 23940
rect 37548 23886 37662 23938
rect 37714 23886 37716 23938
rect 37548 23884 37716 23886
rect 37660 23874 37716 23884
rect 36540 23826 36708 23828
rect 36540 23774 36542 23826
rect 36594 23774 36708 23826
rect 36540 23772 36708 23774
rect 37100 23826 37156 23838
rect 37100 23774 37102 23826
rect 37154 23774 37156 23826
rect 36540 23762 36596 23772
rect 36204 23716 36260 23726
rect 35756 22866 35812 22876
rect 35868 23042 35924 23054
rect 35868 22990 35870 23042
rect 35922 22990 35924 23042
rect 35420 22706 35588 22708
rect 35420 22654 35422 22706
rect 35474 22654 35588 22706
rect 35420 22652 35588 22654
rect 35644 22706 35700 22718
rect 35644 22654 35646 22706
rect 35698 22654 35700 22706
rect 35084 22596 35140 22606
rect 33628 22430 33630 22482
rect 33682 22430 33684 22482
rect 33628 22418 33684 22430
rect 34524 22482 34580 22494
rect 34524 22430 34526 22482
rect 34578 22430 34580 22482
rect 33292 22204 33460 22260
rect 33180 21588 33236 21598
rect 33180 21494 33236 21532
rect 33068 20468 33124 20478
rect 32844 20466 33124 20468
rect 32844 20414 33070 20466
rect 33122 20414 33124 20466
rect 32844 20412 33124 20414
rect 33068 20402 33124 20412
rect 33180 20020 33236 20030
rect 33180 19572 33236 19964
rect 32508 18610 32564 18620
rect 33068 19570 33236 19572
rect 33068 19518 33182 19570
rect 33234 19518 33236 19570
rect 33068 19516 33236 19518
rect 32172 17836 32452 17892
rect 32060 16606 32062 16658
rect 32114 16606 32116 16658
rect 32060 16594 32116 16606
rect 32172 17668 32228 17678
rect 31948 16380 32116 16436
rect 32060 15652 32116 16380
rect 32172 15762 32228 17612
rect 32284 17554 32340 17566
rect 32284 17502 32286 17554
rect 32338 17502 32340 17554
rect 32284 16548 32340 17502
rect 32396 17556 32452 17836
rect 32508 17556 32564 17566
rect 32396 17500 32508 17556
rect 32508 17490 32564 17500
rect 32284 16482 32340 16492
rect 32172 15710 32174 15762
rect 32226 15710 32228 15762
rect 32172 15698 32228 15710
rect 31836 15596 32004 15652
rect 31948 15316 32004 15596
rect 31948 15250 32004 15260
rect 32060 13858 32116 15596
rect 32956 15652 33012 15662
rect 33068 15652 33124 19516
rect 33180 19506 33236 19516
rect 33292 19460 33348 22204
rect 33628 21924 33684 21934
rect 34524 21924 34580 22430
rect 34748 21924 34804 21934
rect 34524 21868 34748 21924
rect 33404 20578 33460 20590
rect 33404 20526 33406 20578
rect 33458 20526 33460 20578
rect 33404 19908 33460 20526
rect 33404 19842 33460 19852
rect 33516 19460 33572 19470
rect 33292 19458 33572 19460
rect 33292 19406 33518 19458
rect 33570 19406 33572 19458
rect 33292 19404 33572 19406
rect 33180 18786 33236 18798
rect 33180 18734 33182 18786
rect 33234 18734 33236 18786
rect 33180 17778 33236 18734
rect 33180 17726 33182 17778
rect 33234 17726 33236 17778
rect 33180 17714 33236 17726
rect 33180 15652 33236 15662
rect 33068 15650 33236 15652
rect 33068 15598 33182 15650
rect 33234 15598 33236 15650
rect 33068 15596 33236 15598
rect 32956 15558 33012 15596
rect 32396 15538 32452 15550
rect 32396 15486 32398 15538
rect 32450 15486 32452 15538
rect 32396 15316 32452 15486
rect 32396 14756 32452 15260
rect 33180 15540 33236 15596
rect 32396 14690 32452 14700
rect 32508 15092 32564 15102
rect 32060 13806 32062 13858
rect 32114 13806 32116 13858
rect 32060 13794 32116 13806
rect 32508 13858 32564 15036
rect 33180 14980 33236 15484
rect 33180 14914 33236 14924
rect 32508 13806 32510 13858
rect 32562 13806 32564 13858
rect 32508 13794 32564 13806
rect 33292 14756 33348 14766
rect 33292 13858 33348 14700
rect 33292 13806 33294 13858
rect 33346 13806 33348 13858
rect 33292 13794 33348 13806
rect 33404 12740 33460 19404
rect 33516 19394 33572 19404
rect 33628 18788 33684 21868
rect 34748 21810 34804 21868
rect 34748 21758 34750 21810
rect 34802 21758 34804 21810
rect 34748 21746 34804 21758
rect 35084 21700 35140 22540
rect 35420 21924 35476 22652
rect 35532 21924 35588 21934
rect 35308 21868 35532 21924
rect 35196 21700 35252 21710
rect 34860 21698 35252 21700
rect 34860 21646 35198 21698
rect 35250 21646 35252 21698
rect 34860 21644 35252 21646
rect 34860 21588 34916 21644
rect 35196 21634 35252 21644
rect 34636 20804 34692 20814
rect 34860 20804 34916 21532
rect 35308 21476 35364 21868
rect 35532 21858 35588 21868
rect 35644 21700 35700 22654
rect 35868 22706 35924 22990
rect 35868 22654 35870 22706
rect 35922 22654 35924 22706
rect 35868 21812 35924 22654
rect 36204 22706 36260 23660
rect 36316 23714 36372 23726
rect 36316 23662 36318 23714
rect 36370 23662 36372 23714
rect 36316 22820 36372 23662
rect 37100 23156 37156 23774
rect 37324 23826 37380 23838
rect 37324 23774 37326 23826
rect 37378 23774 37380 23826
rect 37324 23716 37380 23774
rect 37772 23716 37828 24558
rect 38332 25844 38388 25854
rect 38108 24498 38164 24510
rect 38108 24446 38110 24498
rect 38162 24446 38164 24498
rect 38108 24388 38164 24446
rect 38108 24322 38164 24332
rect 38332 23940 38388 25788
rect 38444 25730 38500 26460
rect 38668 25956 38724 25966
rect 38668 25842 38724 25900
rect 38780 25954 38836 26684
rect 38892 26738 38948 26750
rect 38892 26686 38894 26738
rect 38946 26686 38948 26738
rect 38892 26628 38948 26686
rect 38892 26572 39060 26628
rect 39004 26516 39060 26572
rect 39004 26450 39060 26460
rect 39116 26626 39172 26638
rect 39116 26574 39118 26626
rect 39170 26574 39172 26626
rect 38780 25902 38782 25954
rect 38834 25902 38836 25954
rect 38780 25890 38836 25902
rect 38892 26404 38948 26414
rect 38668 25790 38670 25842
rect 38722 25790 38724 25842
rect 38668 25778 38724 25790
rect 38444 25678 38446 25730
rect 38498 25678 38500 25730
rect 38444 25666 38500 25678
rect 38892 25730 38948 26348
rect 39116 26292 39172 26574
rect 39228 26516 39284 27468
rect 39340 26740 39396 26750
rect 39788 26740 39844 26750
rect 39340 26738 39844 26740
rect 39340 26686 39342 26738
rect 39394 26686 39790 26738
rect 39842 26686 39844 26738
rect 39340 26684 39844 26686
rect 39340 26674 39396 26684
rect 39788 26674 39844 26684
rect 39900 26740 39956 28366
rect 40012 27860 40068 28588
rect 40236 27860 40292 28702
rect 41244 28754 41300 29038
rect 41244 28702 41246 28754
rect 41298 28702 41300 28754
rect 41244 28690 41300 28702
rect 41692 28644 41748 28654
rect 41692 28530 41748 28588
rect 41692 28478 41694 28530
rect 41746 28478 41748 28530
rect 40908 28418 40964 28430
rect 40908 28366 40910 28418
rect 40962 28366 40964 28418
rect 40908 27972 40964 28366
rect 40684 27916 40964 27972
rect 41692 27972 41748 28478
rect 42028 28532 42084 32508
rect 42588 32498 42644 32508
rect 42924 32564 42980 34524
rect 43148 34580 43204 34590
rect 43148 34486 43204 34524
rect 43484 33796 43540 33806
rect 43484 32898 43540 33740
rect 43708 33684 43764 35308
rect 44044 35364 44100 35758
rect 44044 34916 44100 35308
rect 44156 35140 44212 36652
rect 44268 36642 44324 36652
rect 45164 36708 45220 36718
rect 45164 36614 45220 36652
rect 46732 36596 46788 38670
rect 46732 36530 46788 36540
rect 44380 35810 44436 35822
rect 44380 35758 44382 35810
rect 44434 35758 44436 35810
rect 44380 35252 44436 35758
rect 44492 35700 44548 35710
rect 44492 35606 44548 35644
rect 44940 35698 44996 35710
rect 44940 35646 44942 35698
rect 44994 35646 44996 35698
rect 44940 35364 44996 35646
rect 44940 35298 44996 35308
rect 45388 35698 45444 35710
rect 45388 35646 45390 35698
rect 45442 35646 45444 35698
rect 44380 35186 44436 35196
rect 44268 35140 44324 35150
rect 44156 35084 44268 35140
rect 44268 35074 44324 35084
rect 44828 35140 44884 35150
rect 44044 34822 44100 34860
rect 44716 34916 44772 34926
rect 44492 34692 44548 34702
rect 44380 34636 44492 34692
rect 44268 33796 44324 33806
rect 44268 33702 44324 33740
rect 43820 33684 43876 33694
rect 43764 33682 43876 33684
rect 43764 33630 43822 33682
rect 43874 33630 43876 33682
rect 43764 33628 43876 33630
rect 43708 33618 43764 33628
rect 43820 33618 43876 33628
rect 43484 32846 43486 32898
rect 43538 32846 43540 32898
rect 43036 32564 43092 32574
rect 42924 32562 43092 32564
rect 42924 32510 43038 32562
rect 43090 32510 43092 32562
rect 42924 32508 43092 32510
rect 42140 31892 42196 31902
rect 42140 30770 42196 31836
rect 42812 31890 42868 31902
rect 42812 31838 42814 31890
rect 42866 31838 42868 31890
rect 42140 30718 42142 30770
rect 42194 30718 42196 30770
rect 42140 30098 42196 30718
rect 42140 30046 42142 30098
rect 42194 30046 42196 30098
rect 42140 30034 42196 30046
rect 42364 30772 42420 30782
rect 42812 30772 42868 31838
rect 42924 31666 42980 32508
rect 43036 32498 43092 32508
rect 43484 31948 43540 32846
rect 43932 32898 43988 32910
rect 43932 32846 43934 32898
rect 43986 32846 43988 32898
rect 43932 32788 43988 32846
rect 43932 32722 43988 32732
rect 44268 32788 44324 32798
rect 44380 32788 44436 34636
rect 44492 34626 44548 34636
rect 44716 34020 44772 34860
rect 44716 33926 44772 33964
rect 44268 32786 44436 32788
rect 44268 32734 44270 32786
rect 44322 32734 44436 32786
rect 44268 32732 44436 32734
rect 44268 32722 44324 32732
rect 43036 31892 43540 31948
rect 44380 32002 44436 32014
rect 44380 31950 44382 32002
rect 44434 31950 44436 32002
rect 44380 31948 44436 31950
rect 44828 31948 44884 35084
rect 44940 34916 44996 34926
rect 44940 34822 44996 34860
rect 45388 34580 45444 35646
rect 45836 35364 45892 35374
rect 45388 34578 45556 34580
rect 45388 34526 45390 34578
rect 45442 34526 45556 34578
rect 45388 34524 45556 34526
rect 45388 34514 45444 34524
rect 45500 33796 45556 34524
rect 45836 34578 45892 35308
rect 45836 34526 45838 34578
rect 45890 34526 45892 34578
rect 45724 33796 45780 33806
rect 45500 33740 45724 33796
rect 45724 33702 45780 33740
rect 45164 33684 45220 33694
rect 45388 33684 45444 33694
rect 45220 33628 45332 33684
rect 45164 33618 45220 33628
rect 45276 33460 45332 33628
rect 45388 33682 45556 33684
rect 45388 33630 45390 33682
rect 45442 33630 45556 33682
rect 45388 33628 45556 33630
rect 45388 33618 45444 33628
rect 45276 33404 45444 33460
rect 45052 32898 45108 32910
rect 45052 32846 45054 32898
rect 45106 32846 45108 32898
rect 44380 31892 44548 31948
rect 44828 31892 44996 31948
rect 43036 31778 43092 31836
rect 43036 31726 43038 31778
rect 43090 31726 43092 31778
rect 43036 31714 43092 31726
rect 42924 31614 42926 31666
rect 42978 31614 42980 31666
rect 42924 30884 42980 31614
rect 44492 30884 44548 31892
rect 42924 30828 43428 30884
rect 44492 30828 44772 30884
rect 42364 30770 42868 30772
rect 42364 30718 42366 30770
rect 42418 30718 42868 30770
rect 42364 30716 42868 30718
rect 42140 29652 42196 29662
rect 42140 29650 42308 29652
rect 42140 29598 42142 29650
rect 42194 29598 42308 29650
rect 42140 29596 42308 29598
rect 42140 29586 42196 29596
rect 42252 29540 42308 29596
rect 42364 29540 42420 30716
rect 42588 30098 42644 30110
rect 42588 30046 42590 30098
rect 42642 30046 42644 30098
rect 42588 29988 42644 30046
rect 42588 29986 42868 29988
rect 42588 29934 42590 29986
rect 42642 29934 42868 29986
rect 42588 29932 42868 29934
rect 42588 29922 42644 29932
rect 42252 29484 42420 29540
rect 42140 29428 42196 29438
rect 42140 28868 42196 29372
rect 42140 28866 42308 28868
rect 42140 28814 42142 28866
rect 42194 28814 42308 28866
rect 42140 28812 42308 28814
rect 42140 28802 42196 28812
rect 42028 28466 42084 28476
rect 40236 27804 40516 27860
rect 40012 27766 40068 27804
rect 40236 27634 40292 27646
rect 40236 27582 40238 27634
rect 40290 27582 40292 27634
rect 39900 26674 39956 26684
rect 40012 26852 40068 26862
rect 39564 26516 39620 26526
rect 39228 26460 39508 26516
rect 39116 26236 39396 26292
rect 39116 25956 39172 26236
rect 39116 25890 39172 25900
rect 39228 26068 39284 26078
rect 38892 25678 38894 25730
rect 38946 25678 38948 25730
rect 38892 25666 38948 25678
rect 39116 25394 39172 25406
rect 39116 25342 39118 25394
rect 39170 25342 39172 25394
rect 39116 24722 39172 25342
rect 39116 24670 39118 24722
rect 39170 24670 39172 24722
rect 39116 24658 39172 24670
rect 39228 24722 39284 26012
rect 39228 24670 39230 24722
rect 39282 24670 39284 24722
rect 39228 24658 39284 24670
rect 38444 24610 38500 24622
rect 38444 24558 38446 24610
rect 38498 24558 38500 24610
rect 38444 24164 38500 24558
rect 39340 24610 39396 26236
rect 39340 24558 39342 24610
rect 39394 24558 39396 24610
rect 39340 24546 39396 24558
rect 39452 24500 39508 26460
rect 39620 26460 39732 26516
rect 39564 26450 39620 26460
rect 39564 25730 39620 25742
rect 39564 25678 39566 25730
rect 39618 25678 39620 25730
rect 39564 25172 39620 25678
rect 39564 25106 39620 25116
rect 39564 24724 39620 24734
rect 39676 24724 39732 26460
rect 40012 26180 40068 26796
rect 40236 26738 40292 27582
rect 40348 27636 40404 27646
rect 40348 27542 40404 27580
rect 40236 26686 40238 26738
rect 40290 26686 40292 26738
rect 40236 26674 40292 26686
rect 39900 26124 40068 26180
rect 40348 26628 40404 26638
rect 39564 24722 39844 24724
rect 39564 24670 39566 24722
rect 39618 24670 39844 24722
rect 39564 24668 39844 24670
rect 39564 24658 39620 24668
rect 39452 24444 39620 24500
rect 38444 24108 38724 24164
rect 38556 23940 38612 23950
rect 38332 23938 38612 23940
rect 38332 23886 38558 23938
rect 38610 23886 38612 23938
rect 38332 23884 38612 23886
rect 38556 23874 38612 23884
rect 38668 23828 38724 24108
rect 39228 24050 39284 24062
rect 39228 23998 39230 24050
rect 39282 23998 39284 24050
rect 38892 23828 38948 23838
rect 38668 23826 38948 23828
rect 38668 23774 38894 23826
rect 38946 23774 38948 23826
rect 38668 23772 38948 23774
rect 37324 23660 37828 23716
rect 37884 23716 37940 23726
rect 37884 23622 37940 23660
rect 38220 23714 38276 23726
rect 38220 23662 38222 23714
rect 38274 23662 38276 23714
rect 37100 23100 37940 23156
rect 36988 22932 37044 22942
rect 36988 22838 37044 22876
rect 37884 22930 37940 23100
rect 37884 22878 37886 22930
rect 37938 22878 37940 22930
rect 37884 22866 37940 22878
rect 37548 22820 37604 22830
rect 36316 22764 36596 22820
rect 36204 22654 36206 22706
rect 36258 22654 36260 22706
rect 36204 22642 36260 22654
rect 36092 22596 36148 22606
rect 36092 22502 36148 22540
rect 36316 22596 36372 22606
rect 36316 22594 36484 22596
rect 36316 22542 36318 22594
rect 36370 22542 36484 22594
rect 36316 22540 36484 22542
rect 36316 22530 36372 22540
rect 35980 21812 36036 21822
rect 35868 21810 36036 21812
rect 35868 21758 35982 21810
rect 36034 21758 36036 21810
rect 35868 21756 36036 21758
rect 34636 20802 34916 20804
rect 34636 20750 34638 20802
rect 34690 20750 34916 20802
rect 34636 20748 34916 20750
rect 35084 21420 35364 21476
rect 35532 21644 35644 21700
rect 35084 20802 35140 21420
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 20750 35086 20802
rect 35138 20750 35140 20802
rect 34636 20738 34692 20748
rect 34188 20466 34244 20478
rect 34188 20414 34190 20466
rect 34242 20414 34244 20466
rect 34188 20020 34244 20414
rect 34188 19954 34244 19964
rect 34524 19908 34580 19918
rect 34580 19852 34692 19908
rect 34524 19814 34580 19852
rect 33852 19796 33908 19806
rect 34188 19796 34244 19806
rect 33852 19794 34188 19796
rect 33852 19742 33854 19794
rect 33906 19742 34188 19794
rect 33852 19740 34188 19742
rect 33852 19730 33908 19740
rect 34188 19702 34244 19740
rect 33628 18722 33684 18732
rect 34524 18788 34580 18798
rect 34524 18694 34580 18732
rect 34076 18564 34132 18574
rect 34076 18470 34132 18508
rect 34636 17892 34692 19852
rect 34748 18564 34804 20748
rect 35084 20738 35140 20750
rect 35532 20802 35588 21644
rect 35644 21634 35700 21644
rect 35532 20750 35534 20802
rect 35586 20750 35588 20802
rect 35532 20738 35588 20750
rect 35980 20802 36036 21756
rect 36204 21700 36260 21710
rect 36204 21642 36260 21644
rect 36204 21590 36206 21642
rect 36258 21590 36260 21642
rect 36204 21578 36260 21590
rect 36428 21364 36484 22540
rect 36540 21924 36596 22764
rect 37324 22706 37380 22718
rect 37324 22654 37326 22706
rect 37378 22654 37380 22706
rect 36652 21924 36708 21934
rect 36540 21922 36708 21924
rect 36540 21870 36654 21922
rect 36706 21870 36708 21922
rect 36540 21868 36708 21870
rect 36652 21858 36708 21868
rect 35980 20750 35982 20802
rect 36034 20750 36036 20802
rect 35980 20188 36036 20750
rect 36316 21308 36484 21364
rect 37100 21700 37156 21710
rect 36316 20188 36372 21308
rect 36428 20692 36484 20702
rect 36428 20598 36484 20636
rect 35980 20132 36260 20188
rect 35868 20020 35924 20030
rect 35196 19180 35460 19190
rect 35252 19124 35300 19180
rect 35356 19124 35404 19180
rect 35196 19114 35460 19124
rect 35420 18898 35476 18910
rect 35420 18846 35422 18898
rect 35474 18846 35476 18898
rect 35420 18786 35476 18846
rect 35420 18734 35422 18786
rect 35474 18734 35476 18786
rect 35420 18722 35476 18734
rect 35868 18786 35924 19964
rect 35980 18898 36036 20132
rect 36204 20020 36260 20132
rect 36316 20122 36372 20132
rect 37100 20580 37156 21644
rect 36652 20020 36708 20030
rect 36204 19964 36652 20020
rect 36204 19794 36260 19806
rect 36204 19742 36206 19794
rect 36258 19742 36260 19794
rect 36092 19684 36148 19694
rect 36092 19590 36148 19628
rect 35980 18846 35982 18898
rect 36034 18846 36036 18898
rect 35980 18834 36036 18846
rect 35868 18734 35870 18786
rect 35922 18734 35924 18786
rect 35868 18722 35924 18734
rect 36204 18788 36260 19742
rect 36652 19682 36708 19964
rect 36652 19630 36654 19682
rect 36706 19630 36708 19682
rect 36652 19618 36708 19630
rect 37100 19684 37156 20524
rect 37324 20466 37380 22654
rect 37548 22706 37604 22764
rect 38220 22820 38276 23662
rect 38276 22764 38500 22820
rect 38220 22754 38276 22764
rect 37548 22654 37550 22706
rect 37602 22654 37604 22706
rect 37548 22642 37604 22654
rect 38108 22706 38164 22718
rect 38108 22654 38110 22706
rect 38162 22654 38164 22706
rect 37884 21812 37940 21822
rect 37884 21718 37940 21756
rect 37772 21362 37828 21374
rect 37772 21310 37774 21362
rect 37826 21310 37828 21362
rect 37772 20690 37828 21310
rect 37660 20634 37716 20646
rect 37660 20582 37662 20634
rect 37714 20582 37716 20634
rect 37660 20580 37716 20582
rect 37660 20514 37716 20524
rect 37772 20638 37774 20690
rect 37826 20638 37828 20690
rect 37324 20414 37326 20466
rect 37378 20414 37380 20466
rect 37324 20402 37380 20414
rect 37660 20132 37716 20142
rect 37660 19684 37716 20076
rect 37772 20020 37828 20638
rect 38108 20188 38164 22654
rect 38444 22706 38500 22764
rect 38444 22654 38446 22706
rect 38498 22654 38500 22706
rect 38444 22642 38500 22654
rect 38668 21924 38724 21934
rect 38892 21924 38948 23772
rect 39116 23490 39172 23502
rect 39116 23438 39118 23490
rect 39170 23438 39172 23490
rect 39116 22818 39172 23438
rect 39116 22766 39118 22818
rect 39170 22766 39172 22818
rect 39116 22754 39172 22766
rect 38668 21922 38948 21924
rect 38668 21870 38670 21922
rect 38722 21870 38948 21922
rect 38668 21868 38948 21870
rect 38668 21858 38724 21868
rect 38220 21812 38276 21822
rect 38220 20690 38276 21756
rect 38780 21698 38836 21710
rect 38780 21646 38782 21698
rect 38834 21646 38836 21698
rect 38332 21586 38388 21598
rect 38332 21534 38334 21586
rect 38386 21534 38388 21586
rect 38332 21362 38388 21534
rect 38332 21310 38334 21362
rect 38386 21310 38388 21362
rect 38332 21298 38388 21310
rect 38780 20916 38836 21646
rect 38780 20850 38836 20860
rect 39116 21026 39172 21038
rect 39116 20974 39118 21026
rect 39170 20974 39172 21026
rect 38220 20638 38222 20690
rect 38274 20638 38276 20690
rect 38220 20626 38276 20638
rect 38556 20692 38612 20702
rect 38556 20598 38612 20636
rect 39116 20690 39172 20974
rect 39116 20638 39118 20690
rect 39170 20638 39172 20690
rect 39116 20188 39172 20638
rect 38108 20132 38276 20188
rect 37772 19954 37828 19964
rect 38220 19906 38276 20132
rect 38780 20132 39172 20188
rect 39228 20578 39284 23998
rect 39340 23940 39396 23950
rect 39340 23846 39396 23884
rect 39452 22034 39508 22046
rect 39452 21982 39454 22034
rect 39506 21982 39508 22034
rect 39452 21922 39508 21982
rect 39452 21870 39454 21922
rect 39506 21870 39508 21922
rect 39452 21026 39508 21870
rect 39452 20974 39454 21026
rect 39506 20974 39508 21026
rect 39452 20962 39508 20974
rect 39228 20526 39230 20578
rect 39282 20526 39284 20578
rect 38220 19854 38222 19906
rect 38274 19854 38276 19906
rect 38220 19842 38276 19854
rect 38668 20020 38724 20030
rect 37772 19684 37828 19694
rect 37660 19682 37828 19684
rect 37660 19630 37774 19682
rect 37826 19630 37828 19682
rect 37660 19628 37828 19630
rect 36204 18722 36260 18732
rect 36652 18788 36708 18798
rect 34972 18676 35028 18686
rect 34972 18582 35028 18620
rect 36316 18564 36372 18574
rect 34748 18498 34804 18508
rect 36092 18508 36316 18564
rect 33516 17666 33572 17678
rect 33516 17614 33518 17666
rect 33570 17614 33572 17666
rect 33516 17556 33572 17614
rect 33516 17490 33572 17500
rect 33852 17666 33908 17678
rect 33852 17614 33854 17666
rect 33906 17614 33908 17666
rect 33740 15650 33796 15662
rect 33740 15598 33742 15650
rect 33794 15598 33796 15650
rect 33628 15428 33684 15438
rect 33628 13858 33684 15372
rect 33740 15092 33796 15598
rect 33740 14644 33796 15036
rect 33852 14978 33908 17614
rect 34188 17668 34244 17678
rect 34636 17668 34692 17836
rect 35980 17778 36036 17790
rect 35980 17726 35982 17778
rect 36034 17726 36036 17778
rect 34748 17668 34804 17678
rect 34636 17666 34804 17668
rect 34636 17614 34750 17666
rect 34802 17614 34804 17666
rect 34636 17612 34804 17614
rect 34188 17574 34244 17612
rect 34748 17332 34804 17612
rect 35308 17666 35364 17678
rect 35308 17614 35310 17666
rect 35362 17614 35364 17666
rect 35308 17332 35364 17614
rect 35644 17556 35700 17566
rect 35308 17276 35588 17332
rect 34748 17266 34804 17276
rect 35196 17164 35460 17174
rect 35252 17108 35300 17164
rect 35356 17108 35404 17164
rect 35196 17098 35460 17108
rect 35532 16882 35588 17276
rect 35532 16830 35534 16882
rect 35586 16830 35588 16882
rect 35532 16818 35588 16830
rect 34412 16546 34468 16558
rect 34412 16494 34414 16546
rect 34466 16494 34468 16546
rect 34188 15650 34244 15662
rect 34188 15598 34190 15650
rect 34242 15598 34244 15650
rect 34188 15428 34244 15598
rect 34412 15652 34468 16494
rect 34412 15586 34468 15596
rect 34188 15362 34244 15372
rect 35196 15148 35460 15158
rect 35252 15092 35300 15148
rect 35356 15092 35404 15148
rect 35196 15082 35460 15092
rect 33852 14926 33854 14978
rect 33906 14926 33908 14978
rect 33852 14914 33908 14926
rect 33740 14578 33796 14588
rect 35084 14644 35140 14654
rect 35084 14550 35140 14588
rect 35532 14420 35588 14430
rect 35532 14326 35588 14364
rect 33628 13806 33630 13858
rect 33682 13806 33684 13858
rect 33628 13794 33684 13806
rect 35644 13746 35700 17500
rect 35980 15876 36036 17726
rect 35980 15810 36036 15820
rect 35980 14756 36036 14766
rect 36092 14756 36148 18508
rect 36316 18470 36372 18508
rect 35980 14754 36148 14756
rect 35980 14702 35982 14754
rect 36034 14702 36148 14754
rect 35980 14700 36148 14702
rect 36316 15652 36372 15662
rect 35980 14690 36036 14700
rect 36316 13858 36372 15596
rect 36652 15650 36708 18732
rect 37100 18786 37156 19628
rect 37100 18734 37102 18786
rect 37154 18734 37156 18786
rect 37100 18722 37156 18734
rect 37772 18788 37828 19628
rect 37772 18722 37828 18732
rect 38668 18786 38724 19964
rect 38668 18734 38670 18786
rect 38722 18734 38724 18786
rect 38668 18564 38724 18734
rect 38668 18498 38724 18508
rect 38780 19794 38836 20132
rect 38780 19742 38782 19794
rect 38834 19742 38836 19794
rect 38780 18676 38836 19742
rect 39228 19684 39284 20526
rect 39564 20188 39620 24444
rect 39788 23938 39844 24668
rect 39788 23886 39790 23938
rect 39842 23886 39844 23938
rect 39788 23490 39844 23886
rect 39788 23438 39790 23490
rect 39842 23438 39844 23490
rect 39788 23426 39844 23438
rect 39900 22818 39956 26124
rect 40012 25956 40068 25966
rect 40012 23940 40068 25900
rect 40124 25842 40180 25854
rect 40124 25790 40126 25842
rect 40178 25790 40180 25842
rect 40124 24724 40180 25790
rect 40236 25620 40292 25630
rect 40348 25620 40404 26572
rect 40236 25618 40404 25620
rect 40236 25566 40238 25618
rect 40290 25566 40404 25618
rect 40236 25564 40404 25566
rect 40236 25554 40292 25564
rect 40124 24668 40292 24724
rect 40124 24500 40180 24510
rect 40124 24406 40180 24444
rect 40236 24276 40292 24668
rect 40236 24210 40292 24220
rect 40236 23940 40292 23950
rect 40012 23938 40292 23940
rect 40012 23886 40014 23938
rect 40066 23886 40238 23938
rect 40290 23886 40292 23938
rect 40012 23884 40292 23886
rect 40012 23846 40068 23884
rect 40236 23874 40292 23884
rect 39900 22766 39902 22818
rect 39954 22766 39956 22818
rect 39900 22034 39956 22766
rect 39900 21982 39902 22034
rect 39954 21982 39956 22034
rect 39900 21970 39956 21982
rect 40236 23490 40292 23502
rect 40236 23438 40238 23490
rect 40290 23438 40292 23490
rect 40236 21924 40292 23438
rect 40348 23492 40404 25564
rect 40460 25396 40516 27804
rect 40572 26740 40628 26750
rect 40572 26646 40628 26684
rect 40684 26628 40740 27916
rect 41692 27906 41748 27916
rect 42140 27972 42196 27982
rect 42140 27878 42196 27916
rect 41020 27860 41076 27870
rect 40908 27748 40964 27758
rect 41020 27748 41076 27804
rect 40908 27746 41076 27748
rect 40908 27694 40910 27746
rect 40962 27694 41076 27746
rect 40908 27692 41076 27694
rect 41356 27860 41412 27870
rect 40908 27682 40964 27692
rect 41356 27636 41412 27804
rect 41356 27570 41412 27580
rect 42028 27748 42084 27758
rect 42252 27748 42308 28812
rect 42364 28644 42420 29484
rect 42588 28644 42644 28654
rect 42364 28588 42588 28644
rect 42588 28550 42644 28588
rect 42084 27746 42308 27748
rect 42084 27694 42254 27746
rect 42306 27694 42308 27746
rect 42084 27692 42308 27694
rect 41020 27524 41076 27534
rect 40684 26562 40740 26572
rect 40796 27522 41076 27524
rect 40796 27470 41022 27522
rect 41074 27470 41076 27522
rect 40796 27468 41076 27470
rect 40796 26626 40852 27468
rect 41020 27458 41076 27468
rect 40796 26574 40798 26626
rect 40850 26574 40852 26626
rect 40796 26562 40852 26574
rect 41692 26626 41748 26638
rect 41692 26574 41694 26626
rect 41746 26574 41748 26626
rect 41244 26404 41300 26414
rect 41244 26310 41300 26348
rect 41468 25954 41524 25966
rect 41468 25902 41470 25954
rect 41522 25902 41524 25954
rect 41244 25730 41300 25742
rect 41244 25678 41246 25730
rect 41298 25678 41300 25730
rect 40460 25340 40740 25396
rect 40572 25172 40628 25182
rect 40572 24498 40628 25116
rect 40572 24446 40574 24498
rect 40626 24446 40628 24498
rect 40572 24434 40628 24446
rect 40348 23042 40404 23436
rect 40348 22990 40350 23042
rect 40402 22990 40404 23042
rect 40348 22978 40404 22990
rect 40460 24164 40516 24174
rect 40348 22820 40404 22830
rect 40460 22820 40516 24108
rect 40348 22818 40516 22820
rect 40348 22766 40350 22818
rect 40402 22766 40516 22818
rect 40348 22764 40516 22766
rect 40348 22754 40404 22764
rect 40236 21868 40404 21924
rect 39900 21812 39956 21822
rect 39900 21718 39956 21756
rect 40348 21810 40404 21868
rect 40348 21758 40350 21810
rect 40402 21758 40404 21810
rect 40348 21746 40404 21758
rect 40460 21812 40516 22764
rect 40460 21746 40516 21756
rect 40684 21588 40740 25340
rect 41244 24610 41300 25678
rect 41244 24558 41246 24610
rect 41298 24558 41300 24610
rect 40796 24500 40852 24510
rect 40796 22818 40852 24444
rect 41244 23940 41300 24558
rect 41468 24724 41524 25902
rect 41692 25618 41748 26574
rect 42028 25732 42084 27692
rect 42252 27682 42308 27692
rect 42364 27972 42420 27982
rect 42140 26738 42196 26750
rect 42140 26686 42142 26738
rect 42194 26686 42196 26738
rect 42140 26628 42196 26686
rect 42140 26562 42196 26572
rect 42252 26626 42308 26638
rect 42252 26574 42254 26626
rect 42306 26574 42308 26626
rect 42140 25956 42196 25966
rect 42140 25862 42196 25900
rect 42028 25638 42084 25676
rect 41692 25566 41694 25618
rect 41746 25566 41748 25618
rect 41692 25554 41748 25566
rect 41692 24724 41748 24734
rect 41468 24722 41748 24724
rect 41468 24670 41694 24722
rect 41746 24670 41748 24722
rect 41468 24668 41748 24670
rect 41468 24500 41524 24668
rect 41692 24658 41748 24668
rect 41468 24434 41524 24444
rect 42140 24500 42196 24510
rect 41692 24276 41748 24286
rect 41244 23874 41300 23884
rect 41580 24164 41636 24174
rect 41580 23714 41636 24108
rect 41580 23662 41582 23714
rect 41634 23662 41636 23714
rect 41580 23650 41636 23662
rect 41244 23042 41300 23054
rect 41244 22990 41246 23042
rect 41298 22990 41300 23042
rect 40796 22766 40798 22818
rect 40850 22766 40852 22818
rect 40796 22754 40852 22766
rect 41020 22820 41076 22830
rect 41020 22036 41076 22764
rect 41244 22818 41300 22990
rect 41692 22930 41748 24220
rect 41692 22878 41694 22930
rect 41746 22878 41748 22930
rect 41692 22866 41748 22878
rect 41916 23940 41972 23950
rect 41244 22766 41246 22818
rect 41298 22766 41300 22818
rect 41244 22754 41300 22766
rect 41916 22820 41972 23884
rect 42140 23714 42196 24444
rect 42252 23826 42308 26574
rect 42364 25842 42420 27916
rect 42812 27970 42868 29932
rect 43260 29652 43316 30828
rect 43372 30770 43428 30828
rect 43372 30718 43374 30770
rect 43426 30718 43428 30770
rect 43372 30706 43428 30718
rect 44380 30546 44436 30558
rect 44380 30494 44382 30546
rect 44434 30494 44436 30546
rect 44380 29876 44436 30494
rect 44380 29810 44436 29820
rect 44716 29874 44772 30828
rect 44940 30660 44996 31892
rect 45052 31890 45108 32846
rect 45052 31838 45054 31890
rect 45106 31838 45108 31890
rect 45052 31826 45108 31838
rect 45276 32788 45332 32798
rect 45276 31780 45332 32732
rect 45388 32786 45444 33404
rect 45388 32734 45390 32786
rect 45442 32734 45444 32786
rect 45388 32722 45444 32734
rect 45500 31948 45556 33628
rect 45836 33572 45892 34526
rect 46060 34916 46116 34926
rect 46060 33684 46116 34860
rect 47180 34916 47236 34926
rect 46284 34578 46340 34590
rect 46284 34526 46286 34578
rect 46338 34526 46340 34578
rect 46284 33796 46340 34526
rect 47180 34018 47236 34860
rect 47180 33966 47182 34018
rect 47234 33966 47236 34018
rect 47180 33954 47236 33966
rect 46620 33796 46676 33806
rect 45724 33516 45892 33572
rect 45948 33682 46116 33684
rect 45948 33630 46062 33682
rect 46114 33630 46116 33682
rect 45948 33628 46116 33630
rect 45724 32788 45780 33516
rect 45724 32694 45780 32732
rect 45836 32788 45892 32798
rect 45948 32788 46004 33628
rect 46060 33570 46116 33628
rect 46060 33518 46062 33570
rect 46114 33518 46116 33570
rect 46060 33506 46116 33518
rect 46172 33740 46620 33796
rect 45836 32786 46004 32788
rect 45836 32734 45838 32786
rect 45890 32734 46004 32786
rect 45836 32732 46004 32734
rect 45836 32722 45892 32732
rect 45500 31892 45780 31948
rect 45724 31890 45780 31892
rect 45724 31838 45726 31890
rect 45778 31838 45780 31890
rect 45724 31826 45780 31838
rect 45388 31780 45444 31790
rect 45276 31778 45444 31780
rect 45276 31726 45390 31778
rect 45442 31726 45444 31778
rect 45276 31724 45444 31726
rect 45164 30660 45220 30670
rect 44940 30658 45220 30660
rect 44940 30606 45166 30658
rect 45218 30606 45220 30658
rect 44940 30604 45220 30606
rect 45164 30594 45220 30604
rect 44716 29822 44718 29874
rect 44770 29822 44772 29874
rect 44716 29810 44772 29822
rect 45052 29764 45108 29774
rect 45276 29764 45332 31724
rect 45388 31714 45444 31724
rect 45948 30770 46004 32732
rect 46060 32788 46116 32798
rect 46172 32788 46228 33740
rect 46060 32786 46228 32788
rect 46060 32734 46062 32786
rect 46114 32734 46228 32786
rect 46060 32732 46228 32734
rect 46060 32722 46116 32732
rect 46620 32674 46676 33740
rect 46620 32622 46622 32674
rect 46674 32622 46676 32674
rect 46620 31948 46676 32622
rect 46508 31892 46676 31948
rect 46732 33684 46788 33694
rect 46788 33628 47012 33684
rect 46060 31780 46116 31790
rect 46060 31686 46116 31724
rect 45948 30718 45950 30770
rect 46002 30718 46004 30770
rect 45948 30706 46004 30718
rect 46508 30770 46564 31892
rect 46508 30718 46510 30770
rect 46562 30718 46564 30770
rect 45500 30548 45556 30558
rect 45500 30454 45556 30492
rect 46284 30436 46340 30446
rect 45724 29988 45780 29998
rect 45724 29894 45780 29932
rect 45388 29876 45444 29886
rect 45388 29782 45444 29820
rect 46284 29874 46340 30380
rect 46284 29822 46286 29874
rect 46338 29822 46340 29874
rect 45052 29762 45332 29764
rect 45052 29710 45054 29762
rect 45106 29710 45332 29762
rect 45052 29708 45332 29710
rect 45052 29698 45108 29708
rect 43036 29090 43092 29102
rect 43036 29038 43038 29090
rect 43090 29038 43092 29090
rect 43036 28866 43092 29038
rect 43036 28814 43038 28866
rect 43090 28814 43092 28866
rect 43036 28802 43092 28814
rect 42812 27918 42814 27970
rect 42866 27918 42868 27970
rect 42812 27860 42868 27918
rect 43260 28420 43316 29596
rect 44380 29650 44436 29662
rect 44380 29598 44382 29650
rect 44434 29598 44436 29650
rect 43260 27972 43316 28364
rect 43260 27878 43316 27916
rect 44268 29540 44324 29550
rect 42812 27794 42868 27804
rect 43596 27860 43652 27870
rect 43596 27636 43652 27804
rect 43708 27636 43764 27646
rect 43372 27634 43764 27636
rect 43372 27582 43710 27634
rect 43762 27582 43764 27634
rect 43372 27580 43764 27582
rect 43372 26850 43428 27580
rect 43708 27570 43764 27580
rect 43372 26798 43374 26850
rect 43426 26798 43428 26850
rect 43372 26786 43428 26798
rect 44268 26850 44324 29484
rect 44380 29428 44436 29598
rect 44380 29362 44436 29372
rect 44716 28532 44772 28542
rect 44716 27970 44772 28476
rect 44716 27918 44718 27970
rect 44770 27918 44772 27970
rect 44716 27906 44772 27918
rect 45052 28530 45108 28542
rect 45052 28478 45054 28530
rect 45106 28478 45108 28530
rect 45052 28420 45108 28478
rect 45164 28532 45220 29708
rect 45948 28978 46004 28990
rect 45948 28926 45950 28978
rect 46002 28926 46004 28978
rect 45948 28866 46004 28926
rect 45948 28814 45950 28866
rect 46002 28814 46004 28866
rect 45948 28802 46004 28814
rect 45500 28532 45556 28542
rect 45164 28476 45444 28532
rect 45052 27972 45108 28364
rect 45164 27972 45220 27982
rect 45052 27916 45164 27972
rect 45164 27878 45220 27916
rect 44268 26798 44270 26850
rect 44322 26798 44324 26850
rect 44268 26740 44324 26798
rect 44716 26852 44772 26862
rect 44716 26758 44772 26796
rect 44268 26674 44324 26684
rect 42924 26628 42980 26638
rect 45164 26628 45220 26638
rect 42924 26534 42980 26572
rect 44828 26626 45220 26628
rect 44828 26574 45166 26626
rect 45218 26574 45220 26626
rect 44828 26572 45220 26574
rect 43932 26514 43988 26526
rect 43932 26462 43934 26514
rect 43986 26462 43988 26514
rect 42364 25790 42366 25842
rect 42418 25790 42420 25842
rect 42364 24778 42420 25790
rect 43820 25844 43876 25854
rect 43820 25750 43876 25788
rect 42476 25732 42532 25742
rect 42532 25676 42868 25732
rect 42476 25666 42532 25676
rect 42364 24726 42366 24778
rect 42418 24726 42420 24778
rect 42364 24164 42420 24726
rect 42812 24610 42868 25676
rect 43708 25618 43764 25630
rect 43708 25566 43710 25618
rect 43762 25566 43764 25618
rect 43708 25508 43764 25566
rect 43820 25508 43876 25518
rect 43932 25508 43988 26462
rect 44828 26066 44884 26572
rect 45164 26562 45220 26572
rect 44828 26014 44830 26066
rect 44882 26014 44884 26066
rect 44828 26002 44884 26014
rect 45388 25842 45444 28476
rect 45500 27972 45556 28476
rect 45612 27972 45668 27982
rect 45500 27970 45668 27972
rect 45500 27918 45614 27970
rect 45666 27918 45668 27970
rect 45500 27916 45668 27918
rect 45612 27860 45668 27916
rect 46060 27972 46116 27982
rect 46060 27878 46116 27916
rect 46284 27860 46340 29822
rect 46396 29428 46452 29438
rect 46396 28868 46452 29372
rect 46508 28978 46564 30718
rect 46620 31778 46676 31790
rect 46620 31726 46622 31778
rect 46674 31726 46676 31778
rect 46620 30436 46676 31726
rect 46620 30370 46676 30380
rect 46732 30212 46788 33628
rect 46844 33458 46900 33470
rect 46844 33406 46846 33458
rect 46898 33406 46900 33458
rect 46844 32786 46900 33406
rect 46956 33012 47012 33628
rect 47292 33012 47348 40462
rect 48300 40292 48356 40686
rect 49084 40628 49140 40638
rect 48300 40236 48692 40292
rect 48636 40178 48692 40236
rect 48636 40126 48638 40178
rect 48690 40126 48692 40178
rect 48636 40114 48692 40126
rect 49084 39954 49140 40572
rect 49196 40626 49252 40638
rect 49196 40574 49198 40626
rect 49250 40574 49252 40626
rect 49196 40516 49252 40574
rect 49196 40450 49252 40460
rect 49084 39902 49086 39954
rect 49138 39902 49140 39954
rect 49084 39890 49140 39902
rect 48188 39844 48244 39854
rect 49308 39844 49364 40796
rect 49420 40786 49476 40796
rect 49532 40740 49588 40750
rect 49532 40646 49588 40684
rect 49756 40516 49812 42590
rect 50092 41860 50148 45388
rect 50204 44884 50260 47742
rect 50428 47740 50652 47796
rect 50316 45890 50372 45902
rect 50316 45838 50318 45890
rect 50370 45838 50372 45890
rect 50316 45444 50372 45838
rect 50428 45668 50484 47740
rect 50652 47702 50708 47740
rect 52108 47794 52164 47806
rect 52668 47796 52724 47806
rect 52108 47742 52110 47794
rect 52162 47742 52164 47794
rect 52108 47682 52164 47742
rect 52108 47630 52110 47682
rect 52162 47630 52164 47682
rect 50988 46564 51044 46574
rect 50876 46562 51044 46564
rect 50876 46510 50990 46562
rect 51042 46510 51044 46562
rect 50876 46508 51044 46510
rect 50556 46396 50820 46406
rect 50612 46340 50660 46396
rect 50716 46340 50764 46396
rect 50556 46330 50820 46340
rect 50876 46002 50932 46508
rect 50988 46498 51044 46508
rect 50876 45950 50878 46002
rect 50930 45950 50932 46002
rect 50876 45938 50932 45950
rect 51548 46002 51604 46014
rect 51548 45950 51550 46002
rect 51602 45950 51604 46002
rect 50428 45612 50708 45668
rect 50316 45378 50372 45388
rect 50204 43764 50260 44828
rect 50652 44770 50708 45612
rect 50988 44884 51044 44894
rect 50652 44718 50654 44770
rect 50706 44718 50708 44770
rect 50652 44660 50708 44718
rect 50652 44594 50708 44604
rect 50876 44772 50932 44782
rect 50556 44380 50820 44390
rect 50612 44324 50660 44380
rect 50716 44324 50764 44380
rect 50556 44314 50820 44324
rect 50876 43876 50932 44716
rect 50876 43708 50932 43820
rect 50204 43698 50260 43708
rect 50316 43652 50932 43708
rect 50988 43708 51044 44828
rect 51212 44772 51268 44782
rect 51212 44678 51268 44716
rect 51436 44660 51492 44670
rect 51436 44566 51492 44604
rect 50988 43652 51156 43708
rect 50204 42868 50260 42878
rect 50204 42774 50260 42812
rect 49868 41746 49924 41758
rect 49868 41694 49870 41746
rect 49922 41694 49924 41746
rect 49868 41522 49924 41694
rect 49868 41470 49870 41522
rect 49922 41470 49924 41522
rect 49868 41458 49924 41470
rect 49756 40450 49812 40460
rect 49980 40738 50036 40750
rect 49980 40686 49982 40738
rect 50034 40686 50036 40738
rect 47516 39620 47572 39630
rect 47516 39526 47572 39564
rect 48188 38948 48244 39788
rect 48188 38882 48244 38892
rect 49196 39788 49364 39844
rect 49420 40292 49476 40302
rect 49420 39842 49476 40236
rect 49980 40068 50036 40686
rect 49980 40002 50036 40012
rect 49420 39790 49422 39842
rect 49474 39790 49476 39842
rect 47628 38834 47684 38846
rect 47628 38782 47630 38834
rect 47682 38782 47684 38834
rect 47628 38724 47684 38782
rect 48636 38836 48692 38846
rect 47628 38162 47684 38668
rect 48188 38724 48244 38762
rect 48188 38658 48244 38668
rect 48636 38722 48692 38780
rect 48972 38836 49028 38846
rect 49196 38836 49252 39788
rect 49420 39778 49476 39790
rect 49644 39954 49700 39966
rect 49644 39902 49646 39954
rect 49698 39902 49700 39954
rect 48972 38834 49252 38836
rect 48972 38782 48974 38834
rect 49026 38782 49252 38834
rect 48972 38780 49252 38782
rect 48972 38770 49028 38780
rect 48636 38670 48638 38722
rect 48690 38670 48692 38722
rect 48636 38658 48692 38670
rect 49196 38612 49252 38780
rect 49308 39620 49364 39630
rect 49308 38834 49364 39564
rect 49308 38782 49310 38834
rect 49362 38782 49364 38834
rect 49308 38770 49364 38782
rect 49644 38834 49700 39902
rect 49644 38782 49646 38834
rect 49698 38782 49700 38834
rect 49644 38770 49700 38782
rect 50092 38724 50148 41804
rect 50316 41748 50372 43652
rect 50652 43202 50708 43214
rect 50652 43150 50654 43202
rect 50706 43150 50708 43202
rect 50652 42642 50708 43150
rect 50652 42590 50654 42642
rect 50706 42590 50708 42642
rect 50652 42578 50708 42590
rect 51100 42642 51156 43652
rect 51548 43202 51604 45950
rect 52108 45780 52164 47630
rect 52556 47794 52724 47796
rect 52556 47742 52670 47794
rect 52722 47742 52724 47794
rect 52556 47740 52724 47742
rect 52332 45780 52388 45790
rect 52108 45778 52388 45780
rect 52108 45726 52334 45778
rect 52386 45726 52388 45778
rect 52108 45724 52388 45726
rect 52332 45220 52388 45724
rect 52556 45444 52612 47740
rect 52668 47730 52724 47740
rect 53004 47794 53060 47806
rect 53004 47742 53006 47794
rect 53058 47742 53060 47794
rect 53004 47682 53060 47742
rect 53452 47796 53508 47806
rect 53452 47702 53508 47740
rect 53004 47630 53006 47682
rect 53058 47630 53060 47682
rect 53004 47618 53060 47630
rect 52780 46900 52836 46910
rect 53676 46900 53732 46910
rect 52780 46898 53732 46900
rect 52780 46846 52782 46898
rect 52834 46846 53678 46898
rect 53730 46846 53732 46898
rect 52780 46844 53732 46846
rect 52780 46834 52836 46844
rect 53004 46004 53060 46844
rect 53676 46834 53732 46844
rect 53228 46674 53284 46686
rect 53228 46622 53230 46674
rect 53282 46622 53284 46674
rect 53228 46562 53284 46622
rect 54124 46674 54180 46686
rect 54124 46622 54126 46674
rect 54178 46622 54180 46674
rect 53228 46510 53230 46562
rect 53282 46510 53284 46562
rect 53228 46498 53284 46510
rect 53788 46562 53844 46574
rect 53788 46510 53790 46562
rect 53842 46510 53844 46562
rect 53788 46004 53844 46510
rect 53004 46002 53172 46004
rect 53004 45950 53006 46002
rect 53058 45950 53172 46002
rect 53004 45948 53172 45950
rect 53004 45938 53060 45948
rect 52556 45378 52612 45388
rect 52668 45332 52724 45342
rect 52724 45276 53060 45332
rect 52668 45266 52724 45276
rect 51884 44772 51940 44782
rect 51884 44678 51940 44716
rect 51884 43988 51940 43998
rect 51884 43894 51940 43932
rect 52332 43876 52388 45164
rect 53004 44882 53060 45276
rect 53004 44830 53006 44882
rect 53058 44830 53060 44882
rect 52668 44772 52724 44782
rect 52668 44678 52724 44716
rect 52332 43810 52388 43820
rect 52892 43876 52948 43886
rect 52892 43782 52948 43820
rect 51548 43150 51550 43202
rect 51602 43150 51604 43202
rect 51548 43138 51604 43150
rect 51100 42590 51102 42642
rect 51154 42590 51156 42642
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50540 42196 50596 42206
rect 50428 41748 50484 41758
rect 50316 41746 50484 41748
rect 50316 41694 50430 41746
rect 50482 41694 50484 41746
rect 50316 41692 50484 41694
rect 50428 41636 50484 41692
rect 50204 40516 50260 40526
rect 50204 39954 50260 40460
rect 50204 39902 50206 39954
rect 50258 39902 50260 39954
rect 50204 39890 50260 39902
rect 50428 39842 50484 41580
rect 50540 40738 50596 42140
rect 50876 42084 50932 42094
rect 50876 41990 50932 42028
rect 50876 41522 50932 41534
rect 50876 41470 50878 41522
rect 50930 41470 50932 41522
rect 50540 40686 50542 40738
rect 50594 40686 50596 40738
rect 50540 40674 50596 40686
rect 50652 40738 50708 40750
rect 50652 40686 50654 40738
rect 50706 40686 50708 40738
rect 50540 40516 50596 40526
rect 50652 40516 50708 40686
rect 50596 40460 50708 40516
rect 50540 40450 50596 40460
rect 50556 40348 50820 40358
rect 50612 40292 50660 40348
rect 50716 40292 50764 40348
rect 50556 40282 50820 40292
rect 50652 39848 50708 39860
rect 50652 39844 50654 39848
rect 50428 39790 50430 39842
rect 50482 39790 50484 39842
rect 50428 38836 50484 39790
rect 50428 38770 50484 38780
rect 50540 39796 50654 39844
rect 50706 39844 50708 39848
rect 50764 39844 50820 39854
rect 50706 39796 50764 39844
rect 50540 39788 50764 39796
rect 50092 38722 50372 38724
rect 50092 38670 50094 38722
rect 50146 38670 50372 38722
rect 50092 38668 50372 38670
rect 50092 38658 50148 38668
rect 49756 38612 49812 38622
rect 49196 38556 49588 38612
rect 49084 38500 49140 38510
rect 47628 38110 47630 38162
rect 47682 38110 47684 38162
rect 47628 38098 47684 38110
rect 48188 38162 48244 38174
rect 48188 38110 48190 38162
rect 48242 38110 48244 38162
rect 47740 38052 47796 38062
rect 47740 37958 47796 37996
rect 48188 38050 48244 38110
rect 48188 37998 48190 38050
rect 48242 37998 48244 38050
rect 48188 37940 48244 37998
rect 48188 36818 48244 37884
rect 49084 37940 49140 38444
rect 49084 37846 49140 37884
rect 48188 36766 48190 36818
rect 48242 36766 48244 36818
rect 47852 36706 47908 36718
rect 47852 36654 47854 36706
rect 47906 36654 47908 36706
rect 47852 36596 47908 36654
rect 47852 36530 47908 36540
rect 48188 34916 48244 36766
rect 49084 37156 49140 37166
rect 49084 36594 49140 37100
rect 49532 36930 49588 38556
rect 49756 38052 49812 38556
rect 49756 37958 49812 37996
rect 50316 37042 50372 38668
rect 50540 38500 50596 39788
rect 50652 39784 50708 39788
rect 50764 39778 50820 39788
rect 50876 39842 50932 41470
rect 51100 41522 51156 42590
rect 51548 42642 51604 42654
rect 51996 42644 52052 42654
rect 51548 42590 51550 42642
rect 51602 42590 51604 42642
rect 51100 41470 51102 41522
rect 51154 41470 51156 41522
rect 51100 41458 51156 41470
rect 51212 42084 51268 42094
rect 51212 40964 51268 42028
rect 51548 42084 51604 42590
rect 51548 42018 51604 42028
rect 51884 42588 51996 42644
rect 51324 41748 51380 41758
rect 51324 41522 51380 41692
rect 51324 41470 51326 41522
rect 51378 41470 51380 41522
rect 51324 41458 51380 41470
rect 50876 39790 50878 39842
rect 50930 39790 50932 39842
rect 50876 38948 50932 39790
rect 50316 36990 50318 37042
rect 50370 36990 50372 37042
rect 50316 36978 50372 36990
rect 50428 38444 50596 38500
rect 50652 38892 50932 38948
rect 51100 40962 51268 40964
rect 51100 40910 51214 40962
rect 51266 40910 51268 40962
rect 51100 40908 51268 40910
rect 51100 39956 51156 40908
rect 51212 40898 51268 40908
rect 51884 40068 51940 42588
rect 51996 42550 52052 42588
rect 52668 42082 52724 42094
rect 52668 42030 52670 42082
rect 52722 42030 52724 42082
rect 52220 41972 52276 41982
rect 52220 41878 52276 41916
rect 51996 41860 52052 41870
rect 51996 40962 52052 41804
rect 52332 41858 52388 41870
rect 52332 41806 52334 41858
rect 52386 41806 52388 41858
rect 52332 41748 52388 41806
rect 52332 41682 52388 41692
rect 51996 40910 51998 40962
rect 52050 40910 52052 40962
rect 51996 40898 52052 40910
rect 52668 40850 52724 42030
rect 52668 40798 52670 40850
rect 52722 40798 52724 40850
rect 52668 40786 52724 40798
rect 53004 40852 53060 44830
rect 53004 40758 53060 40796
rect 53116 44660 53172 45948
rect 53788 45910 53844 45948
rect 53452 45890 53508 45902
rect 53452 45838 53454 45890
rect 53506 45838 53508 45890
rect 53452 45220 53508 45838
rect 54012 45890 54068 45902
rect 54012 45838 54014 45890
rect 54066 45838 54068 45890
rect 53452 45154 53508 45164
rect 53676 45778 53732 45790
rect 53676 45726 53678 45778
rect 53730 45726 53732 45778
rect 53676 44884 53732 45726
rect 53676 44818 53732 44828
rect 53116 43986 53172 44604
rect 53116 43934 53118 43986
rect 53170 43934 53172 43986
rect 53116 42868 53172 43934
rect 53340 44770 53396 44782
rect 53340 44718 53342 44770
rect 53394 44718 53396 44770
rect 53340 43988 53396 44718
rect 53340 43922 53396 43932
rect 53676 44658 53732 44670
rect 53676 44606 53678 44658
rect 53730 44606 53732 44658
rect 53228 42868 53284 42878
rect 53172 42866 53284 42868
rect 53172 42814 53230 42866
rect 53282 42814 53284 42866
rect 53172 42812 53284 42814
rect 51884 40012 52052 40068
rect 51100 39954 51828 39956
rect 51100 39902 51102 39954
rect 51154 39902 51828 39954
rect 51100 39900 51828 39902
rect 50652 38500 50708 38892
rect 50764 38724 50820 38734
rect 50764 38630 50820 38668
rect 51100 38612 51156 39900
rect 51772 39842 51828 39900
rect 51772 39790 51774 39842
rect 51826 39790 51828 39842
rect 51772 39778 51828 39790
rect 51996 39844 52052 40012
rect 51212 39508 51268 39518
rect 51212 39506 51492 39508
rect 51212 39454 51214 39506
rect 51266 39454 51492 39506
rect 51212 39452 51492 39454
rect 51212 39442 51268 39452
rect 51436 38722 51492 39452
rect 51996 38948 52052 39788
rect 51996 38882 52052 38892
rect 52108 39842 52164 39854
rect 52108 39790 52110 39842
rect 52162 39790 52164 39842
rect 52108 38724 52164 39790
rect 52444 39844 52500 39854
rect 52892 39844 52948 39854
rect 52444 39842 52948 39844
rect 52444 39790 52446 39842
rect 52498 39790 52894 39842
rect 52946 39790 52948 39842
rect 52444 39788 52948 39790
rect 52444 39778 52500 39788
rect 52892 39778 52948 39788
rect 51436 38670 51438 38722
rect 51490 38670 51492 38722
rect 51436 38658 51492 38670
rect 51772 38668 52108 38724
rect 51100 38546 51156 38556
rect 49532 36878 49534 36930
rect 49586 36878 49588 36930
rect 49532 36866 49588 36878
rect 49868 36708 49924 36718
rect 49868 36706 50036 36708
rect 49868 36654 49870 36706
rect 49922 36654 50036 36706
rect 49868 36652 50036 36654
rect 49868 36642 49924 36652
rect 49084 36542 49086 36594
rect 49138 36542 49140 36594
rect 49084 36530 49140 36542
rect 49420 35924 49476 35934
rect 49420 35830 49476 35868
rect 48972 35700 49028 35710
rect 48972 35606 49028 35644
rect 48188 34018 48244 34860
rect 49420 34916 49476 34926
rect 49420 34822 49476 34860
rect 48188 33966 48190 34018
rect 48242 33966 48244 34018
rect 48188 33954 48244 33966
rect 48860 34804 48916 34814
rect 46956 32956 47236 33012
rect 46844 32734 46846 32786
rect 46898 32734 46900 32786
rect 46844 32722 46900 32734
rect 47068 32788 47124 32798
rect 47180 32788 47236 32956
rect 47292 32946 47348 32956
rect 48860 33796 48916 34748
rect 49868 34804 49924 34814
rect 49868 34710 49924 34748
rect 49980 34692 50036 36652
rect 50204 36596 50260 36606
rect 50204 35924 50260 36540
rect 50092 35700 50148 35710
rect 50092 35606 50148 35644
rect 49980 34626 50036 34636
rect 50204 34580 50260 35868
rect 50316 34580 50372 34590
rect 50204 34578 50372 34580
rect 50204 34526 50318 34578
rect 50370 34526 50372 34578
rect 50204 34524 50372 34526
rect 50204 34130 50260 34142
rect 50204 34078 50206 34130
rect 50258 34078 50260 34130
rect 50204 34018 50260 34078
rect 50204 33966 50206 34018
rect 50258 33966 50260 34018
rect 50204 33954 50260 33966
rect 47292 32788 47348 32798
rect 47180 32786 47348 32788
rect 47180 32734 47294 32786
rect 47346 32734 47348 32786
rect 47180 32732 47348 32734
rect 47068 32694 47124 32732
rect 47292 32722 47348 32732
rect 47964 32676 48020 32686
rect 48412 32676 48468 32686
rect 47964 32674 48468 32676
rect 47964 32622 47966 32674
rect 48018 32622 48414 32674
rect 48466 32622 48468 32674
rect 47964 32620 48468 32622
rect 46732 29428 46788 30156
rect 46844 32562 46900 32574
rect 46844 32510 46846 32562
rect 46898 32510 46900 32562
rect 46844 29874 46900 32510
rect 47628 32562 47684 32574
rect 47628 32510 47630 32562
rect 47682 32510 47684 32562
rect 47628 31948 47684 32510
rect 46844 29822 46846 29874
rect 46898 29822 46900 29874
rect 46844 29810 46900 29822
rect 47068 31892 47684 31948
rect 47068 29764 47124 31892
rect 47852 31890 47908 31902
rect 47852 31838 47854 31890
rect 47906 31838 47908 31890
rect 47180 31778 47236 31790
rect 47180 31726 47182 31778
rect 47234 31726 47236 31778
rect 47180 30436 47236 31726
rect 47852 31668 47908 31838
rect 47852 31602 47908 31612
rect 47964 31780 48020 32620
rect 48412 32610 48468 32620
rect 48860 31890 48916 33740
rect 49868 33460 49924 33470
rect 48860 31838 48862 31890
rect 48914 31838 48916 31890
rect 48860 31826 48916 31838
rect 48972 32676 49028 32686
rect 49756 32676 49812 32686
rect 48972 32674 49812 32676
rect 48972 32622 48974 32674
rect 49026 32622 49758 32674
rect 49810 32622 49812 32674
rect 48972 32620 49812 32622
rect 47964 30772 48020 31724
rect 48748 31668 48804 31678
rect 48748 31574 48804 31612
rect 47964 30706 48020 30716
rect 48748 30658 48804 30670
rect 48748 30606 48750 30658
rect 48802 30606 48804 30658
rect 48188 30548 48244 30558
rect 47628 30436 47684 30446
rect 47180 30434 47684 30436
rect 47180 30382 47630 30434
rect 47682 30382 47684 30434
rect 47180 30380 47684 30382
rect 47628 30370 47684 30380
rect 47516 29874 47572 29886
rect 47516 29822 47518 29874
rect 47570 29822 47572 29874
rect 47068 29698 47124 29708
rect 47404 29764 47460 29774
rect 46732 29362 46788 29372
rect 46508 28926 46510 28978
rect 46562 28926 46564 28978
rect 46508 28914 46564 28926
rect 46844 28978 46900 28990
rect 46844 28926 46846 28978
rect 46898 28926 46900 28978
rect 46396 28774 46452 28812
rect 46508 27972 46564 27982
rect 46284 27804 46452 27860
rect 45612 27794 45668 27804
rect 46284 27636 46340 27646
rect 46172 27634 46340 27636
rect 46172 27582 46286 27634
rect 46338 27582 46340 27634
rect 46172 27580 46340 27582
rect 46172 26852 46228 27580
rect 46284 27570 46340 27580
rect 46396 27076 46452 27804
rect 46508 27858 46564 27916
rect 46508 27806 46510 27858
rect 46562 27806 46564 27858
rect 46508 27794 46564 27806
rect 46844 27970 46900 28926
rect 47068 28868 47124 28878
rect 47068 28754 47124 28812
rect 47068 28702 47070 28754
rect 47122 28702 47124 28754
rect 47068 28690 47124 28702
rect 46844 27918 46846 27970
rect 46898 27918 46900 27970
rect 45724 26796 46228 26852
rect 46284 27020 46452 27076
rect 45500 26740 45556 26750
rect 45500 26646 45556 26684
rect 45612 26628 45668 26638
rect 45612 26534 45668 26572
rect 45388 25790 45390 25842
rect 45442 25790 45444 25842
rect 45388 25778 45444 25790
rect 45612 25844 45668 25854
rect 44380 25732 44436 25742
rect 44380 25638 44436 25676
rect 45052 25730 45108 25742
rect 45052 25678 45054 25730
rect 45106 25678 45108 25730
rect 43708 25452 43820 25508
rect 43876 25452 43988 25508
rect 42812 24558 42814 24610
rect 42866 24558 42868 24610
rect 42812 24546 42868 24558
rect 42420 24108 42644 24164
rect 42364 24098 42420 24108
rect 42252 23774 42254 23826
rect 42306 23774 42308 23826
rect 42252 23762 42308 23774
rect 42476 23940 42532 23950
rect 42476 23826 42532 23884
rect 42476 23774 42478 23826
rect 42530 23774 42532 23826
rect 42476 23762 42532 23774
rect 42140 23662 42142 23714
rect 42194 23662 42196 23714
rect 42140 23650 42196 23662
rect 42588 22820 42644 24108
rect 41916 22726 41972 22764
rect 42140 22818 42644 22820
rect 42140 22766 42590 22818
rect 42642 22766 42644 22818
rect 42140 22764 42644 22766
rect 41580 22708 41636 22718
rect 41580 22706 41748 22708
rect 41580 22654 41582 22706
rect 41634 22654 41748 22706
rect 41580 22652 41748 22654
rect 41580 22642 41636 22652
rect 41020 21980 41412 22036
rect 41020 21922 41076 21980
rect 41020 21870 41022 21922
rect 41074 21870 41076 21922
rect 41020 21858 41076 21870
rect 40348 21532 40740 21588
rect 41132 21812 41188 21822
rect 40124 20916 40180 20926
rect 40012 20580 40068 20590
rect 40012 20486 40068 20524
rect 39116 18788 39172 18798
rect 39228 18788 39284 19628
rect 39172 18732 39284 18788
rect 39452 20132 39620 20188
rect 39452 19796 39508 20132
rect 39116 18694 39172 18732
rect 38780 17892 38836 18620
rect 39452 18562 39508 19740
rect 40012 19460 40068 19470
rect 39452 18510 39454 18562
rect 39506 18510 39508 18562
rect 39452 18498 39508 18510
rect 39900 19458 40068 19460
rect 39900 19406 40014 19458
rect 40066 19406 40068 19458
rect 39900 19404 40068 19406
rect 39788 18452 39844 18462
rect 39788 18358 39844 18396
rect 39900 18228 39956 19404
rect 40012 19394 40068 19404
rect 40124 18788 40180 20860
rect 40348 20690 40404 21532
rect 40684 20916 40740 20926
rect 40684 20822 40740 20860
rect 41132 20802 41188 21756
rect 41132 20750 41134 20802
rect 41186 20750 41188 20802
rect 41132 20692 41188 20750
rect 40348 20638 40350 20690
rect 40402 20638 40404 20690
rect 40348 19794 40404 20638
rect 40348 19742 40350 19794
rect 40402 19742 40404 19794
rect 40348 19730 40404 19742
rect 40908 20636 41188 20692
rect 41244 21700 41300 21710
rect 39788 18172 39956 18228
rect 40012 18732 40180 18788
rect 40908 19682 40964 20636
rect 40908 19630 40910 19682
rect 40962 19630 40964 19682
rect 38780 17826 38836 17836
rect 39452 17892 39508 17902
rect 39452 17798 39508 17836
rect 36764 17556 36820 17594
rect 36764 17490 36820 17500
rect 39788 17556 39844 18172
rect 39900 17892 39956 17902
rect 39900 17798 39956 17836
rect 36652 15598 36654 15650
rect 36706 15598 36708 15650
rect 36428 14980 36484 14990
rect 36428 14754 36484 14924
rect 36428 14702 36430 14754
rect 36482 14702 36484 14754
rect 36428 14690 36484 14702
rect 36652 14420 36708 15598
rect 36652 14354 36708 14364
rect 36764 17332 36820 17342
rect 36316 13806 36318 13858
rect 36370 13806 36372 13858
rect 36316 13794 36372 13806
rect 35644 13694 35646 13746
rect 35698 13694 35700 13746
rect 35644 13682 35700 13694
rect 36764 13746 36820 17276
rect 39228 16660 39284 16670
rect 39788 16660 39844 17500
rect 39900 16660 39956 16670
rect 39788 16604 39900 16660
rect 38556 16436 38612 16446
rect 37100 15876 37156 15886
rect 37100 15782 37156 15820
rect 37548 15764 37604 15774
rect 37548 15670 37604 15708
rect 38556 15762 38612 16380
rect 39228 15874 39284 16604
rect 39900 16594 39956 16604
rect 39676 16548 39732 16558
rect 39676 16546 39844 16548
rect 39676 16494 39678 16546
rect 39730 16494 39844 16546
rect 39676 16492 39844 16494
rect 39676 16482 39732 16492
rect 39228 15822 39230 15874
rect 39282 15822 39284 15874
rect 39228 15810 39284 15822
rect 38556 15710 38558 15762
rect 38610 15710 38612 15762
rect 38556 15698 38612 15710
rect 37996 15652 38052 15662
rect 37996 15558 38052 15596
rect 38668 15538 38724 15550
rect 38668 15486 38670 15538
rect 38722 15486 38724 15538
rect 37884 14980 37940 14990
rect 37324 14756 37380 14766
rect 37324 14662 37380 14700
rect 37772 14642 37828 14654
rect 37772 14590 37774 14642
rect 37826 14590 37828 14642
rect 37772 14420 37828 14590
rect 37884 14642 37940 14924
rect 38668 14756 38724 15486
rect 38668 14690 38724 14700
rect 37884 14590 37886 14642
rect 37938 14590 37940 14642
rect 37884 14578 37940 14590
rect 38220 14644 38276 14654
rect 38220 14550 38276 14588
rect 39004 14642 39060 14654
rect 39004 14590 39006 14642
rect 39058 14590 39060 14642
rect 37772 14084 37828 14364
rect 37772 14028 38388 14084
rect 38108 13860 38164 13870
rect 36764 13694 36766 13746
rect 36818 13694 36820 13746
rect 36764 13682 36820 13694
rect 36988 13858 38164 13860
rect 36988 13806 38110 13858
rect 38162 13806 38164 13858
rect 36988 13804 38164 13806
rect 35308 13636 35364 13646
rect 35980 13636 36036 13646
rect 35308 13634 35588 13636
rect 35308 13582 35310 13634
rect 35362 13582 35588 13634
rect 35308 13580 35588 13582
rect 35308 13570 35364 13580
rect 35196 13132 35460 13142
rect 35252 13076 35300 13132
rect 35356 13076 35404 13132
rect 35196 13066 35460 13076
rect 33404 12674 33460 12684
rect 33740 12740 33796 12750
rect 33740 12646 33796 12684
rect 35532 12628 35588 13580
rect 35980 13634 36260 13636
rect 35980 13582 35982 13634
rect 36034 13582 36260 13634
rect 35980 13580 36260 13582
rect 35980 13570 36036 13580
rect 36204 12628 36260 13580
rect 35532 12572 35700 12628
rect 36204 12572 36820 12628
rect 31724 11902 31726 11954
rect 31778 11902 31780 11954
rect 31724 11890 31780 11902
rect 32172 12514 32228 12526
rect 32172 12462 32174 12514
rect 32226 12462 32228 12514
rect 31164 11678 31166 11730
rect 31218 11678 31220 11730
rect 31164 11508 31220 11678
rect 31164 10724 31220 11452
rect 31612 11506 31668 11518
rect 31612 11454 31614 11506
rect 31666 11454 31668 11506
rect 31612 11282 31668 11454
rect 32060 11506 32116 11518
rect 32060 11454 32062 11506
rect 32114 11454 32116 11506
rect 31612 11230 31614 11282
rect 31666 11230 31668 11282
rect 31612 11218 31668 11230
rect 31948 11396 32004 11406
rect 32060 11396 32116 11454
rect 32004 11340 32116 11396
rect 31276 10724 31332 10734
rect 31724 10724 31780 10734
rect 31164 10722 31668 10724
rect 31164 10670 31278 10722
rect 31330 10670 31668 10722
rect 31164 10668 31668 10670
rect 31164 10164 31220 10668
rect 31276 10658 31332 10668
rect 31612 10610 31668 10668
rect 31612 10558 31614 10610
rect 31666 10558 31668 10610
rect 31612 10546 31668 10558
rect 31164 10098 31220 10108
rect 30156 9886 30158 9938
rect 30210 9886 30212 9938
rect 30156 9874 30212 9886
rect 29260 8372 29764 8428
rect 29596 7812 29652 8372
rect 31724 8370 31780 10668
rect 31948 8372 32004 11340
rect 32172 8818 32228 12462
rect 32844 12402 32900 12414
rect 32844 12350 32846 12402
rect 32898 12350 32900 12402
rect 32508 11506 32564 11518
rect 32508 11454 32510 11506
rect 32562 11454 32564 11506
rect 32396 11282 32452 11294
rect 32396 11230 32398 11282
rect 32450 11230 32452 11282
rect 32396 10500 32452 11230
rect 32508 10612 32564 11454
rect 32508 10546 32564 10556
rect 32396 10406 32452 10444
rect 32172 8766 32174 8818
rect 32226 8766 32228 8818
rect 32172 8754 32228 8766
rect 32844 8428 32900 12350
rect 35532 12404 35588 12414
rect 35532 12310 35588 12348
rect 33628 11618 33684 11630
rect 33628 11566 33630 11618
rect 33682 11566 33684 11618
rect 33068 11508 33124 11518
rect 33124 11452 33572 11508
rect 33068 11414 33124 11452
rect 33516 9938 33572 11452
rect 33628 10500 33684 11566
rect 35196 11116 35460 11126
rect 35252 11060 35300 11116
rect 35356 11060 35404 11116
rect 35196 11050 35460 11060
rect 35644 10948 35700 12572
rect 35980 12404 36036 12414
rect 35980 12310 36036 12348
rect 36428 12402 36484 12414
rect 36428 12350 36430 12402
rect 36482 12350 36484 12402
rect 36316 11620 36372 11630
rect 36428 11620 36484 12350
rect 36764 11730 36820 12572
rect 36764 11678 36766 11730
rect 36818 11678 36820 11730
rect 36764 11666 36820 11678
rect 36316 11618 36484 11620
rect 36316 11566 36318 11618
rect 36370 11566 36484 11618
rect 36316 11564 36484 11566
rect 36316 11554 36372 11564
rect 35308 10892 35700 10948
rect 35868 11506 35924 11518
rect 35868 11454 35870 11506
rect 35922 11454 35924 11506
rect 35868 11396 35924 11454
rect 35308 10834 35364 10892
rect 35308 10782 35310 10834
rect 35362 10782 35364 10834
rect 35308 10770 35364 10782
rect 35868 10724 35924 11340
rect 35980 10724 36036 10734
rect 35868 10668 35980 10724
rect 35980 10630 36036 10668
rect 36428 10722 36484 11564
rect 36988 10946 37044 13804
rect 38108 13794 38164 13804
rect 37436 13634 37492 13646
rect 37436 13582 37438 13634
rect 37490 13582 37492 13634
rect 37324 12404 37380 12414
rect 36988 10894 36990 10946
rect 37042 10894 37044 10946
rect 36988 10882 37044 10894
rect 37100 12348 37324 12404
rect 36428 10670 36430 10722
rect 36482 10670 36484 10722
rect 34188 10612 34244 10622
rect 36428 10612 36484 10670
rect 36540 10612 36596 10622
rect 36428 10556 36540 10612
rect 34188 10518 34244 10556
rect 36540 10546 36596 10556
rect 33628 10052 33684 10444
rect 33964 10052 34020 10062
rect 33628 9996 33964 10052
rect 33516 9886 33518 9938
rect 33570 9886 33572 9938
rect 33516 9826 33572 9886
rect 33516 9774 33518 9826
rect 33570 9774 33572 9826
rect 33516 9762 33572 9774
rect 33964 9826 34020 9996
rect 35196 10052 35252 10062
rect 33964 9774 33966 9826
rect 34018 9774 34020 9826
rect 33964 9762 34020 9774
rect 34524 9938 34580 9950
rect 34524 9886 34526 9938
rect 34578 9886 34580 9938
rect 34524 9602 34580 9886
rect 34524 9550 34526 9602
rect 34578 9550 34580 9602
rect 34524 9538 34580 9550
rect 35196 9602 35252 9996
rect 35196 9550 35198 9602
rect 35250 9550 35252 9602
rect 35196 9538 35252 9550
rect 36428 10052 36484 10062
rect 35196 9100 35460 9110
rect 35252 9044 35300 9100
rect 35356 9044 35404 9100
rect 35196 9034 35460 9044
rect 36428 8706 36484 9996
rect 36428 8654 36430 8706
rect 36482 8654 36484 8706
rect 36428 8642 36484 8654
rect 37100 8706 37156 12348
rect 37324 12310 37380 12348
rect 37324 11506 37380 11518
rect 37324 11454 37326 11506
rect 37378 11454 37380 11506
rect 37324 10836 37380 11454
rect 37324 10164 37380 10780
rect 37324 10098 37380 10108
rect 37436 9492 37492 13582
rect 38332 12516 38388 14028
rect 38892 13636 38948 13646
rect 39004 13636 39060 14590
rect 38892 13634 39004 13636
rect 38892 13582 38894 13634
rect 38946 13582 39004 13634
rect 38892 13580 39004 13582
rect 38444 12516 38500 12526
rect 38332 12514 38500 12516
rect 38332 12462 38446 12514
rect 38498 12462 38500 12514
rect 38332 12460 38500 12462
rect 37660 12404 37716 12414
rect 37660 11730 37716 12348
rect 37660 11678 37662 11730
rect 37714 11678 37716 11730
rect 37660 11666 37716 11678
rect 37772 12402 37828 12414
rect 37772 12350 37774 12402
rect 37826 12350 37828 12402
rect 37772 11732 37828 12350
rect 38220 12404 38276 12414
rect 38220 12310 38276 12348
rect 37772 10724 37828 11676
rect 37772 10610 37828 10668
rect 37772 10558 37774 10610
rect 37826 10558 37828 10610
rect 37772 10546 37828 10558
rect 38332 10612 38388 12460
rect 38444 12450 38500 12460
rect 38556 12514 38612 12526
rect 38556 12462 38558 12514
rect 38610 12462 38612 12514
rect 38556 11732 38612 12462
rect 38556 11666 38612 11676
rect 38892 12404 38948 13580
rect 39004 13570 39060 13580
rect 39452 13636 39508 13646
rect 39452 12626 39508 13580
rect 39788 13522 39844 16492
rect 40012 16546 40068 18732
rect 40124 18564 40180 18574
rect 40124 18470 40180 18508
rect 40348 17556 40404 17566
rect 40348 16772 40404 17500
rect 40908 17556 40964 19630
rect 41020 19684 41076 19694
rect 41020 19590 41076 19628
rect 41020 19012 41076 19022
rect 41244 19012 41300 21644
rect 41020 19010 41300 19012
rect 41020 18958 41022 19010
rect 41074 18958 41300 19010
rect 41020 18956 41300 18958
rect 41356 19684 41412 21980
rect 41580 21586 41636 21598
rect 41580 21534 41582 21586
rect 41634 21534 41636 21586
rect 41468 21476 41524 21486
rect 41468 21382 41524 21420
rect 41580 21364 41636 21534
rect 41580 21298 41636 21308
rect 41692 21588 41748 22652
rect 42140 22706 42196 22764
rect 42588 22754 42644 22764
rect 43036 22820 43092 22830
rect 43036 22726 43092 22764
rect 43484 22820 43540 22830
rect 43484 22726 43540 22764
rect 42140 22654 42142 22706
rect 42194 22654 42196 22706
rect 42140 22642 42196 22654
rect 41580 20580 41636 20590
rect 41692 20580 41748 21532
rect 41804 21698 41860 21710
rect 41804 21646 41806 21698
rect 41858 21646 41860 21698
rect 41804 21028 41860 21646
rect 43036 21700 43092 21710
rect 43036 21606 43092 21644
rect 43372 21698 43428 21710
rect 43708 21700 43764 21710
rect 43372 21646 43374 21698
rect 43426 21646 43428 21698
rect 42252 21588 42308 21598
rect 42252 21494 42308 21532
rect 42700 21586 42756 21598
rect 42700 21534 42702 21586
rect 42754 21534 42756 21586
rect 42700 21364 42756 21534
rect 42700 21298 42756 21308
rect 41804 20962 41860 20972
rect 43036 21028 43092 21038
rect 43036 20934 43092 20972
rect 43372 20916 43428 21646
rect 43372 20850 43428 20860
rect 43596 21698 43764 21700
rect 43596 21646 43710 21698
rect 43762 21646 43764 21698
rect 43596 21644 43764 21646
rect 41636 20524 41748 20580
rect 43484 20578 43540 20590
rect 43484 20526 43486 20578
rect 43538 20526 43540 20578
rect 41020 18946 41076 18956
rect 41020 18564 41076 18574
rect 41020 17890 41076 18508
rect 41244 18564 41300 18574
rect 41356 18564 41412 19628
rect 41468 19684 41524 19694
rect 41580 19684 41636 20524
rect 42812 20468 42868 20478
rect 42812 20374 42868 20412
rect 41468 19682 41636 19684
rect 41468 19630 41470 19682
rect 41522 19630 41636 19682
rect 41468 19628 41636 19630
rect 41468 19618 41524 19628
rect 41300 18508 41412 18564
rect 41244 18498 41300 18508
rect 41020 17838 41022 17890
rect 41074 17838 41076 17890
rect 41020 17826 41076 17838
rect 41132 18452 41188 18462
rect 40908 17490 40964 17500
rect 40012 16494 40014 16546
rect 40066 16494 40068 16546
rect 40012 13748 40068 16494
rect 40236 16716 40404 16772
rect 40236 15876 40292 16716
rect 40348 16548 40404 16558
rect 41132 16548 41188 18396
rect 41356 18452 41412 18508
rect 41356 18450 41524 18452
rect 41356 18398 41358 18450
rect 41410 18398 41524 18450
rect 41356 18396 41524 18398
rect 41356 18386 41412 18396
rect 41468 17892 41524 18396
rect 41468 17798 41524 17836
rect 41244 17780 41300 17790
rect 41300 17724 41412 17780
rect 41244 17714 41300 17724
rect 40348 16546 40516 16548
rect 40348 16494 40350 16546
rect 40402 16494 40516 16546
rect 40348 16492 40516 16494
rect 40348 16482 40404 16492
rect 40236 15782 40292 15820
rect 40012 13682 40068 13692
rect 39788 13470 39790 13522
rect 39842 13470 39844 13522
rect 39788 13458 39844 13470
rect 39452 12574 39454 12626
rect 39506 12574 39508 12626
rect 39452 12562 39508 12574
rect 38668 10836 38724 10846
rect 38444 10612 38500 10622
rect 38332 10556 38444 10612
rect 38444 10546 38500 10556
rect 38668 10498 38724 10780
rect 38892 10610 38948 12348
rect 39228 12514 39284 12526
rect 39228 12462 39230 12514
rect 39282 12462 39284 12514
rect 39228 10836 39284 12462
rect 40460 11730 40516 16492
rect 41132 16454 41188 16492
rect 40684 16436 40740 16446
rect 40684 16342 40740 16380
rect 41244 15876 41300 15886
rect 41244 15782 41300 15820
rect 41244 14532 41300 14542
rect 41356 14532 41412 17724
rect 41580 17668 41636 19628
rect 41804 19684 41860 19694
rect 42028 19684 42084 19694
rect 41860 19682 42084 19684
rect 41860 19630 42030 19682
rect 42082 19630 42084 19682
rect 41860 19628 42084 19630
rect 41804 19618 41860 19628
rect 42028 19618 42084 19628
rect 43484 18564 43540 20526
rect 43596 18786 43652 21644
rect 43708 21634 43764 21644
rect 43708 20692 43764 20702
rect 43820 20692 43876 25452
rect 44268 24052 44324 24062
rect 43932 23940 43988 23950
rect 44268 23940 44324 23996
rect 43932 23938 44324 23940
rect 43932 23886 43934 23938
rect 43986 23886 44324 23938
rect 43932 23884 44324 23886
rect 43932 23874 43988 23884
rect 44268 22818 44324 23884
rect 44380 23940 44436 23950
rect 44380 23846 44436 23884
rect 45052 23938 45108 25678
rect 45276 24836 45332 24846
rect 45276 24742 45332 24780
rect 45052 23886 45054 23938
rect 45106 23886 45108 23938
rect 45052 23874 45108 23886
rect 45612 23940 45668 25788
rect 45724 25842 45780 26796
rect 46284 26514 46340 27020
rect 46284 26462 46286 26514
rect 46338 26462 46340 26514
rect 46284 26450 46340 26462
rect 46396 26852 46452 26862
rect 46844 26852 46900 27918
rect 46956 27860 47012 27870
rect 47180 27860 47236 27870
rect 47012 27858 47236 27860
rect 47012 27806 47182 27858
rect 47234 27806 47236 27858
rect 47012 27804 47236 27806
rect 46956 27794 47012 27804
rect 47180 27794 47236 27804
rect 46396 26850 46900 26852
rect 46396 26798 46398 26850
rect 46450 26798 46900 26850
rect 46396 26796 46900 26798
rect 45724 25790 45726 25842
rect 45778 25790 45780 25842
rect 45724 25778 45780 25790
rect 46060 25732 46116 25742
rect 46060 25638 46116 25676
rect 45724 24836 45780 24846
rect 45724 24742 45780 24780
rect 46396 24836 46452 26796
rect 46844 26738 46900 26796
rect 46844 26686 46846 26738
rect 46898 26686 46900 26738
rect 46844 26674 46900 26686
rect 46508 26402 46564 26414
rect 47292 26404 47348 26414
rect 46508 26350 46510 26402
rect 46562 26350 46564 26402
rect 46508 25842 46564 26350
rect 46508 25790 46510 25842
rect 46562 25790 46564 25842
rect 46508 25778 46564 25790
rect 47180 26402 47348 26404
rect 47180 26350 47294 26402
rect 47346 26350 47348 26402
rect 47180 26348 47348 26350
rect 47180 25842 47236 26348
rect 47292 26338 47348 26348
rect 47180 25790 47182 25842
rect 47234 25790 47236 25842
rect 47180 25778 47236 25790
rect 45612 23874 45668 23884
rect 46060 24052 46116 24062
rect 44268 22766 44270 22818
rect 44322 22766 44324 22818
rect 44268 22754 44324 22766
rect 45724 23828 45780 23838
rect 45724 23658 45780 23772
rect 46060 23826 46116 23996
rect 46060 23774 46062 23826
rect 46114 23774 46116 23826
rect 46060 23762 46116 23774
rect 46396 23826 46452 24780
rect 46396 23774 46398 23826
rect 46450 23774 46452 23826
rect 46396 23762 46452 23774
rect 45724 23606 45726 23658
rect 45778 23606 45780 23658
rect 44940 22484 44996 22494
rect 44940 22390 44996 22428
rect 45724 22036 45780 23606
rect 45500 21980 45780 22036
rect 43708 20690 43876 20692
rect 43708 20638 43710 20690
rect 43762 20638 43876 20690
rect 43708 20636 43876 20638
rect 44044 21698 44100 21710
rect 44044 21646 44046 21698
rect 44098 21646 44100 21698
rect 43708 20468 43764 20636
rect 44044 20578 44100 21646
rect 44044 20526 44046 20578
rect 44098 20526 44100 20578
rect 44044 20514 44100 20526
rect 44604 21698 44660 21710
rect 44604 21646 44606 21698
rect 44658 21646 44660 21698
rect 43708 20402 43764 20412
rect 43596 18734 43598 18786
rect 43650 18734 43652 18786
rect 43596 18722 43652 18734
rect 44492 19682 44548 19694
rect 44492 19630 44494 19682
rect 44546 19630 44548 19682
rect 43484 18498 43540 18508
rect 42252 18004 42308 18014
rect 42140 17892 42196 17902
rect 41692 17668 41748 17678
rect 41580 17612 41692 17668
rect 41244 14530 41412 14532
rect 41244 14478 41246 14530
rect 41298 14478 41412 14530
rect 41244 14476 41412 14478
rect 41692 15538 41748 17612
rect 41916 17666 41972 17678
rect 41916 17614 41918 17666
rect 41970 17614 41972 17666
rect 41916 17556 41972 17614
rect 41916 17490 41972 17500
rect 41804 16548 41860 16558
rect 41804 16546 41972 16548
rect 41804 16494 41806 16546
rect 41858 16494 41972 16546
rect 41804 16492 41972 16494
rect 41804 16482 41860 16492
rect 41692 15486 41694 15538
rect 41746 15486 41748 15538
rect 41692 14532 41748 15486
rect 41916 14868 41972 16492
rect 42140 15874 42196 17836
rect 42252 17780 42308 17948
rect 43260 17892 43316 17902
rect 44492 17892 44548 19630
rect 43316 17836 43428 17892
rect 43260 17826 43316 17836
rect 42252 17686 42308 17724
rect 43372 17778 43428 17836
rect 44492 17826 44548 17836
rect 43372 17726 43374 17778
rect 43426 17726 43428 17778
rect 43372 17714 43428 17726
rect 43708 17780 43764 17790
rect 42700 17668 42756 17678
rect 42700 17574 42756 17612
rect 42140 15822 42142 15874
rect 42194 15822 42196 15874
rect 42140 15810 42196 15822
rect 42476 16434 42532 16446
rect 42476 16382 42478 16434
rect 42530 16382 42532 16434
rect 42252 14868 42308 14878
rect 41916 14866 42308 14868
rect 41916 14814 42254 14866
rect 42306 14814 42308 14866
rect 41916 14812 42308 14814
rect 42252 14802 42308 14812
rect 41244 14466 41300 14476
rect 41132 13746 41188 13758
rect 41132 13694 41134 13746
rect 41186 13694 41188 13746
rect 41132 13636 41188 13694
rect 41132 13570 41188 13580
rect 41692 13634 41748 14476
rect 41692 13582 41694 13634
rect 41746 13582 41748 13634
rect 41692 13570 41748 13582
rect 42476 12852 42532 16382
rect 43484 14644 43540 14654
rect 43484 13636 43540 14588
rect 42588 12852 42644 12862
rect 42476 12850 42644 12852
rect 42476 12798 42590 12850
rect 42642 12798 42644 12850
rect 42476 12796 42644 12798
rect 42588 12786 42644 12796
rect 40460 11678 40462 11730
rect 40514 11678 40516 11730
rect 40460 11666 40516 11678
rect 42364 11730 42420 11742
rect 42364 11678 42366 11730
rect 42418 11678 42420 11730
rect 41468 11620 41524 11630
rect 42028 11620 42084 11630
rect 41468 11618 42084 11620
rect 41468 11566 41470 11618
rect 41522 11566 42030 11618
rect 42082 11566 42084 11618
rect 41468 11564 42084 11566
rect 41468 11554 41524 11564
rect 39228 10770 39284 10780
rect 41020 11506 41076 11518
rect 41020 11454 41022 11506
rect 41074 11454 41076 11506
rect 41020 10836 41076 11454
rect 41020 10770 41076 10780
rect 41580 10836 41636 10846
rect 41580 10722 41636 10780
rect 41580 10670 41582 10722
rect 41634 10670 41636 10722
rect 41580 10658 41636 10670
rect 42028 10724 42084 11564
rect 42364 10836 42420 11678
rect 42364 10770 42420 10780
rect 42028 10630 42084 10668
rect 43484 10724 43540 13580
rect 43708 13634 43764 17724
rect 44604 16548 44660 21646
rect 45164 21698 45220 21710
rect 45164 21646 45166 21698
rect 45218 21646 45220 21698
rect 45052 20692 45108 20702
rect 45052 20598 45108 20636
rect 45164 20188 45220 21646
rect 45500 20914 45556 21980
rect 45500 20862 45502 20914
rect 45554 20862 45556 20914
rect 45500 20802 45556 20862
rect 45500 20750 45502 20802
rect 45554 20750 45556 20802
rect 45500 20738 45556 20750
rect 45836 21810 45892 21822
rect 45836 21758 45838 21810
rect 45890 21758 45892 21810
rect 45164 20132 45556 20188
rect 45500 19906 45556 20132
rect 45500 19854 45502 19906
rect 45554 19854 45556 19906
rect 45500 19842 45556 19854
rect 45724 19346 45780 19358
rect 45724 19294 45726 19346
rect 45778 19294 45780 19346
rect 45612 18564 45668 18574
rect 45724 18564 45780 19294
rect 45612 18562 45780 18564
rect 45612 18510 45614 18562
rect 45666 18510 45780 18562
rect 45612 18508 45780 18510
rect 45612 17556 45668 18508
rect 45836 17892 45892 21758
rect 46508 21700 46564 21710
rect 46508 20916 46564 21644
rect 47404 21364 47460 29708
rect 47516 28418 47572 29822
rect 48076 28868 48132 28878
rect 47628 28756 47684 28766
rect 47628 28754 47796 28756
rect 47628 28702 47630 28754
rect 47682 28702 47796 28754
rect 47628 28700 47796 28702
rect 47628 28690 47684 28700
rect 47740 28644 47796 28700
rect 48076 28754 48132 28812
rect 48076 28702 48078 28754
rect 48130 28702 48132 28754
rect 48076 28690 48132 28702
rect 47740 28578 47796 28588
rect 47516 28366 47518 28418
rect 47570 28366 47572 28418
rect 47516 28354 47572 28366
rect 48188 27858 48244 30492
rect 48748 30212 48804 30606
rect 48972 30660 49028 32620
rect 49756 32610 49812 32620
rect 49308 32452 49364 32462
rect 49308 32358 49364 32396
rect 49868 31890 49924 33404
rect 50204 32564 50260 32574
rect 50204 32470 50260 32508
rect 49868 31838 49870 31890
rect 49922 31838 49924 31890
rect 49868 31826 49924 31838
rect 49084 31778 49140 31790
rect 49084 31726 49086 31778
rect 49138 31726 49140 31778
rect 49084 30996 49140 31726
rect 50092 31780 50148 31790
rect 50148 31724 50260 31780
rect 50092 31686 50148 31724
rect 49084 30930 49140 30940
rect 49420 31442 49476 31454
rect 49420 31390 49422 31442
rect 49474 31390 49476 31442
rect 48972 30594 49028 30604
rect 49420 30324 49476 31390
rect 50204 30882 50260 31724
rect 50316 31556 50372 34524
rect 50428 33460 50484 38444
rect 50652 38434 50708 38444
rect 51772 38500 51828 38668
rect 52108 38630 52164 38668
rect 52556 39170 52612 39182
rect 52556 39118 52558 39170
rect 52610 39118 52612 39170
rect 50556 38332 50820 38342
rect 50612 38276 50660 38332
rect 50716 38276 50764 38332
rect 50556 38266 50820 38276
rect 51548 37828 51604 37838
rect 51548 37734 51604 37772
rect 51772 36932 51828 38444
rect 52220 37826 52276 37838
rect 52220 37774 52222 37826
rect 52274 37774 52276 37826
rect 52220 37154 52276 37774
rect 52220 37102 52222 37154
rect 52274 37102 52276 37154
rect 52220 37090 52276 37102
rect 52556 37826 52612 39118
rect 52780 38948 52836 38958
rect 53116 38948 53172 42812
rect 53228 42802 53284 42812
rect 53452 42866 53508 42878
rect 53452 42814 53454 42866
rect 53506 42814 53508 42866
rect 53340 42642 53396 42654
rect 53340 42590 53342 42642
rect 53394 42590 53396 42642
rect 53340 40850 53396 42590
rect 53452 42644 53508 42814
rect 53452 42578 53508 42588
rect 53676 42196 53732 44606
rect 54012 43988 54068 45838
rect 54124 45444 54180 46622
rect 54908 46004 54964 46014
rect 55356 46004 55412 46014
rect 54964 45948 55076 46004
rect 54908 45910 54964 45948
rect 54124 44770 54180 45388
rect 54796 44884 54852 44894
rect 54796 44790 54852 44828
rect 54124 44718 54126 44770
rect 54178 44718 54180 44770
rect 54124 44706 54180 44718
rect 54012 43708 54068 43932
rect 54684 43988 54740 43998
rect 54684 43894 54740 43932
rect 55020 43874 55076 45948
rect 55356 45910 55412 45948
rect 55468 44658 55524 44670
rect 55468 44606 55470 44658
rect 55522 44606 55524 44658
rect 55468 44098 55524 44606
rect 55468 44046 55470 44098
rect 55522 44046 55524 44098
rect 55468 44034 55524 44046
rect 56700 43988 56756 43998
rect 56700 43894 56756 43932
rect 57148 43988 57204 43998
rect 57148 43894 57204 43932
rect 55020 43822 55022 43874
rect 55074 43822 55076 43874
rect 54012 43652 54404 43708
rect 54348 42878 54404 43652
rect 53676 42130 53732 42140
rect 53788 42866 53844 42878
rect 53788 42814 53790 42866
rect 53842 42814 53844 42866
rect 53340 40798 53342 40850
rect 53394 40798 53396 40850
rect 53340 40786 53396 40798
rect 53564 41972 53620 41982
rect 53564 40068 53620 41916
rect 53788 41970 53844 42814
rect 54346 42868 54404 42878
rect 54460 42868 54516 42878
rect 54346 42866 54460 42868
rect 54346 42814 54348 42866
rect 54400 42814 54460 42866
rect 54346 42812 54460 42814
rect 54346 42802 54404 42812
rect 54460 42802 54516 42812
rect 54236 42756 54292 42766
rect 54236 42662 54292 42700
rect 54348 42084 54404 42802
rect 55020 42756 55076 43822
rect 55132 42978 55188 42990
rect 55132 42926 55134 42978
rect 55186 42926 55188 42978
rect 55132 42868 55188 42926
rect 56140 42980 56196 42990
rect 55188 42812 55300 42868
rect 55132 42802 55188 42812
rect 55020 42690 55076 42700
rect 55020 42532 55076 42542
rect 54348 42018 54404 42028
rect 54908 42530 55076 42532
rect 54908 42478 55022 42530
rect 55074 42478 55076 42530
rect 54908 42476 55076 42478
rect 53788 41918 53790 41970
rect 53842 41918 53844 41970
rect 53788 41636 53844 41918
rect 53676 40628 53732 40638
rect 53676 40534 53732 40572
rect 53564 40012 53732 40068
rect 53228 39842 53284 39854
rect 53564 39844 53620 39854
rect 53228 39790 53230 39842
rect 53282 39790 53284 39842
rect 53228 39170 53284 39790
rect 53228 39118 53230 39170
rect 53282 39118 53284 39170
rect 53228 39106 53284 39118
rect 53452 39842 53620 39844
rect 53452 39790 53566 39842
rect 53618 39790 53620 39842
rect 53452 39788 53620 39790
rect 53452 39058 53508 39788
rect 53564 39778 53620 39788
rect 53452 39006 53454 39058
rect 53506 39006 53508 39058
rect 53452 38994 53508 39006
rect 53228 38948 53284 38958
rect 53116 38946 53284 38948
rect 53116 38894 53230 38946
rect 53282 38894 53284 38946
rect 53116 38892 53284 38894
rect 52780 38854 52836 38892
rect 53228 38882 53284 38892
rect 53564 38948 53620 38958
rect 53676 38948 53732 40012
rect 53564 38946 53732 38948
rect 53564 38894 53566 38946
rect 53618 38894 53732 38946
rect 53564 38892 53732 38894
rect 53564 38882 53620 38892
rect 52556 37774 52558 37826
rect 52610 37774 52612 37826
rect 50988 36876 51828 36932
rect 50652 36708 50708 36718
rect 50876 36708 50932 36718
rect 50652 36706 50876 36708
rect 50652 36654 50654 36706
rect 50706 36654 50876 36706
rect 50652 36652 50876 36654
rect 50652 36642 50708 36652
rect 50876 36372 50932 36652
rect 50988 36484 51044 36876
rect 51772 36818 51828 36876
rect 51772 36766 51774 36818
rect 51826 36766 51828 36818
rect 51772 36754 51828 36766
rect 51100 36708 51156 36718
rect 51324 36708 51380 36718
rect 51100 36706 51268 36708
rect 51100 36654 51102 36706
rect 51154 36654 51268 36706
rect 51100 36652 51268 36654
rect 51100 36642 51156 36652
rect 51212 36596 51268 36652
rect 51324 36706 51492 36708
rect 51324 36654 51326 36706
rect 51378 36654 51492 36706
rect 51324 36652 51492 36654
rect 51324 36642 51380 36652
rect 51212 36530 51268 36540
rect 50988 36428 51156 36484
rect 50556 36316 50820 36326
rect 50876 36316 51044 36372
rect 50612 36260 50660 36316
rect 50716 36260 50764 36316
rect 50556 36250 50820 36260
rect 50652 35810 50708 35822
rect 50652 35758 50654 35810
rect 50706 35758 50708 35810
rect 50652 34804 50708 35758
rect 50764 35138 50820 35150
rect 50764 35086 50766 35138
rect 50818 35086 50820 35138
rect 50764 34914 50820 35086
rect 50764 34862 50766 34914
rect 50818 34862 50820 34914
rect 50764 34850 50820 34862
rect 50652 34468 50708 34748
rect 50652 34412 50932 34468
rect 50556 34300 50820 34310
rect 50612 34244 50660 34300
rect 50716 34244 50764 34300
rect 50556 34234 50820 34244
rect 50876 34132 50932 34412
rect 50652 34076 50932 34132
rect 50652 34018 50708 34076
rect 50652 33966 50654 34018
rect 50706 33966 50708 34018
rect 50652 33954 50708 33966
rect 50652 33460 50708 33470
rect 50428 33458 50708 33460
rect 50428 33406 50654 33458
rect 50706 33406 50708 33458
rect 50428 33404 50708 33406
rect 50652 32898 50708 33404
rect 50652 32846 50654 32898
rect 50706 32846 50708 32898
rect 50652 32834 50708 32846
rect 50988 32676 51044 36316
rect 51100 35810 51156 36428
rect 51436 36372 51492 36652
rect 51100 35758 51102 35810
rect 51154 35758 51156 35810
rect 51100 35138 51156 35758
rect 51100 35086 51102 35138
rect 51154 35086 51156 35138
rect 51100 34916 51156 35086
rect 51324 36316 51492 36372
rect 51212 34916 51268 34926
rect 51100 34860 51212 34916
rect 51100 34130 51156 34860
rect 51212 34822 51268 34860
rect 51324 34804 51380 36316
rect 52108 35812 52164 35822
rect 52332 35812 52388 35822
rect 52108 35810 52388 35812
rect 52108 35758 52110 35810
rect 52162 35758 52334 35810
rect 52386 35758 52388 35810
rect 52108 35756 52388 35758
rect 52108 35746 52164 35756
rect 52332 35746 52388 35756
rect 51324 34738 51380 34748
rect 51436 35700 51492 35710
rect 51100 34078 51102 34130
rect 51154 34078 51156 34130
rect 51100 34018 51156 34078
rect 51100 33966 51102 34018
rect 51154 33966 51156 34018
rect 51100 33954 51156 33966
rect 51436 34020 51492 35644
rect 51884 35252 51940 35262
rect 51772 35196 51884 35252
rect 51548 34692 51604 34702
rect 51548 34598 51604 34636
rect 51548 34020 51604 34030
rect 51436 33964 51548 34020
rect 51548 33926 51604 33964
rect 51548 33458 51604 33470
rect 51548 33406 51550 33458
rect 51602 33406 51604 33458
rect 50876 32450 50932 32462
rect 50876 32398 50878 32450
rect 50930 32398 50932 32450
rect 50556 32284 50820 32294
rect 50612 32228 50660 32284
rect 50716 32228 50764 32284
rect 50556 32218 50820 32228
rect 50876 31948 50932 32398
rect 50428 31892 50932 31948
rect 50988 32452 51044 32620
rect 51324 32676 51380 32686
rect 51324 32674 51492 32676
rect 51324 32622 51326 32674
rect 51378 32622 51492 32674
rect 51324 32620 51492 32622
rect 51324 32610 51380 32620
rect 50428 31890 50484 31892
rect 50428 31838 50430 31890
rect 50482 31838 50484 31890
rect 50428 31826 50484 31838
rect 50316 31490 50372 31500
rect 50204 30830 50206 30882
rect 50258 30830 50260 30882
rect 50204 30818 50260 30830
rect 50988 30770 51044 32396
rect 50988 30718 50990 30770
rect 51042 30718 51044 30770
rect 50988 30706 51044 30718
rect 51100 32564 51156 32574
rect 51100 31948 51156 32508
rect 51100 31892 51380 31948
rect 49420 30258 49476 30268
rect 49756 30658 49812 30670
rect 49756 30606 49758 30658
rect 49810 30606 49812 30658
rect 48748 30146 48804 30156
rect 48860 29650 48916 29662
rect 48860 29598 48862 29650
rect 48914 29598 48916 29650
rect 48300 28756 48356 28766
rect 48300 28662 48356 28700
rect 48860 28644 48916 29598
rect 49756 29652 49812 30606
rect 50652 30436 50708 30474
rect 50652 30370 50708 30380
rect 50556 30268 50820 30278
rect 50316 30212 50372 30222
rect 50612 30212 50660 30268
rect 50716 30212 50764 30268
rect 50556 30202 50820 30212
rect 50316 29988 50372 30156
rect 50316 29986 50484 29988
rect 50316 29934 50318 29986
rect 50370 29934 50484 29986
rect 50316 29932 50484 29934
rect 50316 29922 50372 29932
rect 49868 29652 49924 29662
rect 49756 29650 49924 29652
rect 49756 29598 49870 29650
rect 49922 29598 49924 29650
rect 49756 29596 49924 29598
rect 49756 28756 49812 29596
rect 49868 29538 49924 29596
rect 49868 29486 49870 29538
rect 49922 29486 49924 29538
rect 49868 29474 49924 29486
rect 49756 28690 49812 28700
rect 50204 28868 50260 28878
rect 48972 28644 49028 28654
rect 48860 28588 48972 28644
rect 48972 28530 49028 28588
rect 48972 28478 48974 28530
rect 49026 28478 49028 28530
rect 48860 28082 48916 28094
rect 48860 28030 48862 28082
rect 48914 28030 48916 28082
rect 48860 27970 48916 28030
rect 48860 27918 48862 27970
rect 48914 27918 48916 27970
rect 48860 27906 48916 27918
rect 48188 27806 48190 27858
rect 48242 27806 48244 27858
rect 47852 27522 47908 27534
rect 47852 27470 47854 27522
rect 47906 27470 47908 27522
rect 47852 26516 47908 27470
rect 48188 26852 48244 27806
rect 48188 26786 48244 26796
rect 48524 27524 48580 27534
rect 47852 26450 47908 26460
rect 47628 25844 47684 25854
rect 47628 23938 47684 25788
rect 47852 25842 47908 25854
rect 47852 25790 47854 25842
rect 47906 25790 47908 25842
rect 47852 24834 47908 25790
rect 47852 24782 47854 24834
rect 47906 24782 47908 24834
rect 47852 24770 47908 24782
rect 48076 25732 48132 25742
rect 47628 23886 47630 23938
rect 47682 23886 47684 23938
rect 47628 23874 47684 23886
rect 48076 23938 48132 25676
rect 48076 23886 48078 23938
rect 48130 23886 48132 23938
rect 48076 23874 48132 23886
rect 47740 21700 47796 21710
rect 48412 21700 48468 21710
rect 47740 21606 47796 21644
rect 48300 21644 48412 21700
rect 48188 21588 48244 21598
rect 47404 21298 47460 21308
rect 48076 21586 48244 21588
rect 48076 21534 48190 21586
rect 48242 21534 48244 21586
rect 48076 21532 48244 21534
rect 45948 20860 46564 20916
rect 45948 20802 46004 20860
rect 45948 20750 45950 20802
rect 46002 20750 46004 20802
rect 45948 19684 46004 20750
rect 46172 20692 46228 20702
rect 46172 20578 46228 20636
rect 46508 20690 46564 20860
rect 46508 20638 46510 20690
rect 46562 20638 46564 20690
rect 46508 20626 46564 20638
rect 46732 20804 46788 20814
rect 46732 20690 46788 20748
rect 47628 20804 47684 20814
rect 47628 20710 47684 20748
rect 46732 20638 46734 20690
rect 46786 20638 46788 20690
rect 46732 20626 46788 20638
rect 48076 20692 48132 21532
rect 48188 21522 48244 21532
rect 48076 20626 48132 20636
rect 48188 21364 48244 21374
rect 46172 20526 46174 20578
rect 46226 20526 46228 20578
rect 46172 20188 46228 20526
rect 47180 20354 47236 20366
rect 47180 20302 47182 20354
rect 47234 20302 47236 20354
rect 47180 20188 47236 20302
rect 46172 20132 46452 20188
rect 46172 19684 46228 19694
rect 45948 19682 46228 19684
rect 45948 19630 46174 19682
rect 46226 19630 46228 19682
rect 45948 19628 46228 19630
rect 46172 19346 46228 19628
rect 46172 19294 46174 19346
rect 46226 19294 46228 19346
rect 46172 19282 46228 19294
rect 46396 19682 46452 20132
rect 46396 19630 46398 19682
rect 46450 19630 46452 19682
rect 46060 18788 46116 18798
rect 46396 18788 46452 19630
rect 46060 18786 46452 18788
rect 46060 18734 46062 18786
rect 46114 18734 46452 18786
rect 46060 18732 46452 18734
rect 46956 20132 47236 20188
rect 48188 20188 48244 21308
rect 48300 20690 48356 21644
rect 48412 21634 48468 21644
rect 48300 20638 48302 20690
rect 48354 20638 48356 20690
rect 48300 20626 48356 20638
rect 48412 20804 48468 20814
rect 48412 20578 48468 20748
rect 48412 20526 48414 20578
rect 48466 20526 48468 20578
rect 48412 20514 48468 20526
rect 48188 20132 48356 20188
rect 46060 18722 46116 18732
rect 46956 18674 47012 20132
rect 48300 19796 48356 20132
rect 48524 19908 48580 27468
rect 48972 27522 49028 28478
rect 49308 28532 49364 28542
rect 49308 27972 49364 28476
rect 48972 27470 48974 27522
rect 49026 27470 49028 27522
rect 48972 27458 49028 27470
rect 49084 27970 49364 27972
rect 49084 27918 49310 27970
rect 49362 27918 49364 27970
rect 49084 27916 49364 27918
rect 48636 26516 48692 26526
rect 48692 26460 48804 26516
rect 48636 26450 48692 26460
rect 48748 21812 48804 26460
rect 49084 25732 49140 27916
rect 49308 27906 49364 27916
rect 50092 28530 50148 28542
rect 50092 28478 50094 28530
rect 50146 28478 50148 28530
rect 50092 28418 50148 28478
rect 50092 28366 50094 28418
rect 50146 28366 50148 28418
rect 49756 27636 49812 27646
rect 49756 27634 49924 27636
rect 49756 27582 49758 27634
rect 49810 27582 49924 27634
rect 49756 27580 49924 27582
rect 49756 27570 49812 27580
rect 49868 27522 49924 27580
rect 49868 27470 49870 27522
rect 49922 27470 49924 27522
rect 49756 26740 49812 26750
rect 49756 26646 49812 26684
rect 49868 26516 49924 27470
rect 50092 27522 50148 28366
rect 50204 28082 50260 28812
rect 50204 28030 50206 28082
rect 50258 28030 50260 28082
rect 50204 27972 50260 28030
rect 50428 28084 50484 29932
rect 50764 29652 50820 29662
rect 50764 29650 50932 29652
rect 50764 29598 50766 29650
rect 50818 29598 50932 29650
rect 50764 29596 50932 29598
rect 50764 29586 50820 29596
rect 50876 29538 50932 29596
rect 50876 29486 50878 29538
rect 50930 29486 50932 29538
rect 50540 28868 50596 28878
rect 50540 28774 50596 28812
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50428 28028 50708 28084
rect 50204 27970 50372 27972
rect 50204 27918 50206 27970
rect 50258 27918 50372 27970
rect 50204 27916 50372 27918
rect 50204 27906 50260 27916
rect 50092 27470 50094 27522
rect 50146 27470 50148 27522
rect 50092 27458 50148 27470
rect 50204 26516 50260 26526
rect 49868 26514 50260 26516
rect 49868 26462 50206 26514
rect 50258 26462 50260 26514
rect 49868 26460 50260 26462
rect 49644 26402 49700 26414
rect 49644 26350 49646 26402
rect 49698 26350 49700 26402
rect 49644 25844 49700 26350
rect 49644 25750 49700 25788
rect 49084 25638 49140 25676
rect 50204 25732 50260 26460
rect 49532 24722 49588 24734
rect 49532 24670 49534 24722
rect 49586 24670 49588 24722
rect 48860 23828 48916 23838
rect 48860 23734 48916 23772
rect 49420 23828 49476 23838
rect 49420 22820 49476 23772
rect 49532 23716 49588 24670
rect 49532 23622 49588 23660
rect 49980 24052 50036 24062
rect 49980 23938 50036 23996
rect 49980 23886 49982 23938
rect 50034 23886 50036 23938
rect 49532 22820 49588 22830
rect 49980 22820 50036 23886
rect 50204 23716 50260 25676
rect 50316 24836 50372 27916
rect 50428 26740 50484 28028
rect 50652 27972 50708 28028
rect 50652 27878 50708 27916
rect 50876 27860 50932 29486
rect 50988 29426 51044 29438
rect 50988 29374 50990 29426
rect 51042 29374 51044 29426
rect 50988 28530 51044 29374
rect 50988 28478 50990 28530
rect 51042 28478 51044 28530
rect 50988 28418 51044 28478
rect 50988 28366 50990 28418
rect 51042 28366 51044 28418
rect 50988 28354 51044 28366
rect 51100 28084 51156 31892
rect 51324 31778 51380 31892
rect 51324 31726 51326 31778
rect 51378 31726 51380 31778
rect 51324 31714 51380 31726
rect 51436 31780 51492 32620
rect 51436 31714 51492 31724
rect 51548 31892 51604 33406
rect 51772 32674 51828 35196
rect 51884 35186 51940 35196
rect 51884 35028 51940 35038
rect 51884 34934 51940 34972
rect 52556 35028 52612 37774
rect 52892 37828 52948 37838
rect 53228 37828 53284 37838
rect 52892 37734 52948 37772
rect 53004 37826 53284 37828
rect 53004 37774 53230 37826
rect 53282 37774 53284 37826
rect 53004 37772 53284 37774
rect 52780 36708 52836 36718
rect 52780 36614 52836 36652
rect 52892 35810 52948 35822
rect 52892 35758 52894 35810
rect 52946 35758 52948 35810
rect 52892 35698 52948 35758
rect 52892 35646 52894 35698
rect 52946 35646 52948 35698
rect 52892 35634 52948 35646
rect 53004 35252 53060 37772
rect 53228 37762 53284 37772
rect 53116 36932 53172 36942
rect 53116 36838 53172 36876
rect 53676 36708 53732 38892
rect 53788 38946 53844 41580
rect 54796 41970 54852 41982
rect 54796 41918 54798 41970
rect 54850 41918 54852 41970
rect 54796 41636 54852 41918
rect 54796 41570 54852 41580
rect 54796 40852 54852 40862
rect 54908 40852 54964 42476
rect 55020 42466 55076 42476
rect 55244 42084 55300 42812
rect 55356 42866 55412 42878
rect 55356 42814 55358 42866
rect 55410 42814 55412 42866
rect 55356 42756 55412 42814
rect 56028 42868 56084 42878
rect 55356 42690 55412 42700
rect 55692 42756 55748 42766
rect 55692 42662 55748 42700
rect 55804 42642 55860 42654
rect 55804 42590 55806 42642
rect 55858 42590 55860 42642
rect 55804 42532 55860 42590
rect 55244 42028 55412 42084
rect 55356 41972 55412 42028
rect 55692 41972 55748 41982
rect 55356 41970 55748 41972
rect 55356 41918 55694 41970
rect 55746 41918 55748 41970
rect 55356 41916 55748 41918
rect 54796 40850 54964 40852
rect 54796 40798 54798 40850
rect 54850 40798 54964 40850
rect 54796 40796 54964 40798
rect 55468 41634 55524 41646
rect 55468 41582 55470 41634
rect 55522 41582 55524 41634
rect 54796 40786 54852 40796
rect 54236 40738 54292 40750
rect 54236 40686 54238 40738
rect 54290 40686 54292 40738
rect 53900 40068 53956 40078
rect 53900 39974 53956 40012
rect 54236 39956 54292 40686
rect 55468 40738 55524 41582
rect 55692 41188 55748 41916
rect 55804 41636 55860 42476
rect 56028 41860 56084 42812
rect 56140 42866 56196 42924
rect 56140 42814 56142 42866
rect 56194 42814 56196 42866
rect 56140 42644 56196 42814
rect 56476 42868 56532 42878
rect 56476 42774 56532 42812
rect 56924 42756 56980 42766
rect 56924 42662 56980 42700
rect 56140 42578 56196 42588
rect 57372 42644 57428 42654
rect 56700 42532 56756 42542
rect 56700 42082 56756 42476
rect 56700 42030 56702 42082
rect 56754 42030 56756 42082
rect 56700 42018 56756 42030
rect 57372 42084 57428 42588
rect 57820 42642 57876 42654
rect 57820 42590 57822 42642
rect 57874 42590 57876 42642
rect 57820 42530 57876 42590
rect 57820 42478 57822 42530
rect 57874 42478 57876 42530
rect 57820 42466 57876 42478
rect 57372 42028 57764 42084
rect 56028 41858 56196 41860
rect 56028 41806 56030 41858
rect 56082 41806 56196 41858
rect 56028 41804 56196 41806
rect 56028 41794 56084 41804
rect 55804 41570 55860 41580
rect 56140 41748 56196 41804
rect 55916 41188 55972 41198
rect 55692 41186 55972 41188
rect 55692 41134 55918 41186
rect 55970 41134 55972 41186
rect 55692 41132 55972 41134
rect 55916 41122 55972 41132
rect 55468 40686 55470 40738
rect 55522 40686 55524 40738
rect 55468 40674 55524 40686
rect 54348 39956 54404 39966
rect 53788 38894 53790 38946
rect 53842 38894 53844 38946
rect 53788 38882 53844 38894
rect 54012 39954 54404 39956
rect 54012 39902 54350 39954
rect 54402 39902 54404 39954
rect 54012 39900 54404 39902
rect 53788 38724 53844 38734
rect 53788 38630 53844 38668
rect 54012 38164 54068 39900
rect 54348 39890 54404 39900
rect 55692 39954 55748 39966
rect 55692 39902 55694 39954
rect 55746 39902 55748 39954
rect 55020 39844 55076 39854
rect 55020 39842 55412 39844
rect 55020 39790 55022 39842
rect 55074 39790 55412 39842
rect 55020 39788 55412 39790
rect 55020 39778 55076 39788
rect 55356 39058 55412 39788
rect 55692 39172 55748 39902
rect 55804 39172 55860 39182
rect 55692 39170 55860 39172
rect 55692 39118 55806 39170
rect 55858 39118 55860 39170
rect 55692 39116 55860 39118
rect 55804 39106 55860 39116
rect 55356 39006 55358 39058
rect 55410 39006 55412 39058
rect 55356 38994 55412 39006
rect 54124 38946 54180 38958
rect 54124 38894 54126 38946
rect 54178 38894 54180 38946
rect 54124 38836 54180 38894
rect 55580 38948 55636 38958
rect 54236 38836 54292 38846
rect 54124 38834 54292 38836
rect 54124 38782 54238 38834
rect 54290 38782 54292 38834
rect 54124 38780 54292 38782
rect 54236 38770 54292 38780
rect 55580 38836 55636 38892
rect 55580 38834 55860 38836
rect 55580 38782 55582 38834
rect 55634 38782 55860 38834
rect 55580 38780 55860 38782
rect 55580 38770 55636 38780
rect 54684 38724 54740 38734
rect 54684 38630 54740 38668
rect 53788 38108 54068 38164
rect 53788 37938 53844 38108
rect 55804 38050 55860 38780
rect 56028 38724 56084 38734
rect 56140 38724 56196 41692
rect 57148 41748 57204 41758
rect 57148 41654 57204 41692
rect 57596 41746 57652 41758
rect 57596 41694 57598 41746
rect 57650 41694 57652 41746
rect 56252 41186 56308 41198
rect 56252 41134 56254 41186
rect 56306 41134 56308 41186
rect 56252 40962 56308 41134
rect 56252 40910 56254 40962
rect 56306 40910 56308 40962
rect 56252 40898 56308 40910
rect 57260 39844 57316 39854
rect 57596 39844 57652 41694
rect 56924 39842 57652 39844
rect 56924 39790 57262 39842
rect 57314 39790 57652 39842
rect 56924 39788 57652 39790
rect 56812 39506 56868 39518
rect 56812 39454 56814 39506
rect 56866 39454 56868 39506
rect 56812 39170 56868 39454
rect 56812 39118 56814 39170
rect 56866 39118 56868 39170
rect 56812 39106 56868 39118
rect 56476 38948 56532 38958
rect 56924 38948 56980 39788
rect 57260 39778 57316 39788
rect 56532 38946 56980 38948
rect 56532 38894 56926 38946
rect 56978 38894 56980 38946
rect 56532 38892 56980 38894
rect 56476 38854 56532 38892
rect 56924 38882 56980 38892
rect 56084 38668 56196 38724
rect 56028 38630 56084 38668
rect 55804 37998 55806 38050
rect 55858 37998 55860 38050
rect 53788 37886 53790 37938
rect 53842 37886 53844 37938
rect 53788 36932 53844 37886
rect 55020 37938 55076 37950
rect 55020 37886 55022 37938
rect 55074 37886 55076 37938
rect 54348 37826 54404 37838
rect 54348 37774 54350 37826
rect 54402 37774 54404 37826
rect 54348 37156 54404 37774
rect 54348 37090 54404 37100
rect 55020 37044 55076 37886
rect 55132 37044 55188 37054
rect 55020 37042 55188 37044
rect 55020 36990 55134 37042
rect 55186 36990 55188 37042
rect 55020 36988 55188 36990
rect 55132 36978 55188 36988
rect 53788 36866 53844 36876
rect 54124 36930 54180 36942
rect 54124 36878 54126 36930
rect 54178 36878 54180 36930
rect 54124 36708 54180 36878
rect 53676 36652 54124 36708
rect 53004 35186 53060 35196
rect 53116 35812 53172 35822
rect 52556 34962 52612 34972
rect 52780 34916 52836 34926
rect 52108 34804 52164 34814
rect 51996 34020 52052 34030
rect 52108 34020 52164 34748
rect 52780 34802 52836 34860
rect 52780 34750 52782 34802
rect 52834 34750 52836 34802
rect 51996 34018 52164 34020
rect 51996 33966 51998 34018
rect 52050 33966 52164 34018
rect 51996 33964 52164 33966
rect 51996 33954 52052 33964
rect 51772 32622 51774 32674
rect 51826 32622 51828 32674
rect 51772 32610 51828 32622
rect 51884 33796 51940 33806
rect 51884 32786 51940 33740
rect 51884 32734 51886 32786
rect 51938 32734 51940 32786
rect 51884 32452 51940 32734
rect 51548 31778 51604 31836
rect 51548 31726 51550 31778
rect 51602 31726 51604 31778
rect 51548 31714 51604 31726
rect 51660 32396 51940 32452
rect 51324 31556 51380 31566
rect 51212 30882 51268 30894
rect 51212 30830 51214 30882
rect 51266 30830 51268 30882
rect 51212 29652 51268 30830
rect 51212 29426 51268 29596
rect 51324 30658 51380 31500
rect 51324 30606 51326 30658
rect 51378 30606 51380 30658
rect 51324 29538 51380 30606
rect 51324 29486 51326 29538
rect 51378 29486 51380 29538
rect 51324 29474 51380 29486
rect 51548 30996 51604 31006
rect 51548 30882 51604 30940
rect 51548 30830 51550 30882
rect 51602 30830 51604 30882
rect 51548 29988 51604 30830
rect 51660 30548 51716 32396
rect 52108 31948 52164 33964
rect 52332 34692 52388 34702
rect 52220 33460 52276 33470
rect 52220 33366 52276 33404
rect 51884 31892 51940 31902
rect 51660 30482 51716 30492
rect 51772 31778 51828 31790
rect 51772 31726 51774 31778
rect 51826 31726 51828 31778
rect 51772 30100 51828 31726
rect 51772 30034 51828 30044
rect 51660 29988 51716 29998
rect 51548 29986 51716 29988
rect 51548 29934 51662 29986
rect 51714 29934 51716 29986
rect 51548 29932 51716 29934
rect 51212 29374 51214 29426
rect 51266 29374 51268 29426
rect 51212 29362 51268 29374
rect 51548 28868 51604 29932
rect 51660 29922 51716 29932
rect 51548 28802 51604 28812
rect 51884 28868 51940 31836
rect 51996 31892 52164 31948
rect 51996 31890 52052 31892
rect 51996 31838 51998 31890
rect 52050 31838 52052 31890
rect 51996 29652 52052 31838
rect 52220 31666 52276 31678
rect 52220 31614 52222 31666
rect 52274 31614 52276 31666
rect 52220 30996 52276 31614
rect 52332 31332 52388 34636
rect 52780 33908 52836 34750
rect 52668 33794 52724 33806
rect 52668 33742 52670 33794
rect 52722 33742 52724 33794
rect 52668 32900 52724 33742
rect 52668 32834 52724 32844
rect 52780 32788 52836 33852
rect 53004 34916 53060 34926
rect 53004 34802 53060 34860
rect 53004 34750 53006 34802
rect 53058 34750 53060 34802
rect 52892 33796 52948 33806
rect 52892 33702 52948 33740
rect 52892 32788 52948 32798
rect 52780 32786 52948 32788
rect 52780 32734 52894 32786
rect 52946 32734 52948 32786
rect 52780 32732 52948 32734
rect 53004 32788 53060 34750
rect 53116 33906 53172 35756
rect 53228 35812 53284 35822
rect 53228 35810 53396 35812
rect 53228 35758 53230 35810
rect 53282 35758 53396 35810
rect 53228 35756 53396 35758
rect 53228 35746 53284 35756
rect 53116 33854 53118 33906
rect 53170 33854 53172 33906
rect 53116 33842 53172 33854
rect 53340 35028 53396 35756
rect 53228 32788 53284 32798
rect 53004 32786 53284 32788
rect 53004 32734 53230 32786
rect 53282 32734 53284 32786
rect 53004 32732 53284 32734
rect 52892 32722 52948 32732
rect 53228 32722 53284 32732
rect 52892 32562 52948 32574
rect 52892 32510 52894 32562
rect 52946 32510 52948 32562
rect 52556 32002 52612 32014
rect 52556 31950 52558 32002
rect 52610 31950 52612 32002
rect 52444 31778 52500 31790
rect 52444 31726 52446 31778
rect 52498 31726 52500 31778
rect 52444 31556 52500 31726
rect 52556 31668 52612 31950
rect 52892 31890 52948 32510
rect 53340 31948 53396 34972
rect 53564 35810 53620 35822
rect 53564 35758 53566 35810
rect 53618 35758 53620 35810
rect 53564 34580 53620 35758
rect 53788 34916 53844 36652
rect 54124 36614 54180 36652
rect 54348 36932 54404 36942
rect 54348 35922 54404 36876
rect 54348 35870 54350 35922
rect 54402 35870 54404 35922
rect 54348 35858 54404 35870
rect 54572 36706 54628 36718
rect 54572 36654 54574 36706
rect 54626 36654 54628 36706
rect 53900 35812 53956 35822
rect 53900 35718 53956 35756
rect 53788 34850 53844 34860
rect 54572 35140 54628 36654
rect 55804 36708 55860 37998
rect 55804 36642 55860 36652
rect 56028 36818 56084 36830
rect 56028 36766 56030 36818
rect 56082 36766 56084 36818
rect 55692 36036 55748 36046
rect 55916 36036 55972 36046
rect 55692 36034 55916 36036
rect 55692 35982 55694 36034
rect 55746 35982 55916 36034
rect 55692 35980 55916 35982
rect 55692 35970 55748 35980
rect 55916 35970 55972 35980
rect 55020 35810 55076 35822
rect 55020 35758 55022 35810
rect 55074 35758 55076 35810
rect 54572 35084 54964 35140
rect 54012 34580 54068 34590
rect 53564 34578 54068 34580
rect 53564 34526 54014 34578
rect 54066 34526 54068 34578
rect 53564 34524 54068 34526
rect 54012 34514 54068 34524
rect 54012 34020 54068 34030
rect 53900 33684 53956 33694
rect 52892 31838 52894 31890
rect 52946 31838 52948 31890
rect 52892 31826 52948 31838
rect 53228 31892 53396 31948
rect 53788 32900 53844 32910
rect 53228 31890 53284 31892
rect 53228 31838 53230 31890
rect 53282 31838 53284 31890
rect 53228 31826 53284 31838
rect 53564 31778 53620 31790
rect 53564 31726 53566 31778
rect 53618 31726 53620 31778
rect 53564 31668 53620 31726
rect 52556 31612 53620 31668
rect 52444 31490 52500 31500
rect 52332 31276 52724 31332
rect 52220 30930 52276 30940
rect 52668 30770 52724 31276
rect 52668 30718 52670 30770
rect 52722 30718 52724 30770
rect 52668 30706 52724 30718
rect 52108 30548 52164 30558
rect 52108 30546 52612 30548
rect 52108 30494 52110 30546
rect 52162 30494 52612 30546
rect 52108 30492 52612 30494
rect 52108 30482 52164 30492
rect 52556 30100 52612 30492
rect 53004 30436 53060 30446
rect 53004 30434 53284 30436
rect 53004 30382 53006 30434
rect 53058 30382 53284 30434
rect 53004 30380 53284 30382
rect 52556 30044 52948 30100
rect 52892 29874 52948 30044
rect 52892 29822 52894 29874
rect 52946 29822 52948 29874
rect 52892 29810 52948 29822
rect 51996 29586 52052 29596
rect 52332 29652 52388 29662
rect 52332 29558 52388 29596
rect 51660 28532 51716 28542
rect 51884 28532 51940 28812
rect 52780 28868 52836 28878
rect 51660 28530 51828 28532
rect 51660 28478 51662 28530
rect 51714 28478 51828 28530
rect 51660 28476 51828 28478
rect 51660 28466 51716 28476
rect 51100 28028 51268 28084
rect 51100 27860 51156 27870
rect 50876 27804 51100 27860
rect 51100 27766 51156 27804
rect 51212 26964 51268 28028
rect 51660 27972 51716 27982
rect 51660 27858 51716 27916
rect 51660 27806 51662 27858
rect 51714 27806 51716 27858
rect 51660 27794 51716 27806
rect 51772 27748 51828 28476
rect 51884 28466 51940 28476
rect 52108 28532 52164 28542
rect 52108 28530 52276 28532
rect 52108 28478 52110 28530
rect 52162 28478 52276 28530
rect 52108 28476 52276 28478
rect 52108 28466 52164 28476
rect 52108 27972 52164 27982
rect 52108 27858 52164 27916
rect 52108 27806 52110 27858
rect 52162 27806 52164 27858
rect 52108 27794 52164 27806
rect 52220 27860 52276 28476
rect 52332 27860 52388 27870
rect 52220 27804 52332 27860
rect 52332 27766 52388 27804
rect 51884 27748 51940 27758
rect 51772 27746 51940 27748
rect 51772 27694 51886 27746
rect 51938 27694 51940 27746
rect 51772 27692 51940 27694
rect 51884 27634 51940 27692
rect 51884 27582 51886 27634
rect 51938 27582 51940 27634
rect 51884 27570 51940 27582
rect 50428 26674 50484 26684
rect 50652 26908 51268 26964
rect 50652 26850 50708 26908
rect 50652 26798 50654 26850
rect 50706 26798 50708 26850
rect 50652 26402 50708 26798
rect 50988 26740 51044 26750
rect 50876 26628 50932 26638
rect 50876 26534 50932 26572
rect 50652 26350 50654 26402
rect 50706 26350 50708 26402
rect 50652 26338 50708 26350
rect 50556 26236 50820 26246
rect 50612 26180 50660 26236
rect 50716 26180 50764 26236
rect 50556 26170 50820 26180
rect 50988 25730 51044 26684
rect 51212 26628 51268 26908
rect 51996 27522 52052 27534
rect 51996 27470 51998 27522
rect 52050 27470 52052 27522
rect 51548 26852 51604 26862
rect 51996 26852 52052 27470
rect 51996 26796 52724 26852
rect 51324 26740 51380 26750
rect 51324 26646 51380 26684
rect 51548 26738 51604 26796
rect 51548 26686 51550 26738
rect 51602 26686 51604 26738
rect 51548 26674 51604 26686
rect 52668 26738 52724 26796
rect 52668 26686 52670 26738
rect 52722 26686 52724 26738
rect 52668 26674 52724 26686
rect 51212 26562 51268 26572
rect 51884 26626 51940 26638
rect 51884 26574 51886 26626
rect 51938 26574 51940 26626
rect 50988 25678 50990 25730
rect 51042 25678 51044 25730
rect 50988 25666 51044 25678
rect 51660 25172 51716 25182
rect 50316 24780 50708 24836
rect 50204 23650 50260 23660
rect 50428 24052 50484 24780
rect 50652 24666 50708 24780
rect 50652 24614 50654 24666
rect 50706 24614 50708 24666
rect 50652 24602 50708 24614
rect 51212 24498 51268 24510
rect 51212 24446 51214 24498
rect 51266 24446 51268 24498
rect 50556 24220 50820 24230
rect 50612 24164 50660 24220
rect 50716 24164 50764 24220
rect 50556 24154 50820 24164
rect 50428 23602 50484 23996
rect 50428 23550 50430 23602
rect 50482 23550 50484 23602
rect 50428 23538 50484 23550
rect 50652 23826 50708 23838
rect 50652 23774 50654 23826
rect 50706 23774 50708 23826
rect 50652 23716 50708 23774
rect 49420 22818 49812 22820
rect 49420 22766 49534 22818
rect 49586 22766 49812 22818
rect 49420 22764 49812 22766
rect 49532 22754 49588 22764
rect 49756 21922 49812 22764
rect 49980 22818 50260 22820
rect 49980 22766 49982 22818
rect 50034 22766 50260 22818
rect 49980 22764 50260 22766
rect 49980 22754 50036 22764
rect 49756 21870 49758 21922
rect 49810 21870 49812 21922
rect 48860 21812 48916 21822
rect 48748 21810 48916 21812
rect 48748 21758 48862 21810
rect 48914 21758 48916 21810
rect 48748 21756 48916 21758
rect 48860 20188 48916 21756
rect 49756 21812 49812 21870
rect 49756 21746 49812 21756
rect 50204 21922 50260 22764
rect 50428 22484 50484 22494
rect 50652 22484 50708 23660
rect 51212 22484 51268 24446
rect 50428 22482 51268 22484
rect 50428 22430 50430 22482
rect 50482 22430 51214 22482
rect 51266 22430 51268 22482
rect 50428 22428 51268 22430
rect 50428 22418 50484 22428
rect 50556 22204 50820 22214
rect 50612 22148 50660 22204
rect 50716 22148 50764 22204
rect 50556 22138 50820 22148
rect 50204 21870 50206 21922
rect 50258 21870 50260 21922
rect 50204 21812 50260 21870
rect 50652 21812 50708 21822
rect 50204 21810 50708 21812
rect 50204 21758 50654 21810
rect 50706 21758 50708 21810
rect 50204 21756 50708 21758
rect 50204 21700 50260 21756
rect 50204 21634 50260 21644
rect 49308 21586 49364 21598
rect 49308 21534 49310 21586
rect 49362 21534 49364 21586
rect 49308 20692 49364 21534
rect 50652 21588 50708 21756
rect 50764 21812 50820 21822
rect 50764 21718 50820 21756
rect 50652 21522 50708 21532
rect 50988 21700 51044 21710
rect 51212 21700 51268 22428
rect 51660 22818 51716 25116
rect 51884 24724 51940 26574
rect 52108 26628 52164 26638
rect 52108 25284 52164 26572
rect 52220 25732 52276 25742
rect 52220 25638 52276 25676
rect 51884 24658 51940 24668
rect 51996 25228 52164 25284
rect 51884 24500 51940 24510
rect 51884 24406 51940 24444
rect 51772 23828 51828 23838
rect 51772 23714 51828 23772
rect 51772 23662 51774 23714
rect 51826 23662 51828 23714
rect 51772 23650 51828 23662
rect 51660 22766 51662 22818
rect 51714 22766 51716 22818
rect 50988 21698 51268 21700
rect 50988 21646 50990 21698
rect 51042 21646 51268 21698
rect 50988 21644 51268 21646
rect 51436 21812 51492 21822
rect 50092 21028 50148 21038
rect 48860 20132 49140 20188
rect 48524 19842 48580 19852
rect 47964 19684 48020 19694
rect 47516 19572 47572 19582
rect 47516 19570 47684 19572
rect 47516 19518 47518 19570
rect 47570 19518 47684 19570
rect 47516 19516 47684 19518
rect 47516 19506 47572 19516
rect 46956 18622 46958 18674
rect 47010 18622 47012 18674
rect 46956 18610 47012 18622
rect 47628 18674 47684 19516
rect 47628 18622 47630 18674
rect 47682 18622 47684 18674
rect 47628 18610 47684 18622
rect 47964 18674 48020 19628
rect 47964 18622 47966 18674
rect 48018 18622 48020 18674
rect 47964 18610 48020 18622
rect 46172 18564 46228 18574
rect 46060 17892 46116 17902
rect 45836 17890 46116 17892
rect 45836 17838 46062 17890
rect 46114 17838 46116 17890
rect 45836 17836 46116 17838
rect 46060 17826 46116 17836
rect 45612 17490 45668 17500
rect 45724 16770 45780 16782
rect 45724 16718 45726 16770
rect 45778 16718 45780 16770
rect 45052 16660 45108 16670
rect 45388 16660 45444 16670
rect 45108 16658 45444 16660
rect 45108 16606 45390 16658
rect 45442 16606 45444 16658
rect 45108 16604 45444 16606
rect 45052 16566 45108 16604
rect 45388 16594 45444 16604
rect 45724 16660 45780 16718
rect 45724 16594 45780 16604
rect 44604 16482 44660 16492
rect 45164 15092 45220 15102
rect 43820 14644 43876 14654
rect 43820 14550 43876 14588
rect 44940 14644 44996 14654
rect 45164 14644 45220 15036
rect 44996 14588 45220 14644
rect 44940 14550 44996 14588
rect 44268 14532 44324 14542
rect 44268 14438 44324 14476
rect 43708 13582 43710 13634
rect 43762 13582 43764 13634
rect 43708 13570 43764 13582
rect 45052 13634 45108 13646
rect 45052 13582 45054 13634
rect 45106 13582 45108 13634
rect 44492 13524 44548 13534
rect 45052 13524 45108 13582
rect 44492 13522 45108 13524
rect 44492 13470 44494 13522
rect 44546 13470 45108 13522
rect 44492 13468 45108 13470
rect 45164 13524 45220 14588
rect 45500 14532 45556 14542
rect 45388 13748 45444 13758
rect 45388 13654 45444 13692
rect 45164 13468 45444 13524
rect 44492 13458 44548 13468
rect 45388 12404 45444 13468
rect 44380 11730 44436 11742
rect 45388 11732 45444 12348
rect 44380 11678 44382 11730
rect 44434 11678 44436 11730
rect 43484 10658 43540 10668
rect 43596 10836 43652 10846
rect 43596 10722 43652 10780
rect 43596 10670 43598 10722
rect 43650 10670 43652 10722
rect 43596 10658 43652 10670
rect 38892 10558 38894 10610
rect 38946 10558 38948 10610
rect 38892 10546 38948 10558
rect 39116 10612 39172 10622
rect 39116 10518 39172 10556
rect 41132 10612 41188 10622
rect 41132 10518 41188 10556
rect 44044 10612 44100 10622
rect 44044 10518 44100 10556
rect 44380 10612 44436 11678
rect 45276 11676 45444 11732
rect 44380 10546 44436 10556
rect 44492 10724 44548 10734
rect 38668 10446 38670 10498
rect 38722 10446 38724 10498
rect 38668 10434 38724 10446
rect 44492 9826 44548 10668
rect 45164 10612 45220 10622
rect 45276 10612 45332 11676
rect 45388 10836 45444 10846
rect 45500 10836 45556 14476
rect 46060 13860 46116 13870
rect 46172 13860 46228 18508
rect 47292 18564 47348 18574
rect 47292 18562 47460 18564
rect 47292 18510 47294 18562
rect 47346 18510 47460 18562
rect 47292 18508 47460 18510
rect 47292 18498 47348 18508
rect 47180 17556 47236 17566
rect 47292 17556 47348 17566
rect 47236 17554 47348 17556
rect 47236 17502 47294 17554
rect 47346 17502 47348 17554
rect 47236 17500 47348 17502
rect 46060 13858 46228 13860
rect 46060 13806 46062 13858
rect 46114 13806 46228 13858
rect 46060 13804 46228 13806
rect 46956 16548 47012 16558
rect 46060 13794 46116 13804
rect 46620 13748 46676 13758
rect 46956 13748 47012 16492
rect 47180 15540 47236 17500
rect 47292 17490 47348 17500
rect 47404 16660 47460 18508
rect 48300 17890 48356 19740
rect 49084 19794 49140 20132
rect 49084 19742 49086 19794
rect 49138 19742 49140 19794
rect 49084 19730 49140 19742
rect 48748 19684 48804 19694
rect 48748 19590 48804 19628
rect 48300 17838 48302 17890
rect 48354 17838 48356 17890
rect 48300 17826 48356 17838
rect 48524 18562 48580 18574
rect 48524 18510 48526 18562
rect 48578 18510 48580 18562
rect 47292 16548 47348 16558
rect 47292 16434 47348 16492
rect 47292 16382 47294 16434
rect 47346 16382 47348 16434
rect 47292 16370 47348 16382
rect 47404 15764 47460 16604
rect 47740 17554 47796 17566
rect 47740 17502 47742 17554
rect 47794 17502 47796 17554
rect 47628 16436 47684 16446
rect 47516 15764 47572 15774
rect 47404 15708 47516 15764
rect 47516 15698 47572 15708
rect 47292 15540 47348 15550
rect 47068 15538 47348 15540
rect 47068 15486 47294 15538
rect 47346 15486 47348 15538
rect 47068 15484 47348 15486
rect 47068 14532 47124 15484
rect 47292 15474 47348 15484
rect 47628 15204 47684 16380
rect 47740 15876 47796 17502
rect 48524 16548 48580 18510
rect 49084 18562 49140 18574
rect 49084 18510 49086 18562
rect 49138 18510 49140 18562
rect 49084 18002 49140 18510
rect 49084 17950 49086 18002
rect 49138 17950 49140 18002
rect 49084 17938 49140 17950
rect 48972 17666 49028 17678
rect 48972 17614 48974 17666
rect 49026 17614 49028 17666
rect 48972 17556 49028 17614
rect 48972 17490 49028 17500
rect 49308 17666 49364 20636
rect 49868 21026 50148 21028
rect 49868 20974 50094 21026
rect 50146 20974 50148 21026
rect 49868 20972 50148 20974
rect 49756 19908 49812 19918
rect 49756 19814 49812 19852
rect 49308 17614 49310 17666
rect 49362 17614 49364 17666
rect 49308 16884 49364 17614
rect 48412 16436 48468 16446
rect 48412 16342 48468 16380
rect 48524 16212 48580 16492
rect 49084 16828 49364 16884
rect 49420 19682 49476 19694
rect 49420 19630 49422 19682
rect 49474 19630 49476 19682
rect 48860 16436 48916 16446
rect 49084 16436 49140 16828
rect 49420 16772 49476 19630
rect 49756 18564 49812 18574
rect 49868 18564 49924 20972
rect 50092 20962 50148 20972
rect 50092 20692 50148 20702
rect 50092 20578 50148 20636
rect 50764 20692 50820 20702
rect 50988 20692 51044 21644
rect 51436 20804 51492 21756
rect 50820 20636 51044 20692
rect 51324 20802 51492 20804
rect 51324 20750 51438 20802
rect 51490 20750 51492 20802
rect 51324 20748 51492 20750
rect 50764 20626 50820 20636
rect 50092 20526 50094 20578
rect 50146 20526 50148 20578
rect 50092 20514 50148 20526
rect 50556 20188 50820 20198
rect 51324 20188 51380 20748
rect 51436 20738 51492 20748
rect 50612 20132 50660 20188
rect 50716 20132 50764 20188
rect 50556 20122 50820 20132
rect 51212 20132 51380 20188
rect 50204 19796 50260 19806
rect 50204 19702 50260 19740
rect 50876 19682 50932 19694
rect 50876 19630 50878 19682
rect 50930 19630 50932 19682
rect 49756 18562 49924 18564
rect 49756 18510 49758 18562
rect 49810 18510 49924 18562
rect 49756 18508 49924 18510
rect 50540 18564 50596 18574
rect 49756 18498 49812 18508
rect 50540 18470 50596 18508
rect 50556 18172 50820 18182
rect 50612 18116 50660 18172
rect 50716 18116 50764 18172
rect 50556 18106 50820 18116
rect 50876 17668 50932 19630
rect 50876 17602 50932 17612
rect 50988 18898 51044 18910
rect 50988 18846 50990 18898
rect 51042 18846 51044 18898
rect 50988 18450 51044 18846
rect 50988 18398 50990 18450
rect 51042 18398 51044 18450
rect 49308 16716 49476 16772
rect 49532 17556 49588 17566
rect 48916 16380 49140 16436
rect 49196 16436 49252 16446
rect 48860 16342 48916 16380
rect 48412 16156 48580 16212
rect 48300 15876 48356 15886
rect 47740 15820 48300 15876
rect 48188 15762 48244 15820
rect 48300 15810 48356 15820
rect 48188 15710 48190 15762
rect 48242 15710 48244 15762
rect 48188 15698 48244 15710
rect 48412 15652 48468 16156
rect 49084 15988 49140 15998
rect 48972 15932 49084 15988
rect 48636 15764 48692 15774
rect 48412 15586 48468 15596
rect 48524 15708 48636 15764
rect 47740 15540 47796 15550
rect 47740 15446 47796 15484
rect 47628 15138 47684 15148
rect 48524 14644 48580 15708
rect 48636 15698 48692 15708
rect 48972 15650 49028 15932
rect 49084 15922 49140 15932
rect 49196 15876 49252 16380
rect 49196 15782 49252 15820
rect 48972 15598 48974 15650
rect 49026 15598 49028 15650
rect 48972 15540 49028 15598
rect 48972 15474 49028 15484
rect 48636 15426 48692 15438
rect 48636 15374 48638 15426
rect 48690 15374 48692 15426
rect 48636 14980 48692 15374
rect 48636 14924 49028 14980
rect 48636 14644 48692 14654
rect 48524 14642 48692 14644
rect 48524 14590 48638 14642
rect 48690 14590 48692 14642
rect 48524 14588 48692 14590
rect 48636 14578 48692 14588
rect 48972 14642 49028 14924
rect 48972 14590 48974 14642
rect 49026 14590 49028 14642
rect 48972 14578 49028 14590
rect 49308 14642 49364 16716
rect 49420 16324 49476 16334
rect 49420 15652 49476 16268
rect 49532 15876 49588 17500
rect 49868 17554 49924 17566
rect 49868 17502 49870 17554
rect 49922 17502 49924 17554
rect 49644 16434 49700 16446
rect 49644 16382 49646 16434
rect 49698 16382 49700 16434
rect 49644 16324 49700 16382
rect 49868 16436 49924 17502
rect 50764 17554 50820 17566
rect 50764 17502 50766 17554
rect 50818 17502 50820 17554
rect 50764 17332 50820 17502
rect 50988 17332 51044 18398
rect 51212 18338 51268 20132
rect 51548 19794 51604 19806
rect 51548 19742 51550 19794
rect 51602 19742 51604 19794
rect 51436 19010 51492 19022
rect 51436 18958 51438 19010
rect 51490 18958 51492 19010
rect 51436 18786 51492 18958
rect 51436 18734 51438 18786
rect 51490 18734 51492 18786
rect 51436 18722 51492 18734
rect 51212 18286 51214 18338
rect 51266 18286 51268 18338
rect 51212 17554 51268 18286
rect 51548 17892 51604 19742
rect 51548 17826 51604 17836
rect 51660 19796 51716 22766
rect 51996 21812 52052 25228
rect 52780 25172 52836 28812
rect 53004 26740 53060 30380
rect 53116 30100 53172 30110
rect 53116 28868 53172 30044
rect 53228 29874 53284 30380
rect 53788 29988 53844 32844
rect 53900 32564 53956 33628
rect 53900 32498 53956 32508
rect 54012 32786 54068 33964
rect 54348 33908 54404 33918
rect 54572 33908 54628 35084
rect 54684 34916 54740 34926
rect 54740 34860 54852 34916
rect 54684 34822 54740 34860
rect 54796 34468 54852 34860
rect 54908 34804 54964 35084
rect 54908 34710 54964 34748
rect 55020 34580 55076 35758
rect 55692 34692 55748 34702
rect 55244 34580 55300 34590
rect 55020 34578 55300 34580
rect 55020 34526 55246 34578
rect 55298 34526 55300 34578
rect 55020 34524 55300 34526
rect 55244 34514 55300 34524
rect 54796 34412 55076 34468
rect 55020 34132 55076 34412
rect 55020 34018 55076 34076
rect 55692 34132 55748 34636
rect 55692 34066 55748 34076
rect 55020 33966 55022 34018
rect 55074 33966 55076 34018
rect 55020 33954 55076 33966
rect 54404 33852 54628 33908
rect 54348 33814 54404 33852
rect 55804 33684 55860 33694
rect 55804 33590 55860 33628
rect 54012 32734 54014 32786
rect 54066 32734 54068 32786
rect 53900 31780 53956 31790
rect 53900 31686 53956 31724
rect 54012 30996 54068 32734
rect 54124 32786 54180 32798
rect 54124 32734 54126 32786
rect 54178 32734 54180 32786
rect 54124 32564 54180 32734
rect 55020 32676 55076 32686
rect 55020 32582 55076 32620
rect 54124 32004 54180 32508
rect 54684 32450 54740 32462
rect 54684 32398 54686 32450
rect 54738 32398 54740 32450
rect 54684 31948 54740 32398
rect 54124 31556 54180 31948
rect 54124 31490 54180 31500
rect 54348 31892 54740 31948
rect 55580 32450 55636 32462
rect 55580 32398 55582 32450
rect 55634 32398 55636 32450
rect 54348 31890 54404 31892
rect 54348 31838 54350 31890
rect 54402 31838 54404 31890
rect 53900 30940 54068 30996
rect 53900 30324 53956 30940
rect 53900 30258 53956 30268
rect 54012 30770 54068 30782
rect 54012 30718 54014 30770
rect 54066 30718 54068 30770
rect 53900 29988 53956 29998
rect 53788 29986 53956 29988
rect 53788 29934 53902 29986
rect 53954 29934 53956 29986
rect 53788 29932 53956 29934
rect 53900 29922 53956 29932
rect 53228 29822 53230 29874
rect 53282 29822 53284 29874
rect 53228 29810 53284 29822
rect 53564 29762 53620 29774
rect 53564 29710 53566 29762
rect 53618 29710 53620 29762
rect 53564 29092 53620 29710
rect 54012 29652 54068 30718
rect 54236 30436 54292 30446
rect 54068 29596 54180 29652
rect 54012 29586 54068 29596
rect 53788 29092 53844 29102
rect 53564 29090 53844 29092
rect 53564 29038 53790 29090
rect 53842 29038 53844 29090
rect 53564 29036 53844 29038
rect 53788 29026 53844 29036
rect 53228 28868 53284 28878
rect 53116 28866 53284 28868
rect 53116 28814 53230 28866
rect 53282 28814 53284 28866
rect 53116 28812 53284 28814
rect 53228 28532 53284 28812
rect 53228 28466 53284 28476
rect 53340 28868 53396 28878
rect 53116 27972 53172 27982
rect 53172 27916 53284 27972
rect 53116 27878 53172 27916
rect 53004 26738 53172 26740
rect 53004 26686 53006 26738
rect 53058 26686 53172 26738
rect 53004 26684 53172 26686
rect 53004 26674 53060 26684
rect 51660 17890 51716 19740
rect 51884 21756 51996 21812
rect 51884 20802 51940 21756
rect 51996 21746 52052 21756
rect 52108 25116 52836 25172
rect 52892 25172 52948 25182
rect 52108 22818 52164 25116
rect 52780 24836 52836 24846
rect 52892 24836 52948 25116
rect 52780 24834 52948 24836
rect 52780 24782 52782 24834
rect 52834 24782 52948 24834
rect 52780 24780 52948 24782
rect 52780 24770 52836 24780
rect 52892 24500 52948 24510
rect 52556 24386 52612 24398
rect 52556 24334 52558 24386
rect 52610 24334 52612 24386
rect 52556 23602 52612 24334
rect 52892 23826 52948 24444
rect 53116 23828 53172 26684
rect 53228 25732 53284 27916
rect 53340 27746 53396 28812
rect 54124 28868 54180 29596
rect 54124 28774 54180 28812
rect 53340 27694 53342 27746
rect 53394 27694 53396 27746
rect 53340 27682 53396 27694
rect 53452 27858 53508 27870
rect 53452 27806 53454 27858
rect 53506 27806 53508 27858
rect 53340 26626 53396 26638
rect 53340 26574 53342 26626
rect 53394 26574 53396 26626
rect 53340 25954 53396 26574
rect 53452 26628 53508 27806
rect 53676 26740 53732 26750
rect 53676 26646 53732 26684
rect 54236 26738 54292 30380
rect 54348 29764 54404 31838
rect 55020 31778 55076 31790
rect 55020 31726 55022 31778
rect 55074 31726 55076 31778
rect 54460 30660 54516 30670
rect 54516 30604 54628 30660
rect 54460 30566 54516 30604
rect 54460 29764 54516 29774
rect 54348 29762 54516 29764
rect 54348 29710 54462 29762
rect 54514 29710 54516 29762
rect 54348 29708 54516 29710
rect 54348 28532 54404 28542
rect 54348 27858 54404 28476
rect 54348 27806 54350 27858
rect 54402 27806 54404 27858
rect 54348 27794 54404 27806
rect 54460 27636 54516 29708
rect 54572 28642 54628 30604
rect 55020 30546 55076 31726
rect 55468 31780 55524 31790
rect 55468 30660 55524 31724
rect 55468 30594 55524 30604
rect 55020 30494 55022 30546
rect 55074 30494 55076 30546
rect 55020 30482 55076 30494
rect 55580 29988 55636 32398
rect 56028 31948 56084 36766
rect 57484 36818 57540 36830
rect 57484 36766 57486 36818
rect 57538 36766 57540 36818
rect 57148 36708 57204 36718
rect 56700 36036 56756 36046
rect 56700 35942 56756 35980
rect 57148 35810 57204 36652
rect 57148 35758 57150 35810
rect 57202 35758 57204 35810
rect 57148 35746 57204 35758
rect 56812 35700 56868 35710
rect 56700 35698 56868 35700
rect 56700 35646 56814 35698
rect 56866 35646 56868 35698
rect 56700 35644 56868 35646
rect 56140 35026 56196 35038
rect 56140 34974 56142 35026
rect 56194 34974 56196 35026
rect 56140 34916 56196 34974
rect 56700 35026 56756 35644
rect 56812 35634 56868 35644
rect 56700 34974 56702 35026
rect 56754 34974 56756 35026
rect 56700 34962 56756 34974
rect 56140 34822 56196 34860
rect 56588 34692 56644 34702
rect 56588 32788 56644 34636
rect 56588 32786 56868 32788
rect 56588 32734 56590 32786
rect 56642 32734 56868 32786
rect 56588 32732 56868 32734
rect 56588 32722 56644 32732
rect 56812 32002 56868 32732
rect 56812 31950 56814 32002
rect 56866 31950 56868 32002
rect 56812 31948 56868 31950
rect 55692 31890 55748 31902
rect 55692 31838 55694 31890
rect 55746 31838 55748 31890
rect 55692 31668 55748 31838
rect 56028 31892 56196 31948
rect 56028 31826 56084 31836
rect 55692 31602 55748 31612
rect 56140 30770 56196 31892
rect 56700 31892 56868 31948
rect 57036 32562 57092 32574
rect 57036 32510 57038 32562
rect 57090 32510 57092 32562
rect 56700 31826 56756 31836
rect 56476 31780 56532 31790
rect 56476 31686 56532 31724
rect 57036 31780 57092 32510
rect 57036 31714 57092 31724
rect 57148 32004 57204 32042
rect 57484 31948 57540 36766
rect 57596 36708 57652 36718
rect 57708 36708 57764 42028
rect 57596 36706 57764 36708
rect 57596 36654 57598 36706
rect 57650 36654 57764 36706
rect 57596 36652 57764 36654
rect 57596 36642 57652 36652
rect 57148 31892 57540 31948
rect 58156 31892 58212 31902
rect 56588 31668 56644 31678
rect 56812 31668 56868 31678
rect 56644 31666 56868 31668
rect 56644 31614 56814 31666
rect 56866 31614 56868 31666
rect 56644 31612 56868 31614
rect 56588 31602 56644 31612
rect 56812 31602 56868 31612
rect 56140 30718 56142 30770
rect 56194 30718 56196 30770
rect 56140 30706 56196 30718
rect 57148 30660 57204 31892
rect 58156 31798 58212 31836
rect 57372 31778 57428 31790
rect 57372 31726 57374 31778
rect 57426 31726 57428 31778
rect 57372 31668 57428 31726
rect 57708 31668 57764 31678
rect 57372 31666 57764 31668
rect 57372 31614 57710 31666
rect 57762 31614 57764 31666
rect 57372 31612 57764 31614
rect 57372 30772 57428 31612
rect 57708 31602 57764 31612
rect 57596 30772 57652 30782
rect 57372 30770 57652 30772
rect 57372 30718 57598 30770
rect 57650 30718 57652 30770
rect 57372 30716 57652 30718
rect 57260 30660 57316 30670
rect 57148 30658 57316 30660
rect 57148 30606 57262 30658
rect 57314 30606 57316 30658
rect 57148 30604 57316 30606
rect 57260 30594 57316 30604
rect 57596 30324 57652 30716
rect 57596 30258 57652 30268
rect 55692 29988 55748 29998
rect 55580 29986 55748 29988
rect 55580 29934 55694 29986
rect 55746 29934 55748 29986
rect 55580 29932 55748 29934
rect 55692 29922 55748 29932
rect 55020 29762 55076 29774
rect 55020 29710 55022 29762
rect 55074 29710 55076 29762
rect 55020 29092 55076 29710
rect 55580 29092 55636 29102
rect 55020 29090 55636 29092
rect 55020 29038 55582 29090
rect 55634 29038 55636 29090
rect 55020 29036 55636 29038
rect 55580 29026 55636 29036
rect 54572 28590 54574 28642
rect 54626 28590 54628 28642
rect 54572 27972 54628 28590
rect 55692 28756 55748 28766
rect 54572 27906 54628 27916
rect 54684 28532 54740 28542
rect 54236 26686 54238 26738
rect 54290 26686 54292 26738
rect 54236 26674 54292 26686
rect 54348 27580 54516 27636
rect 53452 26562 53508 26572
rect 53340 25902 53342 25954
rect 53394 25902 53396 25954
rect 53340 25890 53396 25902
rect 53900 25956 53956 25966
rect 53900 25844 53956 25900
rect 53788 25842 53956 25844
rect 53788 25790 53902 25842
rect 53954 25790 53956 25842
rect 53788 25788 53956 25790
rect 53228 25730 53732 25732
rect 53228 25678 53230 25730
rect 53282 25678 53732 25730
rect 53228 25676 53732 25678
rect 53228 25666 53284 25676
rect 53228 25058 53284 25070
rect 53228 25006 53230 25058
rect 53282 25006 53284 25058
rect 53228 24834 53284 25006
rect 53228 24782 53230 24834
rect 53282 24782 53284 24834
rect 53228 24770 53284 24782
rect 53676 24836 53732 25676
rect 53788 25058 53844 25788
rect 53900 25778 53956 25788
rect 53788 25006 53790 25058
rect 53842 25006 53844 25058
rect 53788 24994 53844 25006
rect 53676 24834 54180 24836
rect 53676 24782 53678 24834
rect 53730 24782 54180 24834
rect 53676 24780 54180 24782
rect 53676 24770 53732 24780
rect 53452 24724 53508 24734
rect 53228 23828 53284 23838
rect 52892 23774 52894 23826
rect 52946 23774 52948 23826
rect 52892 23762 52948 23774
rect 53004 23826 53284 23828
rect 53004 23774 53230 23826
rect 53282 23774 53284 23826
rect 53004 23772 53284 23774
rect 52556 23550 52558 23602
rect 52610 23550 52612 23602
rect 52556 23538 52612 23550
rect 52108 22766 52110 22818
rect 52162 22766 52164 22818
rect 51884 20750 51886 20802
rect 51938 20750 51940 20802
rect 51884 18898 51940 20750
rect 51996 21588 52052 21598
rect 51996 20580 52052 21532
rect 51996 19572 52052 20524
rect 52108 20468 52164 22766
rect 53004 22706 53060 23772
rect 53228 23762 53284 23772
rect 53004 22654 53006 22706
rect 53058 22654 53060 22706
rect 53004 22642 53060 22654
rect 53452 22708 53508 24668
rect 53564 24386 53620 24398
rect 53564 24334 53566 24386
rect 53618 24334 53620 24386
rect 53564 23826 53620 24334
rect 54124 24386 54180 24780
rect 54124 24334 54126 24386
rect 54178 24334 54180 24386
rect 53900 23940 53956 23950
rect 53900 23846 53956 23884
rect 54124 23940 54180 24334
rect 54124 23874 54180 23884
rect 53564 23774 53566 23826
rect 53618 23774 53620 23826
rect 53564 23762 53620 23774
rect 54348 23826 54404 27580
rect 54460 25732 54516 25742
rect 54684 25732 54740 28476
rect 54796 27970 54852 27982
rect 54796 27918 54798 27970
rect 54850 27918 54852 27970
rect 54796 26738 54852 27918
rect 55356 27972 55412 27982
rect 54796 26686 54798 26738
rect 54850 26686 54852 26738
rect 54796 26674 54852 26686
rect 54908 27860 54964 27870
rect 54908 25956 54964 27804
rect 55356 26852 55412 27916
rect 55692 27860 55748 28700
rect 56700 28530 56756 28542
rect 56700 28478 56702 28530
rect 56754 28478 56756 28530
rect 55804 27860 55860 27870
rect 56700 27860 56756 28478
rect 55692 27858 56756 27860
rect 55692 27806 55806 27858
rect 55858 27806 56756 27858
rect 55692 27804 56756 27806
rect 55804 27794 55860 27804
rect 56700 27634 56756 27804
rect 56700 27582 56702 27634
rect 56754 27582 56756 27634
rect 56700 26964 56756 27582
rect 56700 26908 57204 26964
rect 55356 26796 55860 26852
rect 55468 26514 55524 26526
rect 55468 26462 55470 26514
rect 55522 26462 55524 26514
rect 54908 25890 54964 25900
rect 55356 25956 55412 25966
rect 55356 25862 55412 25900
rect 54908 25732 54964 25742
rect 54684 25730 54964 25732
rect 54684 25678 54910 25730
rect 54962 25678 54964 25730
rect 54684 25676 54964 25678
rect 54460 24722 54516 25676
rect 54908 25172 54964 25676
rect 55468 25396 55524 26462
rect 55804 25954 55860 26796
rect 55804 25902 55806 25954
rect 55858 25902 55860 25954
rect 55804 25890 55860 25902
rect 56700 25956 56756 25966
rect 54908 25106 54964 25116
rect 55356 25340 55524 25396
rect 55356 24834 55412 25340
rect 55356 24782 55358 24834
rect 55410 24782 55412 24834
rect 55356 24770 55412 24782
rect 55804 25172 55860 25182
rect 54460 24670 54462 24722
rect 54514 24670 54516 24722
rect 54460 24658 54516 24670
rect 55804 24722 55860 25116
rect 55804 24670 55806 24722
rect 55858 24670 55860 24722
rect 55804 24658 55860 24670
rect 56700 24724 56756 25900
rect 56700 24630 56756 24668
rect 57148 25618 57204 26908
rect 57148 25566 57150 25618
rect 57202 25566 57204 25618
rect 57148 24612 57204 25566
rect 57820 24722 57876 24734
rect 57820 24670 57822 24722
rect 57874 24670 57876 24722
rect 57596 24612 57652 24622
rect 57148 24610 57652 24612
rect 57148 24558 57598 24610
rect 57650 24558 57652 24610
rect 57148 24556 57652 24558
rect 55692 24388 55748 24398
rect 55692 23938 55748 24332
rect 57484 24388 57540 24398
rect 57484 24294 57540 24332
rect 55692 23886 55694 23938
rect 55746 23886 55748 23938
rect 55692 23874 55748 23886
rect 57148 23940 57204 23950
rect 57148 23846 57204 23884
rect 54348 23774 54350 23826
rect 54402 23774 54404 23826
rect 53676 22708 53732 22718
rect 53452 22706 53732 22708
rect 53452 22654 53678 22706
rect 53730 22654 53732 22706
rect 53452 22652 53732 22654
rect 53676 22642 53732 22652
rect 54236 22708 54292 22718
rect 54348 22708 54404 23774
rect 54236 22706 54404 22708
rect 54236 22654 54238 22706
rect 54290 22654 54404 22706
rect 54236 22652 54404 22654
rect 55020 23714 55076 23726
rect 55020 23662 55022 23714
rect 55074 23662 55076 23714
rect 54236 22642 54292 22652
rect 52668 22596 52724 22606
rect 53340 22596 53396 22606
rect 52668 22594 52836 22596
rect 52668 22542 52670 22594
rect 52722 22542 52836 22594
rect 52668 22540 52836 22542
rect 52668 22530 52724 22540
rect 52780 20692 52836 22540
rect 53116 22594 53396 22596
rect 53116 22542 53342 22594
rect 53394 22542 53396 22594
rect 53116 22540 53396 22542
rect 52892 21924 52948 21934
rect 53116 21924 53172 22540
rect 53340 22530 53396 22540
rect 54796 22594 54852 22606
rect 54796 22542 54798 22594
rect 54850 22542 54852 22594
rect 52892 21922 53172 21924
rect 52892 21870 52894 21922
rect 52946 21870 53172 21922
rect 52892 21868 53172 21870
rect 53452 21980 53732 22036
rect 52892 21858 52948 21868
rect 52892 20692 52948 20702
rect 52780 20690 52948 20692
rect 52780 20638 52894 20690
rect 52946 20638 52948 20690
rect 52780 20636 52948 20638
rect 52892 20626 52948 20636
rect 53452 20468 53508 21980
rect 53676 21924 53732 21980
rect 53676 21868 54068 21924
rect 53564 21812 53620 21822
rect 53620 21756 53732 21812
rect 53564 21718 53620 21756
rect 53564 20580 53620 20590
rect 53564 20486 53620 20524
rect 52108 20412 53508 20468
rect 52780 20020 52836 20030
rect 52668 19682 52724 19694
rect 52668 19630 52670 19682
rect 52722 19630 52724 19682
rect 52332 19572 52388 19582
rect 51996 19570 52388 19572
rect 51996 19518 52334 19570
rect 52386 19518 52388 19570
rect 51996 19516 52388 19518
rect 52220 19012 52276 19022
rect 52332 19012 52388 19516
rect 52220 19010 52388 19012
rect 52220 18958 52222 19010
rect 52274 18958 52388 19010
rect 52220 18956 52388 18958
rect 52220 18946 52276 18956
rect 51884 18846 51886 18898
rect 51938 18846 51940 18898
rect 51884 18834 51940 18846
rect 51884 18676 51940 18686
rect 51884 18450 51940 18620
rect 52668 18676 52724 19630
rect 52668 18610 52724 18620
rect 51884 18398 51886 18450
rect 51938 18398 51940 18450
rect 51884 18338 51940 18398
rect 51884 18286 51886 18338
rect 51938 18286 51940 18338
rect 51884 18274 51940 18286
rect 51996 18564 52052 18574
rect 51660 17838 51662 17890
rect 51714 17838 51716 17890
rect 51212 17502 51214 17554
rect 51266 17502 51268 17554
rect 50764 17276 51044 17332
rect 51100 17330 51156 17342
rect 51100 17278 51102 17330
rect 51154 17278 51156 17330
rect 50092 16436 50148 16446
rect 49868 16380 50092 16436
rect 50092 16342 50148 16380
rect 50540 16434 50596 16446
rect 50540 16382 50542 16434
rect 50594 16382 50596 16434
rect 49644 16258 49700 16268
rect 50540 16324 50596 16382
rect 50540 16258 50596 16268
rect 50556 16156 50820 16166
rect 50612 16100 50660 16156
rect 50716 16100 50764 16156
rect 50556 16090 50820 16100
rect 50092 15876 50148 15886
rect 49532 15874 50092 15876
rect 49532 15822 49534 15874
rect 49586 15822 50092 15874
rect 49532 15820 50092 15822
rect 49532 15810 49588 15820
rect 50092 15782 50148 15820
rect 49644 15652 49700 15662
rect 49420 15650 49700 15652
rect 49420 15598 49646 15650
rect 49698 15598 49700 15650
rect 49420 15596 49700 15598
rect 49644 15586 49700 15596
rect 49868 15652 49924 15662
rect 49308 14590 49310 14642
rect 49362 14590 49364 14642
rect 49308 14578 49364 14590
rect 49868 14642 49924 15596
rect 49868 14590 49870 14642
rect 49922 14590 49924 14642
rect 49868 14578 49924 14590
rect 50540 15540 50596 15550
rect 50876 15540 50932 17276
rect 50988 16772 51044 16782
rect 51100 16772 51156 17278
rect 50988 16770 51156 16772
rect 50988 16718 50990 16770
rect 51042 16718 51156 16770
rect 50988 16716 51156 16718
rect 50988 16706 51044 16716
rect 51100 15988 51156 16716
rect 51100 15894 51156 15932
rect 51212 16436 51268 17502
rect 51660 17330 51716 17838
rect 51660 17278 51662 17330
rect 51714 17278 51716 17330
rect 51660 17266 51716 17278
rect 50540 15538 50932 15540
rect 50540 15486 50542 15538
rect 50594 15486 50932 15538
rect 50540 15484 50932 15486
rect 50988 15876 51044 15886
rect 50540 14644 50596 15484
rect 50540 14578 50596 14588
rect 47852 14532 47908 14542
rect 47068 14466 47124 14476
rect 47180 14530 47908 14532
rect 47180 14478 47854 14530
rect 47906 14478 47908 14530
rect 47180 14476 47908 14478
rect 46620 13746 47012 13748
rect 46620 13694 46622 13746
rect 46674 13694 47012 13746
rect 46620 13692 47012 13694
rect 47180 13746 47236 14476
rect 47852 14466 47908 14476
rect 48300 14530 48356 14542
rect 48300 14478 48302 14530
rect 48354 14478 48356 14530
rect 47180 13694 47182 13746
rect 47234 13694 47236 13746
rect 46620 13682 46676 13692
rect 47180 13682 47236 13694
rect 47852 13746 47908 13758
rect 47852 13694 47854 13746
rect 47906 13694 47908 13746
rect 45724 13634 45780 13646
rect 45724 13582 45726 13634
rect 45778 13582 45780 13634
rect 45612 11508 45668 11518
rect 45724 11508 45780 13582
rect 46732 12626 46788 12638
rect 46732 12574 46734 12626
rect 46786 12574 46788 12626
rect 46396 12404 46452 12414
rect 46732 12404 46788 12574
rect 46452 12348 46788 12404
rect 46396 12310 46452 12348
rect 45612 11506 45780 11508
rect 45612 11454 45614 11506
rect 45666 11454 45780 11506
rect 45612 11452 45780 11454
rect 45612 11442 45668 11452
rect 45444 10780 45556 10836
rect 45388 10770 45444 10780
rect 45388 10612 45444 10622
rect 45276 10610 45444 10612
rect 45276 10558 45390 10610
rect 45442 10558 45444 10610
rect 45276 10556 45444 10558
rect 45164 10518 45220 10556
rect 45388 10546 45444 10556
rect 45500 10610 45556 10780
rect 47852 10834 47908 13694
rect 48300 12738 48356 14478
rect 50428 14530 50484 14542
rect 50428 14478 50430 14530
rect 50482 14478 50484 14530
rect 50428 13748 50484 14478
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50540 13748 50596 13758
rect 50428 13746 50596 13748
rect 50428 13694 50542 13746
rect 50594 13694 50596 13746
rect 50428 13692 50596 13694
rect 50540 13682 50596 13692
rect 48300 12686 48302 12738
rect 48354 12686 48356 12738
rect 48300 12674 48356 12686
rect 50988 12738 51044 15820
rect 51212 15540 51268 16380
rect 51436 16434 51492 16446
rect 51436 16382 51438 16434
rect 51490 16382 51492 16434
rect 51436 16324 51492 16382
rect 51996 16324 52052 18508
rect 52668 17780 52724 17790
rect 52780 17780 52836 19964
rect 53004 19684 53060 20412
rect 53676 20188 53732 21756
rect 54012 21810 54068 21868
rect 54012 21758 54014 21810
rect 54066 21758 54068 21810
rect 54012 21746 54068 21758
rect 54572 21698 54628 21710
rect 54572 21646 54574 21698
rect 54626 21646 54628 21698
rect 54348 21586 54404 21598
rect 54348 21534 54350 21586
rect 54402 21534 54404 21586
rect 54348 20690 54404 21534
rect 54348 20638 54350 20690
rect 54402 20638 54404 20690
rect 54124 20468 54180 20478
rect 54124 20374 54180 20412
rect 53676 20132 54180 20188
rect 53340 19796 53396 19806
rect 53340 19702 53396 19740
rect 54124 19794 54180 20132
rect 54124 19742 54126 19794
rect 54178 19742 54180 19794
rect 53676 19684 53732 19694
rect 52892 19682 53060 19684
rect 52892 19630 53006 19682
rect 53058 19630 53060 19682
rect 52892 19628 53060 19630
rect 52892 18730 52948 19628
rect 53004 19618 53060 19628
rect 53564 19682 53732 19684
rect 53564 19630 53678 19682
rect 53730 19630 53732 19682
rect 53564 19628 53732 19630
rect 52892 18678 52894 18730
rect 52946 18678 52948 18730
rect 52892 18564 52948 18678
rect 53564 18676 53620 19628
rect 53676 19618 53732 19628
rect 53340 18620 53620 18676
rect 52892 18498 52948 18508
rect 53228 18564 53284 18574
rect 53228 18470 53284 18508
rect 52668 17778 52836 17780
rect 52668 17726 52670 17778
rect 52722 17726 52836 17778
rect 52668 17724 52836 17726
rect 53340 17778 53396 18620
rect 54124 18564 54180 19742
rect 54348 18676 54404 20638
rect 54348 18610 54404 18620
rect 54572 19796 54628 21646
rect 54796 21028 54852 22542
rect 55020 22484 55076 23662
rect 56700 23604 56756 23614
rect 56700 23510 56756 23548
rect 57596 23604 57652 24556
rect 57820 23940 57876 24670
rect 57932 24724 57988 24734
rect 57988 24710 58100 24724
rect 57988 24668 58046 24710
rect 57932 24658 57988 24668
rect 58044 24658 58046 24668
rect 58098 24658 58100 24710
rect 58044 24646 58100 24658
rect 57596 22706 57652 23548
rect 57596 22654 57598 22706
rect 57650 22654 57652 22706
rect 55468 22484 55524 22494
rect 55020 22418 55076 22428
rect 55132 22482 55524 22484
rect 55132 22430 55470 22482
rect 55522 22430 55524 22482
rect 55132 22428 55524 22430
rect 55132 21362 55188 22428
rect 55468 22418 55524 22428
rect 56476 22484 56532 22494
rect 56476 22390 56532 22428
rect 56700 21812 56756 21822
rect 55132 21310 55134 21362
rect 55186 21310 55188 21362
rect 55132 21298 55188 21310
rect 55468 21698 55524 21710
rect 55468 21646 55470 21698
rect 55522 21646 55524 21698
rect 54796 20962 54852 20972
rect 55356 20690 55412 20702
rect 55356 20638 55358 20690
rect 55410 20638 55412 20690
rect 54908 20580 54964 20590
rect 54796 20466 54852 20478
rect 54796 20414 54798 20466
rect 54850 20414 54852 20466
rect 54796 20020 54852 20414
rect 54796 19954 54852 19964
rect 54124 18498 54180 18508
rect 53676 17892 53732 17902
rect 53676 17798 53732 17836
rect 53340 17726 53342 17778
rect 53394 17726 53396 17778
rect 52668 17714 52724 17724
rect 53340 17714 53396 17726
rect 53004 17666 53060 17678
rect 53004 17614 53006 17666
rect 53058 17614 53060 17666
rect 52332 17554 52388 17566
rect 52332 17502 52334 17554
rect 52386 17502 52388 17554
rect 51436 16268 52052 16324
rect 51436 15986 51492 15998
rect 51436 15934 51438 15986
rect 51490 15934 51492 15986
rect 51436 15874 51492 15934
rect 51436 15822 51438 15874
rect 51490 15822 51492 15874
rect 51436 15810 51492 15822
rect 51772 15986 51828 15998
rect 51772 15934 51774 15986
rect 51826 15934 51828 15986
rect 51212 15474 51268 15484
rect 51772 15316 51828 15934
rect 51884 15540 51940 15550
rect 51884 15446 51940 15484
rect 51772 15260 51940 15316
rect 51772 14756 51828 14766
rect 51660 14754 51828 14756
rect 51660 14702 51774 14754
rect 51826 14702 51828 14754
rect 51660 14700 51828 14702
rect 51660 14644 51716 14700
rect 51772 14690 51828 14700
rect 51100 14588 51716 14644
rect 51100 14530 51156 14588
rect 51100 14478 51102 14530
rect 51154 14478 51156 14530
rect 51100 14466 51156 14478
rect 50988 12686 50990 12738
rect 51042 12686 51044 12738
rect 50988 12674 51044 12686
rect 51548 14308 51604 14318
rect 51548 12738 51604 14252
rect 51548 12686 51550 12738
rect 51602 12686 51604 12738
rect 51548 12674 51604 12686
rect 51884 12738 51940 15260
rect 51996 14308 52052 16268
rect 52108 16436 52164 16446
rect 52108 15876 52164 16380
rect 52332 16324 52388 17502
rect 52388 16268 52612 16324
rect 52332 16258 52388 16268
rect 52332 15876 52388 15886
rect 52164 15874 52388 15876
rect 52164 15822 52334 15874
rect 52386 15822 52388 15874
rect 52164 15820 52388 15822
rect 52108 15810 52164 15820
rect 52332 15810 52388 15820
rect 51996 14242 52052 14252
rect 52556 13860 52612 16268
rect 53004 15764 53060 17614
rect 53452 17668 53508 17678
rect 53508 17612 53620 17668
rect 53452 17602 53508 17612
rect 53228 16658 53284 16670
rect 53228 16606 53230 16658
rect 53282 16606 53284 16658
rect 53228 16436 53284 16606
rect 53228 16370 53284 16380
rect 53452 16434 53508 16446
rect 53452 16382 53454 16434
rect 53506 16382 53508 16434
rect 53004 15670 53060 15708
rect 53340 15764 53396 15774
rect 53452 15764 53508 16382
rect 53564 15876 53620 17612
rect 54236 17666 54292 17678
rect 54236 17614 54238 17666
rect 54290 17614 54292 17666
rect 53676 16658 53732 16670
rect 53676 16606 53678 16658
rect 53730 16606 53732 16658
rect 53676 16324 53732 16606
rect 54124 16658 54180 16670
rect 54124 16606 54126 16658
rect 54178 16606 54180 16658
rect 54124 16548 54180 16606
rect 54124 16482 54180 16492
rect 53676 16258 53732 16268
rect 53900 16436 53956 16446
rect 53676 15876 53732 15886
rect 53564 15874 53732 15876
rect 53564 15822 53678 15874
rect 53730 15822 53732 15874
rect 53564 15820 53732 15822
rect 53676 15810 53732 15820
rect 53340 15762 53508 15764
rect 53340 15710 53342 15762
rect 53394 15710 53508 15762
rect 53340 15708 53508 15710
rect 53340 15698 53396 15708
rect 52668 15650 52724 15662
rect 52668 15598 52670 15650
rect 52722 15598 52724 15650
rect 52668 14756 52724 15598
rect 52668 14690 52724 14700
rect 52892 14644 52948 14654
rect 52892 14550 52948 14588
rect 52668 14530 52724 14542
rect 52668 14478 52670 14530
rect 52722 14478 52724 14530
rect 52668 14308 52724 14478
rect 52668 14242 52724 14252
rect 52556 13636 52612 13804
rect 53900 13748 53956 16380
rect 54236 15762 54292 17614
rect 54572 16660 54628 19740
rect 54796 19796 54852 19806
rect 54908 19796 54964 20524
rect 55356 20244 55412 20638
rect 55468 20580 55524 21646
rect 55468 20514 55524 20524
rect 55692 21698 55748 21710
rect 55692 21646 55694 21698
rect 55746 21646 55748 21698
rect 55692 20468 55748 21646
rect 56476 21028 56532 21038
rect 56476 20934 56532 20972
rect 56700 20804 56756 21756
rect 57148 21588 57204 21598
rect 57596 21588 57652 22654
rect 57708 23884 57820 23940
rect 57708 22818 57764 23884
rect 57820 23874 57876 23884
rect 57708 22766 57710 22818
rect 57762 22766 57764 22818
rect 57708 21812 57764 22766
rect 57708 21746 57764 21756
rect 57148 21586 57652 21588
rect 57148 21534 57150 21586
rect 57202 21534 57652 21586
rect 57148 21532 57652 21534
rect 56812 20804 56868 20814
rect 56700 20802 56868 20804
rect 56700 20750 56814 20802
rect 56866 20750 56868 20802
rect 56700 20748 56868 20750
rect 57148 20804 57204 21532
rect 57260 20804 57316 20814
rect 57148 20802 57316 20804
rect 57148 20750 57262 20802
rect 57314 20750 57316 20802
rect 57148 20748 57316 20750
rect 55916 20692 55972 20702
rect 55916 20598 55972 20636
rect 56812 20692 56868 20748
rect 57260 20738 57316 20748
rect 55356 20188 55524 20244
rect 55468 20132 55524 20188
rect 55692 20132 55748 20412
rect 55468 20076 55748 20132
rect 56700 20468 56756 20478
rect 55468 19906 55524 20076
rect 55468 19854 55470 19906
rect 55522 19854 55524 19906
rect 55468 19842 55524 19854
rect 54796 19794 54964 19796
rect 54796 19742 54798 19794
rect 54850 19742 54964 19794
rect 54796 19740 54964 19742
rect 55132 19796 55188 19806
rect 54796 19730 54852 19740
rect 54796 18898 54852 18910
rect 54796 18846 54798 18898
rect 54850 18846 54852 18898
rect 54684 18786 54740 18798
rect 54684 18734 54686 18786
rect 54738 18734 54740 18786
rect 54684 18676 54740 18734
rect 54684 18610 54740 18620
rect 54796 17778 54852 18846
rect 55132 18562 55188 19740
rect 55132 18510 55134 18562
rect 55186 18510 55188 18562
rect 55132 18498 55188 18510
rect 56700 19570 56756 20412
rect 56812 20188 56868 20636
rect 56812 20132 57204 20188
rect 56700 19518 56702 19570
rect 56754 19518 56756 19570
rect 56700 18564 56756 19518
rect 57148 18674 57204 20132
rect 57148 18622 57150 18674
rect 57202 18622 57204 18674
rect 56924 18564 56980 18574
rect 57148 18564 57204 18622
rect 56700 18508 56924 18564
rect 56924 18498 56980 18508
rect 57036 18508 57204 18564
rect 57708 18564 57764 18574
rect 54796 17726 54798 17778
rect 54850 17726 54852 17778
rect 54796 17714 54852 17726
rect 55468 17780 55524 17790
rect 55468 17778 55748 17780
rect 55468 17726 55470 17778
rect 55522 17726 55748 17778
rect 55468 17724 55748 17726
rect 55468 17714 55524 17724
rect 55692 16994 55748 17724
rect 55692 16942 55694 16994
rect 55746 16942 55748 16994
rect 55692 16930 55748 16942
rect 54572 16566 54628 16604
rect 54908 16658 54964 16670
rect 54908 16606 54910 16658
rect 54962 16606 54964 16658
rect 54236 15710 54238 15762
rect 54290 15710 54292 15762
rect 54236 15652 54292 15710
rect 54236 15586 54292 15596
rect 54460 16548 54516 16558
rect 54460 15540 54516 16492
rect 54908 16436 54964 16606
rect 54908 16370 54964 16380
rect 55020 16660 55076 16670
rect 54460 14532 54516 15484
rect 54796 15650 54852 15662
rect 54796 15598 54798 15650
rect 54850 15598 54852 15650
rect 54460 14530 54740 14532
rect 54460 14478 54462 14530
rect 54514 14478 54740 14530
rect 54460 14476 54740 14478
rect 54460 14466 54516 14476
rect 54572 13860 54628 13870
rect 54572 13766 54628 13804
rect 54236 13748 54292 13758
rect 53900 13746 54292 13748
rect 53900 13694 54238 13746
rect 54290 13694 54292 13746
rect 53900 13692 54292 13694
rect 54684 13748 54740 14476
rect 54796 13970 54852 15598
rect 54908 14532 54964 14542
rect 55020 14532 55076 16604
rect 55132 16658 55188 16670
rect 55132 16606 55134 16658
rect 55186 16606 55188 16658
rect 55132 16324 55188 16606
rect 55356 16658 55412 16670
rect 55356 16606 55358 16658
rect 55410 16606 55412 16658
rect 55356 16548 55412 16606
rect 55580 16660 55636 16670
rect 55580 16566 55636 16604
rect 56140 16660 56196 16670
rect 56140 16566 56196 16604
rect 55356 16482 55412 16492
rect 56588 16548 56644 16558
rect 56588 16454 56644 16492
rect 55132 16258 55188 16268
rect 57036 16434 57092 18508
rect 57036 16382 57038 16434
rect 57090 16382 57092 16434
rect 55468 15764 55524 15774
rect 55468 15762 55972 15764
rect 55468 15710 55470 15762
rect 55522 15710 55972 15762
rect 55468 15708 55972 15710
rect 55468 15698 55524 15708
rect 54908 14530 55076 14532
rect 54908 14478 54910 14530
rect 54962 14478 55076 14530
rect 54908 14476 55076 14478
rect 54908 14466 54964 14476
rect 54796 13918 54798 13970
rect 54850 13918 54852 13970
rect 54796 13906 54852 13918
rect 54908 13748 54964 13758
rect 54684 13746 54964 13748
rect 54684 13694 54910 13746
rect 54962 13694 54964 13746
rect 54684 13692 54964 13694
rect 52668 13636 52724 13646
rect 52556 13634 52724 13636
rect 52556 13582 52670 13634
rect 52722 13582 52724 13634
rect 52556 13580 52724 13582
rect 52668 13570 52724 13580
rect 51884 12686 51886 12738
rect 51938 12686 51940 12738
rect 48860 12404 48916 12414
rect 48860 11730 48916 12348
rect 50556 12124 50820 12134
rect 50612 12068 50660 12124
rect 50716 12068 50764 12124
rect 50556 12058 50820 12068
rect 48860 11678 48862 11730
rect 48914 11678 48916 11730
rect 48860 11620 48916 11678
rect 51884 11732 51940 12686
rect 52780 12740 52836 12750
rect 53900 12740 53956 13692
rect 54236 13682 54292 13692
rect 54908 13524 54964 13692
rect 55020 13746 55076 14476
rect 55020 13694 55022 13746
rect 55074 13694 55076 13746
rect 55020 13682 55076 13694
rect 55580 13524 55636 13534
rect 54908 13522 55636 13524
rect 54908 13470 55582 13522
rect 55634 13470 55636 13522
rect 54908 13468 55636 13470
rect 52780 11842 52836 12684
rect 53788 12738 53956 12740
rect 53788 12686 53902 12738
rect 53954 12686 53956 12738
rect 53788 12684 53956 12686
rect 52780 11790 52782 11842
rect 52834 11790 52836 11842
rect 52780 11778 52836 11790
rect 53676 12514 53732 12526
rect 53676 12462 53678 12514
rect 53730 12462 53732 12514
rect 51884 11666 51940 11676
rect 53340 11732 53396 11742
rect 53340 11638 53396 11676
rect 48860 11554 48916 11564
rect 52332 11620 52388 11630
rect 52332 11526 52388 11564
rect 53116 11620 53172 11630
rect 47852 10782 47854 10834
rect 47906 10782 47908 10834
rect 47852 10770 47908 10782
rect 53116 10722 53172 11564
rect 53676 11620 53732 12462
rect 53788 11842 53844 12684
rect 53900 12674 53956 12684
rect 55356 12740 55412 13468
rect 55580 13458 55636 13468
rect 55916 12850 55972 15708
rect 56252 14756 56308 14766
rect 56252 14662 56308 14700
rect 57036 14642 57092 16382
rect 57484 16436 57540 16446
rect 57708 16436 57764 18508
rect 57484 16434 57764 16436
rect 57484 16382 57486 16434
rect 57538 16382 57764 16434
rect 57484 16380 57764 16382
rect 57484 16324 57540 16380
rect 57484 16258 57540 16268
rect 57036 14590 57038 14642
rect 57090 14590 57092 14642
rect 57036 14578 57092 14590
rect 56140 14532 56196 14542
rect 56028 14530 56196 14532
rect 56028 14478 56142 14530
rect 56194 14478 56196 14530
rect 56028 14476 56196 14478
rect 56028 13860 56084 14476
rect 56140 14466 56196 14476
rect 56028 13766 56084 13804
rect 55916 12798 55918 12850
rect 55970 12798 55972 12850
rect 55916 12786 55972 12798
rect 55356 12626 55412 12684
rect 55356 12574 55358 12626
rect 55410 12574 55412 12626
rect 55356 12562 55412 12574
rect 53788 11790 53790 11842
rect 53842 11790 53844 11842
rect 53788 11778 53844 11790
rect 53676 11554 53732 11564
rect 53116 10670 53118 10722
rect 53170 10670 53172 10722
rect 53116 10658 53172 10670
rect 45500 10558 45502 10610
rect 45554 10558 45556 10610
rect 45500 10546 45556 10558
rect 50556 10108 50820 10118
rect 50612 10052 50660 10108
rect 50716 10052 50764 10108
rect 50556 10042 50820 10052
rect 44492 9774 44494 9826
rect 44546 9774 44548 9826
rect 44492 9762 44548 9774
rect 37548 9492 37604 9502
rect 37436 9490 37604 9492
rect 37436 9438 37550 9490
rect 37602 9438 37604 9490
rect 37436 9436 37604 9438
rect 37548 9426 37604 9436
rect 37100 8654 37102 8706
rect 37154 8654 37156 8706
rect 37100 8642 37156 8654
rect 31724 8318 31726 8370
rect 31778 8318 31780 8370
rect 31612 7924 31668 7934
rect 29596 7718 29652 7756
rect 30380 7812 30436 7822
rect 29148 7606 29204 7644
rect 30268 7588 30324 7598
rect 30268 7494 30324 7532
rect 30380 7586 30436 7756
rect 30604 7700 30660 7710
rect 30604 7606 30660 7644
rect 31612 7698 31668 7868
rect 31612 7646 31614 7698
rect 31666 7646 31668 7698
rect 31612 7634 31668 7646
rect 30380 7534 30382 7586
rect 30434 7534 30436 7586
rect 30380 7522 30436 7534
rect 31724 7588 31780 8318
rect 31836 8316 32004 8372
rect 32284 8372 32900 8428
rect 31836 7924 31892 8316
rect 31836 7858 31892 7868
rect 32284 7810 32340 8372
rect 50556 8092 50820 8102
rect 50612 8036 50660 8092
rect 50716 8036 50764 8092
rect 50556 8026 50820 8036
rect 32284 7758 32286 7810
rect 32338 7758 32340 7810
rect 32284 7746 32340 7758
rect 31724 7522 31780 7532
rect 4284 7410 4340 7420
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 3836 6738 3892 6748
rect 19836 6076 20100 6086
rect 19892 6020 19940 6076
rect 19996 6020 20044 6076
rect 19836 6010 20100 6020
rect 50556 6076 50820 6086
rect 50612 6020 50660 6076
rect 50716 6020 50764 6076
rect 50556 6010 50820 6020
rect 4476 5068 4740 5078
rect 4532 5012 4580 5068
rect 4636 5012 4684 5068
rect 4476 5002 4740 5012
rect 35196 5068 35460 5078
rect 35252 5012 35300 5068
rect 35356 5012 35404 5068
rect 35196 5002 35460 5012
rect 19836 4060 20100 4070
rect 19892 4004 19940 4060
rect 19996 4004 20044 4060
rect 19836 3994 20100 4004
rect 50556 4060 50820 4070
rect 50612 4004 50660 4060
rect 50716 4004 50764 4060
rect 50556 3994 50820 4004
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
<< via2 >>
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 4476 55466 4532 55468
rect 4476 55414 4478 55466
rect 4478 55414 4530 55466
rect 4530 55414 4532 55466
rect 4476 55412 4532 55414
rect 4580 55466 4636 55468
rect 4580 55414 4582 55466
rect 4582 55414 4634 55466
rect 4634 55414 4636 55466
rect 4580 55412 4636 55414
rect 4684 55466 4740 55468
rect 4684 55414 4686 55466
rect 4686 55414 4738 55466
rect 4738 55414 4740 55466
rect 4684 55412 4740 55414
rect 35196 55466 35252 55468
rect 35196 55414 35198 55466
rect 35198 55414 35250 55466
rect 35250 55414 35252 55466
rect 35196 55412 35252 55414
rect 35300 55466 35356 55468
rect 35300 55414 35302 55466
rect 35302 55414 35354 55466
rect 35354 55414 35356 55466
rect 35300 55412 35356 55414
rect 35404 55466 35460 55468
rect 35404 55414 35406 55466
rect 35406 55414 35458 55466
rect 35458 55414 35460 55466
rect 35404 55412 35460 55414
rect 19836 54458 19892 54460
rect 19836 54406 19838 54458
rect 19838 54406 19890 54458
rect 19890 54406 19892 54458
rect 19836 54404 19892 54406
rect 19940 54458 19996 54460
rect 19940 54406 19942 54458
rect 19942 54406 19994 54458
rect 19994 54406 19996 54458
rect 19940 54404 19996 54406
rect 20044 54458 20100 54460
rect 20044 54406 20046 54458
rect 20046 54406 20098 54458
rect 20098 54406 20100 54458
rect 20044 54404 20100 54406
rect 50556 54458 50612 54460
rect 50556 54406 50558 54458
rect 50558 54406 50610 54458
rect 50610 54406 50612 54458
rect 50556 54404 50612 54406
rect 50660 54458 50716 54460
rect 50660 54406 50662 54458
rect 50662 54406 50714 54458
rect 50714 54406 50716 54458
rect 50660 54404 50716 54406
rect 50764 54458 50820 54460
rect 50764 54406 50766 54458
rect 50766 54406 50818 54458
rect 50818 54406 50820 54458
rect 50764 54404 50820 54406
rect 3836 53788 3892 53844
rect 56140 53788 56196 53844
rect 4476 53450 4532 53452
rect 4476 53398 4478 53450
rect 4478 53398 4530 53450
rect 4530 53398 4532 53450
rect 4476 53396 4532 53398
rect 4580 53450 4636 53452
rect 4580 53398 4582 53450
rect 4582 53398 4634 53450
rect 4634 53398 4636 53450
rect 4580 53396 4636 53398
rect 4684 53450 4740 53452
rect 4684 53398 4686 53450
rect 4686 53398 4738 53450
rect 4738 53398 4740 53450
rect 4684 53396 4740 53398
rect 35196 53450 35252 53452
rect 35196 53398 35198 53450
rect 35198 53398 35250 53450
rect 35250 53398 35252 53450
rect 35196 53396 35252 53398
rect 35300 53450 35356 53452
rect 35300 53398 35302 53450
rect 35302 53398 35354 53450
rect 35354 53398 35356 53450
rect 35300 53396 35356 53398
rect 35404 53450 35460 53452
rect 35404 53398 35406 53450
rect 35406 53398 35458 53450
rect 35458 53398 35460 53450
rect 35404 53396 35460 53398
rect 19836 52442 19892 52444
rect 19836 52390 19838 52442
rect 19838 52390 19890 52442
rect 19890 52390 19892 52442
rect 19836 52388 19892 52390
rect 19940 52442 19996 52444
rect 19940 52390 19942 52442
rect 19942 52390 19994 52442
rect 19994 52390 19996 52442
rect 19940 52388 19996 52390
rect 20044 52442 20100 52444
rect 20044 52390 20046 52442
rect 20046 52390 20098 52442
rect 20098 52390 20100 52442
rect 20044 52388 20100 52390
rect 50556 52442 50612 52444
rect 50556 52390 50558 52442
rect 50558 52390 50610 52442
rect 50610 52390 50612 52442
rect 50556 52388 50612 52390
rect 50660 52442 50716 52444
rect 50660 52390 50662 52442
rect 50662 52390 50714 52442
rect 50714 52390 50716 52442
rect 50660 52388 50716 52390
rect 50764 52442 50820 52444
rect 50764 52390 50766 52442
rect 50766 52390 50818 52442
rect 50818 52390 50820 52442
rect 50764 52388 50820 52390
rect 4476 51434 4532 51436
rect 4476 51382 4478 51434
rect 4478 51382 4530 51434
rect 4530 51382 4532 51434
rect 4476 51380 4532 51382
rect 4580 51434 4636 51436
rect 4580 51382 4582 51434
rect 4582 51382 4634 51434
rect 4634 51382 4636 51434
rect 4580 51380 4636 51382
rect 4684 51434 4740 51436
rect 4684 51382 4686 51434
rect 4686 51382 4738 51434
rect 4738 51382 4740 51434
rect 4684 51380 4740 51382
rect 35196 51434 35252 51436
rect 35196 51382 35198 51434
rect 35198 51382 35250 51434
rect 35250 51382 35252 51434
rect 35196 51380 35252 51382
rect 35300 51434 35356 51436
rect 35300 51382 35302 51434
rect 35302 51382 35354 51434
rect 35354 51382 35356 51434
rect 35300 51380 35356 51382
rect 35404 51434 35460 51436
rect 35404 51382 35406 51434
rect 35406 51382 35458 51434
rect 35458 51382 35460 51434
rect 35404 51380 35460 51382
rect 19836 50426 19892 50428
rect 19836 50374 19838 50426
rect 19838 50374 19890 50426
rect 19890 50374 19892 50426
rect 19836 50372 19892 50374
rect 19940 50426 19996 50428
rect 19940 50374 19942 50426
rect 19942 50374 19994 50426
rect 19994 50374 19996 50426
rect 19940 50372 19996 50374
rect 20044 50426 20100 50428
rect 20044 50374 20046 50426
rect 20046 50374 20098 50426
rect 20098 50374 20100 50426
rect 20044 50372 20100 50374
rect 50556 50426 50612 50428
rect 50556 50374 50558 50426
rect 50558 50374 50610 50426
rect 50610 50374 50612 50426
rect 50556 50372 50612 50374
rect 50660 50426 50716 50428
rect 50660 50374 50662 50426
rect 50662 50374 50714 50426
rect 50714 50374 50716 50426
rect 50660 50372 50716 50374
rect 50764 50426 50820 50428
rect 50764 50374 50766 50426
rect 50766 50374 50818 50426
rect 50818 50374 50820 50426
rect 50764 50372 50820 50374
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 19836 48410 19892 48412
rect 19836 48358 19838 48410
rect 19838 48358 19890 48410
rect 19890 48358 19892 48410
rect 19836 48356 19892 48358
rect 19940 48410 19996 48412
rect 19940 48358 19942 48410
rect 19942 48358 19994 48410
rect 19994 48358 19996 48410
rect 19940 48356 19996 48358
rect 20044 48410 20100 48412
rect 20044 48358 20046 48410
rect 20046 48358 20098 48410
rect 20098 48358 20100 48410
rect 20044 48356 20100 48358
rect 19516 47906 19572 47908
rect 19516 47854 19518 47906
rect 19518 47854 19570 47906
rect 19570 47854 19572 47906
rect 19516 47852 19572 47854
rect 20188 47852 20244 47908
rect 4476 47402 4532 47404
rect 4476 47350 4478 47402
rect 4478 47350 4530 47402
rect 4530 47350 4532 47402
rect 4476 47348 4532 47350
rect 4580 47402 4636 47404
rect 4580 47350 4582 47402
rect 4582 47350 4634 47402
rect 4634 47350 4636 47402
rect 4580 47348 4636 47350
rect 4684 47402 4740 47404
rect 4684 47350 4686 47402
rect 4686 47350 4738 47402
rect 4738 47350 4740 47402
rect 4684 47348 4740 47350
rect 20188 47180 20244 47236
rect 23100 48748 23156 48804
rect 21644 47180 21700 47236
rect 4476 45386 4532 45388
rect 4476 45334 4478 45386
rect 4478 45334 4530 45386
rect 4530 45334 4532 45386
rect 4476 45332 4532 45334
rect 4580 45386 4636 45388
rect 4580 45334 4582 45386
rect 4582 45334 4634 45386
rect 4634 45334 4636 45386
rect 4580 45332 4636 45334
rect 4684 45386 4740 45388
rect 4684 45334 4686 45386
rect 4686 45334 4738 45386
rect 4738 45334 4740 45386
rect 4684 45332 4740 45334
rect 17500 45276 17556 45332
rect 17164 44882 17220 44884
rect 17164 44830 17166 44882
rect 17166 44830 17218 44882
rect 17218 44830 17220 44882
rect 17164 44828 17220 44830
rect 17948 45276 18004 45332
rect 19836 46394 19892 46396
rect 19836 46342 19838 46394
rect 19838 46342 19890 46394
rect 19890 46342 19892 46394
rect 19836 46340 19892 46342
rect 19940 46394 19996 46396
rect 19940 46342 19942 46394
rect 19942 46342 19994 46394
rect 19994 46342 19996 46394
rect 19940 46340 19996 46342
rect 20044 46394 20100 46396
rect 20044 46342 20046 46394
rect 20046 46342 20098 46394
rect 20098 46342 20100 46394
rect 20044 46340 20100 46342
rect 17612 44828 17668 44884
rect 20636 47068 20692 47124
rect 21868 46956 21924 47012
rect 20524 46060 20580 46116
rect 20188 45276 20244 45332
rect 18060 44882 18116 44884
rect 18060 44830 18062 44882
rect 18062 44830 18114 44882
rect 18114 44830 18116 44882
rect 18060 44828 18116 44830
rect 21308 45276 21364 45332
rect 19836 44378 19892 44380
rect 19836 44326 19838 44378
rect 19838 44326 19890 44378
rect 19890 44326 19892 44378
rect 19836 44324 19892 44326
rect 19940 44378 19996 44380
rect 19940 44326 19942 44378
rect 19942 44326 19994 44378
rect 19994 44326 19996 44378
rect 19940 44324 19996 44326
rect 20044 44378 20100 44380
rect 20044 44326 20046 44378
rect 20046 44326 20098 44378
rect 20098 44326 20100 44378
rect 20044 44324 20100 44326
rect 18060 43708 18116 43764
rect 19628 43820 19684 43876
rect 4476 43370 4532 43372
rect 4476 43318 4478 43370
rect 4478 43318 4530 43370
rect 4530 43318 4532 43370
rect 4476 43316 4532 43318
rect 4580 43370 4636 43372
rect 4580 43318 4582 43370
rect 4582 43318 4634 43370
rect 4634 43318 4636 43370
rect 4580 43316 4636 43318
rect 4684 43370 4740 43372
rect 4684 43318 4686 43370
rect 4686 43318 4738 43370
rect 4738 43318 4740 43370
rect 4684 43316 4740 43318
rect 1820 41746 1876 41748
rect 1820 41694 1822 41746
rect 1822 41694 1874 41746
rect 1874 41694 1876 41746
rect 1820 41692 1876 41694
rect 3724 41746 3780 41748
rect 3724 41694 3726 41746
rect 3726 41694 3778 41746
rect 3778 41694 3780 41746
rect 3724 41692 3780 41694
rect 1820 40460 1876 40516
rect 1708 40348 1764 40404
rect 3724 40684 3780 40740
rect 2380 40348 2436 40404
rect 2716 40460 2772 40516
rect 4620 41858 4676 41860
rect 4620 41806 4622 41858
rect 4622 41806 4674 41858
rect 4674 41806 4676 41858
rect 4620 41804 4676 41806
rect 6188 41804 6244 41860
rect 4476 41354 4532 41356
rect 4476 41302 4478 41354
rect 4478 41302 4530 41354
rect 4530 41302 4532 41354
rect 4476 41300 4532 41302
rect 4580 41354 4636 41356
rect 4580 41302 4582 41354
rect 4582 41302 4634 41354
rect 4634 41302 4636 41354
rect 4580 41300 4636 41302
rect 4684 41354 4740 41356
rect 4684 41302 4686 41354
rect 4686 41302 4738 41354
rect 4738 41302 4740 41354
rect 4684 41300 4740 41302
rect 4620 40684 4676 40740
rect 4060 40348 4116 40404
rect 4476 39338 4532 39340
rect 4476 39286 4478 39338
rect 4478 39286 4530 39338
rect 4530 39286 4532 39338
rect 4476 39284 4532 39286
rect 4580 39338 4636 39340
rect 4580 39286 4582 39338
rect 4582 39286 4634 39338
rect 4634 39286 4636 39338
rect 4580 39284 4636 39286
rect 4684 39338 4740 39340
rect 4684 39286 4686 39338
rect 4686 39286 4738 39338
rect 4738 39286 4740 39338
rect 4684 39284 4740 39286
rect 2380 38892 2436 38948
rect 5628 40514 5684 40516
rect 5628 40462 5630 40514
rect 5630 40462 5682 40514
rect 5682 40462 5684 40514
rect 5628 40460 5684 40462
rect 6300 41580 6356 41636
rect 7196 41634 7252 41636
rect 7196 41582 7198 41634
rect 7198 41582 7250 41634
rect 7250 41582 7252 41634
rect 7196 41580 7252 41582
rect 6860 40572 6916 40628
rect 6300 40460 6356 40516
rect 6076 40348 6132 40404
rect 4956 39564 5012 39620
rect 9772 42588 9828 42644
rect 8092 41916 8148 41972
rect 8988 41916 9044 41972
rect 9660 41970 9716 41972
rect 9660 41918 9662 41970
rect 9662 41918 9714 41970
rect 9714 41918 9716 41970
rect 9660 41916 9716 41918
rect 9548 41468 9604 41524
rect 7532 40460 7588 40516
rect 7868 40514 7924 40516
rect 7868 40462 7870 40514
rect 7870 40462 7922 40514
rect 7922 40462 7924 40514
rect 7868 40460 7924 40462
rect 8652 40626 8708 40628
rect 8652 40574 8654 40626
rect 8654 40574 8706 40626
rect 8706 40574 8708 40626
rect 8652 40572 8708 40574
rect 7980 40012 8036 40068
rect 6188 39564 6244 39620
rect 5628 38946 5684 38948
rect 5628 38894 5630 38946
rect 5630 38894 5682 38946
rect 5682 38894 5684 38946
rect 5628 38892 5684 38894
rect 4956 38722 5012 38724
rect 4956 38670 4958 38722
rect 4958 38670 5010 38722
rect 5010 38670 5012 38722
rect 4956 38668 5012 38670
rect 5740 38722 5796 38724
rect 5740 38670 5742 38722
rect 5742 38670 5794 38722
rect 5794 38670 5796 38722
rect 5740 38668 5796 38670
rect 8876 40066 8932 40068
rect 8876 40014 8878 40066
rect 8878 40014 8930 40066
rect 8930 40014 8932 40066
rect 8876 40012 8932 40014
rect 10668 42642 10724 42644
rect 10668 42590 10670 42642
rect 10670 42590 10722 42642
rect 10722 42590 10724 42642
rect 10668 42588 10724 42590
rect 19292 41970 19348 41972
rect 19292 41918 19294 41970
rect 19294 41918 19346 41970
rect 19346 41918 19348 41970
rect 19292 41916 19348 41918
rect 11004 41858 11060 41860
rect 11004 41806 11006 41858
rect 11006 41806 11058 41858
rect 11058 41806 11060 41858
rect 11004 41804 11060 41806
rect 12124 41804 12180 41860
rect 10892 41522 10948 41524
rect 10892 41470 10894 41522
rect 10894 41470 10946 41522
rect 10946 41470 10948 41522
rect 10892 41468 10948 41470
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19516 41580 19572 41636
rect 19852 40962 19908 40964
rect 19852 40910 19854 40962
rect 19854 40910 19906 40962
rect 19906 40910 19908 40962
rect 19852 40908 19908 40910
rect 20188 40908 20244 40964
rect 10220 40572 10276 40628
rect 18284 40796 18340 40852
rect 11788 40012 11844 40068
rect 12572 40066 12628 40068
rect 12572 40014 12574 40066
rect 12574 40014 12626 40066
rect 12626 40014 12628 40066
rect 12572 40012 12628 40014
rect 9660 39564 9716 39620
rect 10332 39564 10388 39620
rect 10220 38892 10276 38948
rect 8652 38668 8708 38724
rect 1820 36876 1876 36932
rect 6636 38610 6692 38612
rect 6636 38558 6638 38610
rect 6638 38558 6690 38610
rect 6690 38558 6692 38610
rect 6636 38556 6692 38558
rect 4844 37996 4900 38052
rect 5740 38050 5796 38052
rect 5740 37998 5742 38050
rect 5742 37998 5794 38050
rect 5794 37998 5796 38050
rect 5740 37996 5796 37998
rect 6300 37996 6356 38052
rect 2716 36876 2772 36932
rect 4476 37322 4532 37324
rect 4476 37270 4478 37322
rect 4478 37270 4530 37322
rect 4530 37270 4532 37322
rect 4476 37268 4532 37270
rect 4580 37322 4636 37324
rect 4580 37270 4582 37322
rect 4582 37270 4634 37322
rect 4634 37270 4636 37322
rect 4580 37268 4636 37270
rect 4684 37322 4740 37324
rect 4684 37270 4686 37322
rect 4686 37270 4738 37322
rect 4738 37270 4740 37322
rect 4684 37268 4740 37270
rect 3612 36764 3668 36820
rect 4508 36876 4564 36932
rect 5068 36818 5124 36820
rect 5068 36766 5070 36818
rect 5070 36766 5122 36818
rect 5122 36766 5124 36818
rect 5068 36764 5124 36766
rect 6076 36764 6132 36820
rect 3052 36652 3108 36708
rect 3836 36652 3892 36708
rect 5628 36706 5684 36708
rect 5628 36654 5630 36706
rect 5630 36654 5682 36706
rect 5682 36654 5684 36706
rect 5628 36652 5684 36654
rect 4172 36316 4228 36372
rect 3388 35084 3444 35140
rect 6636 37996 6692 38052
rect 17164 39900 17220 39956
rect 13356 39618 13412 39620
rect 13356 39566 13358 39618
rect 13358 39566 13410 39618
rect 13410 39566 13412 39618
rect 13356 39564 13412 39566
rect 13468 38946 13524 38948
rect 13468 38894 13470 38946
rect 13470 38894 13522 38946
rect 13522 38894 13524 38946
rect 13468 38892 13524 38894
rect 12796 38722 12852 38724
rect 12796 38670 12798 38722
rect 12798 38670 12850 38722
rect 12850 38670 12852 38722
rect 12796 38668 12852 38670
rect 13580 38722 13636 38724
rect 13580 38670 13582 38722
rect 13582 38670 13634 38722
rect 13634 38670 13636 38722
rect 13580 38668 13636 38670
rect 16828 38668 16884 38724
rect 9324 36930 9380 36932
rect 9324 36878 9326 36930
rect 9326 36878 9378 36930
rect 9378 36878 9380 36930
rect 9324 36876 9380 36878
rect 9660 37548 9716 37604
rect 10780 37548 10836 37604
rect 9884 36876 9940 36932
rect 12796 36594 12852 36596
rect 12796 36542 12798 36594
rect 12798 36542 12850 36594
rect 12850 36542 12852 36594
rect 12796 36540 12852 36542
rect 10220 36428 10276 36484
rect 11340 36428 11396 36484
rect 9884 35868 9940 35924
rect 11004 35922 11060 35924
rect 11004 35870 11006 35922
rect 11006 35870 11058 35922
rect 11058 35870 11060 35922
rect 11004 35868 11060 35870
rect 13804 37602 13860 37604
rect 13804 37550 13806 37602
rect 13806 37550 13858 37602
rect 13858 37550 13860 37602
rect 13804 37548 13860 37550
rect 16716 36930 16772 36932
rect 16716 36878 16718 36930
rect 16718 36878 16770 36930
rect 16770 36878 16772 36930
rect 16716 36876 16772 36878
rect 13580 36594 13636 36596
rect 13580 36542 13582 36594
rect 13582 36542 13634 36594
rect 13634 36542 13636 36594
rect 13580 36540 13636 36542
rect 13468 36482 13524 36484
rect 13468 36430 13470 36482
rect 13470 36430 13522 36482
rect 13522 36430 13524 36482
rect 13468 36428 13524 36430
rect 13020 35868 13076 35924
rect 14140 35868 14196 35924
rect 15260 35868 15316 35924
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 5628 35138 5684 35140
rect 5628 35086 5630 35138
rect 5630 35086 5682 35138
rect 5682 35086 5684 35138
rect 5628 35084 5684 35086
rect 6300 35084 6356 35140
rect 4172 34636 4228 34692
rect 3724 34524 3780 34580
rect 3276 34018 3332 34020
rect 3276 33966 3278 34018
rect 3278 33966 3330 34018
rect 3330 33966 3332 34018
rect 3276 33964 3332 33966
rect 5740 34578 5796 34580
rect 5740 34526 5742 34578
rect 5742 34526 5794 34578
rect 5794 34526 5796 34578
rect 5740 34524 5796 34526
rect 4060 34018 4116 34020
rect 4060 33966 4062 34018
rect 4062 33966 4114 34018
rect 4114 33966 4116 34018
rect 4060 33964 4116 33966
rect 5740 33740 5796 33796
rect 4476 33290 4532 33292
rect 4476 33238 4478 33290
rect 4478 33238 4530 33290
rect 4530 33238 4532 33290
rect 4476 33236 4532 33238
rect 4580 33290 4636 33292
rect 4580 33238 4582 33290
rect 4582 33238 4634 33290
rect 4634 33238 4636 33290
rect 4580 33236 4636 33238
rect 4684 33290 4740 33292
rect 4684 33238 4686 33290
rect 4686 33238 4738 33290
rect 4738 33238 4740 33290
rect 4684 33236 4740 33238
rect 11900 35084 11956 35140
rect 13468 35138 13524 35140
rect 13468 35086 13470 35138
rect 13470 35086 13522 35138
rect 13522 35086 13524 35138
rect 13468 35084 13524 35086
rect 6412 33740 6468 33796
rect 3836 32508 3892 32564
rect 5628 32562 5684 32564
rect 5628 32510 5630 32562
rect 5630 32510 5682 32562
rect 5682 32510 5684 32562
rect 5628 32508 5684 32510
rect 3388 31778 3444 31780
rect 3388 31726 3390 31778
rect 3390 31726 3442 31778
rect 3442 31726 3444 31778
rect 3388 31724 3444 31726
rect 4172 31724 4228 31780
rect 1820 29986 1876 29988
rect 1820 29934 1822 29986
rect 1822 29934 1874 29986
rect 1874 29934 1876 29986
rect 1820 29932 1876 29934
rect 2380 30604 2436 30660
rect 3724 30716 3780 30772
rect 2828 29986 2884 29988
rect 2828 29934 2830 29986
rect 2830 29934 2882 29986
rect 2882 29934 2884 29986
rect 2828 29932 2884 29934
rect 4476 31274 4532 31276
rect 4476 31222 4478 31274
rect 4478 31222 4530 31274
rect 4530 31222 4532 31274
rect 4476 31220 4532 31222
rect 4580 31274 4636 31276
rect 4580 31222 4582 31274
rect 4582 31222 4634 31274
rect 4634 31222 4636 31274
rect 4580 31220 4636 31222
rect 4684 31274 4740 31276
rect 4684 31222 4686 31274
rect 4686 31222 4738 31274
rect 4738 31222 4740 31274
rect 4684 31220 4740 31222
rect 6300 31724 6356 31780
rect 6076 30716 6132 30772
rect 6188 31388 6244 31444
rect 5516 30604 5572 30660
rect 4060 30492 4116 30548
rect 4620 30546 4676 30548
rect 4620 30494 4622 30546
rect 4622 30494 4674 30546
rect 4674 30494 4676 30546
rect 4620 30492 4676 30494
rect 4060 29986 4116 29988
rect 4060 29934 4062 29986
rect 4062 29934 4114 29986
rect 4114 29934 4116 29986
rect 4060 29932 4116 29934
rect 2380 28754 2436 28756
rect 2380 28702 2382 28754
rect 2382 28702 2434 28754
rect 2434 28702 2436 28754
rect 2380 28700 2436 28702
rect 1932 28476 1988 28532
rect 3164 28476 3220 28532
rect 1820 25954 1876 25956
rect 1820 25902 1822 25954
rect 1822 25902 1874 25954
rect 1874 25902 1876 25954
rect 1820 25900 1876 25902
rect 4956 29484 5012 29540
rect 4476 29258 4532 29260
rect 4476 29206 4478 29258
rect 4478 29206 4530 29258
rect 4530 29206 4532 29258
rect 4476 29204 4532 29206
rect 4580 29258 4636 29260
rect 4580 29206 4582 29258
rect 4582 29206 4634 29258
rect 4634 29206 4636 29258
rect 4580 29204 4636 29206
rect 4684 29258 4740 29260
rect 4684 29206 4686 29258
rect 4686 29206 4738 29258
rect 4738 29206 4740 29258
rect 4684 29204 4740 29206
rect 6860 33794 6916 33796
rect 6860 33742 6862 33794
rect 6862 33742 6914 33794
rect 6914 33742 6916 33794
rect 6860 33740 6916 33742
rect 7532 32284 7588 32340
rect 6972 31778 7028 31780
rect 6972 31726 6974 31778
rect 6974 31726 7026 31778
rect 7026 31726 7028 31778
rect 6972 31724 7028 31726
rect 7420 31778 7476 31780
rect 7420 31726 7422 31778
rect 7422 31726 7474 31778
rect 7474 31726 7476 31778
rect 7420 31724 7476 31726
rect 6860 31388 6916 31444
rect 7308 31442 7364 31444
rect 7308 31390 7310 31442
rect 7310 31390 7362 31442
rect 7362 31390 7364 31442
rect 7308 31388 7364 31390
rect 8876 32002 8932 32004
rect 8876 31950 8878 32002
rect 8878 31950 8930 32002
rect 8930 31950 8932 32002
rect 8876 31948 8932 31950
rect 10892 32562 10948 32564
rect 10892 32510 10894 32562
rect 10894 32510 10946 32562
rect 10946 32510 10948 32562
rect 10892 32508 10948 32510
rect 9772 31948 9828 32004
rect 12236 33570 12292 33572
rect 12236 33518 12238 33570
rect 12238 33518 12290 33570
rect 12290 33518 12292 33570
rect 12236 33516 12292 33518
rect 7532 31388 7588 31444
rect 8764 31724 8820 31780
rect 7308 30492 7364 30548
rect 9996 30940 10052 30996
rect 8316 30546 8372 30548
rect 8316 30494 8318 30546
rect 8318 30494 8370 30546
rect 8370 30494 8372 30546
rect 8316 30492 8372 30494
rect 5740 29484 5796 29540
rect 6188 28700 6244 28756
rect 4956 28642 5012 28644
rect 4956 28590 4958 28642
rect 4958 28590 5010 28642
rect 5010 28590 5012 28642
rect 4956 28588 5012 28590
rect 6076 28642 6132 28644
rect 6076 28590 6078 28642
rect 6078 28590 6130 28642
rect 6130 28590 6132 28642
rect 6076 28588 6132 28590
rect 6748 28700 6804 28756
rect 2716 26796 2772 26852
rect 5740 28476 5796 28532
rect 6748 27580 6804 27636
rect 4476 27242 4532 27244
rect 4476 27190 4478 27242
rect 4478 27190 4530 27242
rect 4530 27190 4532 27242
rect 4476 27188 4532 27190
rect 4580 27242 4636 27244
rect 4580 27190 4582 27242
rect 4582 27190 4634 27242
rect 4634 27190 4636 27242
rect 4580 27188 4636 27190
rect 4684 27242 4740 27244
rect 4684 27190 4686 27242
rect 4686 27190 4738 27242
rect 4738 27190 4740 27242
rect 4684 27188 4740 27190
rect 4956 26850 5012 26852
rect 4956 26798 4958 26850
rect 4958 26798 5010 26850
rect 5010 26798 5012 26850
rect 4956 26796 5012 26798
rect 9996 30044 10052 30100
rect 10556 30546 10612 30548
rect 10556 30494 10558 30546
rect 10558 30494 10610 30546
rect 10610 30494 10612 30546
rect 10556 30492 10612 30494
rect 11116 30492 11172 30548
rect 11676 30156 11732 30212
rect 14028 33516 14084 33572
rect 13580 32620 13636 32676
rect 13468 32562 13524 32564
rect 13468 32510 13470 32562
rect 13470 32510 13522 32562
rect 13522 32510 13524 32562
rect 13468 32508 13524 32510
rect 14140 32002 14196 32004
rect 14140 31950 14142 32002
rect 14142 31950 14194 32002
rect 14194 31950 14196 32002
rect 14140 31948 14196 31950
rect 12908 31836 12964 31892
rect 16380 35868 16436 35924
rect 16380 35698 16436 35700
rect 16380 35646 16382 35698
rect 16382 35646 16434 35698
rect 16434 35646 16436 35698
rect 16380 35644 16436 35646
rect 16828 35084 16884 35140
rect 16604 34690 16660 34692
rect 16604 34638 16606 34690
rect 16606 34638 16658 34690
rect 16658 34638 16660 34690
rect 16604 34636 16660 34638
rect 17612 38668 17668 38724
rect 18172 37100 18228 37156
rect 17724 35644 17780 35700
rect 16380 33906 16436 33908
rect 16380 33854 16382 33906
rect 16382 33854 16434 33906
rect 16434 33854 16436 33906
rect 16380 33852 16436 33854
rect 16380 33628 16436 33684
rect 13804 31890 13860 31892
rect 13804 31838 13806 31890
rect 13806 31838 13858 31890
rect 13858 31838 13860 31890
rect 13804 31836 13860 31838
rect 12908 30828 12964 30884
rect 12460 30770 12516 30772
rect 12460 30718 12462 30770
rect 12462 30718 12514 30770
rect 12514 30718 12516 30770
rect 12460 30716 12516 30718
rect 12124 30546 12180 30548
rect 12124 30494 12126 30546
rect 12126 30494 12178 30546
rect 12178 30494 12180 30546
rect 12124 30492 12180 30494
rect 15372 31890 15428 31892
rect 15372 31838 15374 31890
rect 15374 31838 15426 31890
rect 15426 31838 15428 31890
rect 15372 31836 15428 31838
rect 14364 31666 14420 31668
rect 14364 31614 14366 31666
rect 14366 31614 14418 31666
rect 14418 31614 14420 31666
rect 14364 31612 14420 31614
rect 13244 30492 13300 30548
rect 12124 30098 12180 30100
rect 12124 30046 12126 30098
rect 12126 30046 12178 30098
rect 12178 30046 12180 30098
rect 12124 30044 12180 30046
rect 11564 29820 11620 29876
rect 12572 29874 12628 29876
rect 12572 29822 12574 29874
rect 12574 29822 12626 29874
rect 12626 29822 12628 29874
rect 12572 29820 12628 29822
rect 14028 30492 14084 30548
rect 14924 30882 14980 30884
rect 14924 30830 14926 30882
rect 14926 30830 14978 30882
rect 14978 30830 14980 30882
rect 14924 30828 14980 30830
rect 14140 30268 14196 30324
rect 13132 29148 13188 29204
rect 12908 29036 12964 29092
rect 12460 28588 12516 28644
rect 13468 28642 13524 28644
rect 13468 28590 13470 28642
rect 13470 28590 13522 28642
rect 13522 28590 13524 28642
rect 13468 28588 13524 28590
rect 13692 28588 13748 28644
rect 8316 26796 8372 26852
rect 9324 26850 9380 26852
rect 9324 26798 9326 26850
rect 9326 26798 9378 26850
rect 9378 26798 9380 26850
rect 9324 26796 9380 26798
rect 2716 25954 2772 25956
rect 2716 25902 2718 25954
rect 2718 25902 2770 25954
rect 2770 25902 2772 25954
rect 2716 25900 2772 25902
rect 2268 25564 2324 25620
rect 1820 25340 1876 25396
rect 1820 23938 1876 23940
rect 1820 23886 1822 23938
rect 1822 23886 1874 23938
rect 1874 23886 1876 23938
rect 1820 23884 1876 23886
rect 1932 23548 1988 23604
rect 2604 23938 2660 23940
rect 2604 23886 2606 23938
rect 2606 23886 2658 23938
rect 2658 23886 2660 23938
rect 2604 23884 2660 23886
rect 3500 25394 3556 25396
rect 3500 25342 3502 25394
rect 3502 25342 3554 25394
rect 3554 25342 3556 25394
rect 3500 25340 3556 25342
rect 3948 25618 4004 25620
rect 3948 25566 3950 25618
rect 3950 25566 4002 25618
rect 4002 25566 4004 25618
rect 3948 25564 4004 25566
rect 4476 25226 4532 25228
rect 4476 25174 4478 25226
rect 4478 25174 4530 25226
rect 4530 25174 4532 25226
rect 4476 25172 4532 25174
rect 4580 25226 4636 25228
rect 4580 25174 4582 25226
rect 4582 25174 4634 25226
rect 4634 25174 4636 25226
rect 4580 25172 4636 25174
rect 4684 25226 4740 25228
rect 4684 25174 4686 25226
rect 4686 25174 4738 25226
rect 4738 25174 4740 25226
rect 4684 25172 4740 25174
rect 4844 24668 4900 24724
rect 5740 25676 5796 25732
rect 7196 25730 7252 25732
rect 7196 25678 7198 25730
rect 7198 25678 7250 25730
rect 7250 25678 7252 25730
rect 7196 25676 7252 25678
rect 6188 25564 6244 25620
rect 5068 24444 5124 24500
rect 3164 23548 3220 23604
rect 4844 23548 4900 23604
rect 4476 23210 4532 23212
rect 4476 23158 4478 23210
rect 4478 23158 4530 23210
rect 4530 23158 4532 23210
rect 4476 23156 4532 23158
rect 4580 23210 4636 23212
rect 4580 23158 4582 23210
rect 4582 23158 4634 23210
rect 4634 23158 4636 23210
rect 4580 23156 4636 23158
rect 4684 23210 4740 23212
rect 4684 23158 4686 23210
rect 4686 23158 4738 23210
rect 4738 23158 4740 23210
rect 4684 23156 4740 23158
rect 5852 25228 5908 25284
rect 5628 24722 5684 24724
rect 5628 24670 5630 24722
rect 5630 24670 5682 24722
rect 5682 24670 5684 24722
rect 5628 24668 5684 24670
rect 6188 24444 6244 24500
rect 6524 24498 6580 24500
rect 6524 24446 6526 24498
rect 6526 24446 6578 24498
rect 6578 24446 6580 24498
rect 6524 24444 6580 24446
rect 4620 22764 4676 22820
rect 8764 25730 8820 25732
rect 8764 25678 8766 25730
rect 8766 25678 8818 25730
rect 8818 25678 8820 25730
rect 8764 25676 8820 25678
rect 8204 25228 8260 25284
rect 9324 24722 9380 24724
rect 9324 24670 9326 24722
rect 9326 24670 9378 24722
rect 9378 24670 9380 24722
rect 9324 24668 9380 24670
rect 10108 26796 10164 26852
rect 9772 26626 9828 26628
rect 9772 26574 9774 26626
rect 9774 26574 9826 26626
rect 9826 26574 9828 26626
rect 9772 26572 9828 26574
rect 11228 26796 11284 26852
rect 11452 26572 11508 26628
rect 11004 26348 11060 26404
rect 14028 28754 14084 28756
rect 14028 28702 14030 28754
rect 14030 28702 14082 28754
rect 14082 28702 14084 28754
rect 14028 28700 14084 28702
rect 13916 28252 13972 28308
rect 12796 26796 12852 26852
rect 9660 25340 9716 25396
rect 10220 24722 10276 24724
rect 10220 24670 10222 24722
rect 10222 24670 10274 24722
rect 10274 24670 10276 24722
rect 10220 24668 10276 24670
rect 11340 25394 11396 25396
rect 11340 25342 11342 25394
rect 11342 25342 11394 25394
rect 11394 25342 11396 25394
rect 11340 25340 11396 25342
rect 13468 26796 13524 26852
rect 12908 26738 12964 26740
rect 12908 26686 12910 26738
rect 12910 26686 12962 26738
rect 12962 26686 12964 26738
rect 12908 26684 12964 26686
rect 12796 26348 12852 26404
rect 12124 25340 12180 25396
rect 14028 26738 14084 26740
rect 14028 26686 14030 26738
rect 14030 26686 14082 26738
rect 14082 26686 14084 26738
rect 14028 26684 14084 26686
rect 14252 26684 14308 26740
rect 13580 26460 13636 26516
rect 10892 24668 10948 24724
rect 14700 30492 14756 30548
rect 15036 30044 15092 30100
rect 14924 29874 14980 29876
rect 14924 29822 14926 29874
rect 14926 29822 14978 29874
rect 14978 29822 14980 29874
rect 14924 29820 14980 29822
rect 16940 32956 16996 33012
rect 15708 31724 15764 31780
rect 16380 31778 16436 31780
rect 16380 31726 16382 31778
rect 16382 31726 16434 31778
rect 16434 31726 16436 31778
rect 16380 31724 16436 31726
rect 16268 30380 16324 30436
rect 15932 30044 15988 30100
rect 14924 29036 14980 29092
rect 14700 28588 14756 28644
rect 14476 26572 14532 26628
rect 14364 26348 14420 26404
rect 9548 24444 9604 24500
rect 12348 24498 12404 24500
rect 12348 24446 12350 24498
rect 12350 24446 12402 24498
rect 12402 24446 12404 24498
rect 12348 24444 12404 24446
rect 14028 24498 14084 24500
rect 14028 24446 14030 24498
rect 14030 24446 14082 24498
rect 14082 24446 14084 24498
rect 14028 24444 14084 24446
rect 15484 29596 15540 29652
rect 16380 29762 16436 29764
rect 16380 29710 16382 29762
rect 16382 29710 16434 29762
rect 16434 29710 16436 29762
rect 16380 29708 16436 29710
rect 16940 28978 16996 28980
rect 16940 28926 16942 28978
rect 16942 28926 16994 28978
rect 16994 28926 16996 28978
rect 16940 28924 16996 28926
rect 16604 28866 16660 28868
rect 16604 28814 16606 28866
rect 16606 28814 16658 28866
rect 16658 28814 16660 28866
rect 16604 28812 16660 28814
rect 15036 28700 15092 28756
rect 15036 26908 15092 26964
rect 15932 28642 15988 28644
rect 15932 28590 15934 28642
rect 15934 28590 15986 28642
rect 15986 28590 15988 28642
rect 15932 28588 15988 28590
rect 16492 28642 16548 28644
rect 16492 28590 16494 28642
rect 16494 28590 16546 28642
rect 16546 28590 16548 28642
rect 16492 28588 16548 28590
rect 16044 27858 16100 27860
rect 16044 27806 16046 27858
rect 16046 27806 16098 27858
rect 16098 27806 16100 27858
rect 16044 27804 16100 27806
rect 15484 26460 15540 26516
rect 16156 26684 16212 26740
rect 16604 26514 16660 26516
rect 16604 26462 16606 26514
rect 16606 26462 16658 26514
rect 16658 26462 16660 26514
rect 16604 26460 16660 26462
rect 16828 25618 16884 25620
rect 16828 25566 16830 25618
rect 16830 25566 16882 25618
rect 16882 25566 16884 25618
rect 16828 25564 16884 25566
rect 16268 24722 16324 24724
rect 16268 24670 16270 24722
rect 16270 24670 16322 24722
rect 16322 24670 16324 24722
rect 16268 24668 16324 24670
rect 14588 24444 14644 24500
rect 16828 23602 16884 23604
rect 16828 23550 16830 23602
rect 16830 23550 16882 23602
rect 16882 23550 16884 23602
rect 16828 23548 16884 23550
rect 5740 22818 5796 22820
rect 5740 22766 5742 22818
rect 5742 22766 5794 22818
rect 5794 22766 5796 22818
rect 5740 22764 5796 22766
rect 15260 22370 15316 22372
rect 15260 22318 15262 22370
rect 15262 22318 15314 22370
rect 15314 22318 15316 22370
rect 15260 22316 15316 22318
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 16940 21868 16996 21924
rect 16268 20748 16324 20804
rect 14700 20188 14756 20244
rect 15260 20188 15316 20244
rect 16940 20802 16996 20804
rect 16940 20750 16942 20802
rect 16942 20750 16994 20802
rect 16994 20750 16996 20802
rect 16940 20748 16996 20750
rect 16828 20188 16884 20244
rect 4476 19178 4532 19180
rect 4476 19126 4478 19178
rect 4478 19126 4530 19178
rect 4530 19126 4532 19178
rect 4476 19124 4532 19126
rect 4580 19178 4636 19180
rect 4580 19126 4582 19178
rect 4582 19126 4634 19178
rect 4634 19126 4636 19178
rect 4580 19124 4636 19126
rect 4684 19178 4740 19180
rect 4684 19126 4686 19178
rect 4686 19126 4738 19178
rect 4738 19126 4740 19178
rect 4684 19124 4740 19126
rect 16716 19906 16772 19908
rect 16716 19854 16718 19906
rect 16718 19854 16770 19906
rect 16770 19854 16772 19906
rect 16716 19852 16772 19854
rect 17388 31778 17444 31780
rect 17388 31726 17390 31778
rect 17390 31726 17442 31778
rect 17442 31726 17444 31778
rect 17388 31724 17444 31726
rect 17388 29596 17444 29652
rect 17388 29036 17444 29092
rect 19292 40850 19348 40852
rect 19292 40798 19294 40850
rect 19294 40798 19346 40850
rect 19346 40798 19348 40850
rect 19292 40796 19348 40798
rect 19836 40346 19892 40348
rect 19836 40294 19838 40346
rect 19838 40294 19890 40346
rect 19890 40294 19892 40346
rect 19836 40292 19892 40294
rect 19940 40346 19996 40348
rect 19940 40294 19942 40346
rect 19942 40294 19994 40346
rect 19994 40294 19996 40346
rect 19940 40292 19996 40294
rect 20044 40346 20100 40348
rect 20044 40294 20046 40346
rect 20046 40294 20098 40346
rect 20098 40294 20100 40346
rect 20044 40292 20100 40294
rect 21756 44604 21812 44660
rect 22428 46898 22484 46900
rect 22428 46846 22430 46898
rect 22430 46846 22482 46898
rect 22482 46846 22484 46898
rect 22428 46844 22484 46846
rect 22876 46956 22932 47012
rect 23660 47068 23716 47124
rect 23548 46956 23604 47012
rect 23996 46844 24052 46900
rect 22652 46114 22708 46116
rect 22652 46062 22654 46114
rect 22654 46062 22706 46114
rect 22706 46062 22708 46114
rect 22652 46060 22708 46062
rect 23324 46114 23380 46116
rect 23324 46062 23326 46114
rect 23326 46062 23378 46114
rect 23378 46062 23380 46114
rect 23324 46060 23380 46062
rect 23772 44604 23828 44660
rect 20636 42812 20692 42868
rect 21532 43708 21588 43764
rect 20412 41692 20468 41748
rect 20300 40796 20356 40852
rect 20412 41020 20468 41076
rect 20188 40012 20244 40068
rect 19852 38668 19908 38724
rect 18732 36594 18788 36596
rect 18732 36542 18734 36594
rect 18734 36542 18786 36594
rect 18786 36542 18788 36594
rect 18732 36540 18788 36542
rect 21644 41970 21700 41972
rect 21644 41918 21646 41970
rect 21646 41918 21698 41970
rect 21698 41918 21700 41970
rect 21644 41916 21700 41918
rect 23436 43596 23492 43652
rect 23100 42866 23156 42868
rect 23100 42814 23102 42866
rect 23102 42814 23154 42866
rect 23154 42814 23156 42866
rect 23100 42812 23156 42814
rect 24332 48802 24388 48804
rect 24332 48750 24334 48802
rect 24334 48750 24386 48802
rect 24386 48750 24388 48802
rect 24332 48748 24388 48750
rect 25228 48802 25284 48804
rect 25228 48750 25230 48802
rect 25230 48750 25282 48802
rect 25282 48750 25284 48802
rect 25228 48748 25284 48750
rect 24220 46844 24276 46900
rect 24220 46114 24276 46116
rect 24220 46062 24222 46114
rect 24222 46062 24274 46114
rect 24274 46062 24276 46114
rect 24220 46060 24276 46062
rect 24108 43596 24164 43652
rect 21980 42140 22036 42196
rect 21868 41804 21924 41860
rect 20748 41580 20804 41636
rect 21980 41692 22036 41748
rect 21308 40796 21364 40852
rect 20748 40738 20804 40740
rect 20748 40686 20750 40738
rect 20750 40686 20802 40738
rect 20802 40686 20804 40738
rect 20748 40684 20804 40686
rect 20860 39954 20916 39956
rect 20860 39902 20862 39954
rect 20862 39902 20914 39954
rect 20914 39902 20916 39954
rect 20860 39900 20916 39902
rect 22092 41916 22148 41972
rect 22764 42140 22820 42196
rect 24108 41916 24164 41972
rect 22092 41020 22148 41076
rect 22316 41804 22372 41860
rect 22764 41580 22820 41636
rect 23884 41634 23940 41636
rect 23884 41582 23886 41634
rect 23886 41582 23938 41634
rect 23938 41582 23940 41634
rect 23884 41580 23940 41582
rect 22316 40738 22372 40740
rect 22316 40686 22318 40738
rect 22318 40686 22370 40738
rect 22370 40686 22372 40738
rect 22316 40684 22372 40686
rect 24332 43820 24388 43876
rect 31948 48748 32004 48804
rect 26012 48018 26068 48020
rect 26012 47966 26014 48018
rect 26014 47966 26066 48018
rect 26066 47966 26068 48018
rect 26012 47964 26068 47966
rect 26908 46956 26964 47012
rect 24556 46172 24612 46228
rect 25116 46172 25172 46228
rect 26460 46172 26516 46228
rect 25452 46114 25508 46116
rect 25452 46062 25454 46114
rect 25454 46062 25506 46114
rect 25506 46062 25508 46114
rect 25452 46060 25508 46062
rect 25228 45724 25284 45780
rect 24220 40796 24276 40852
rect 21644 40012 21700 40068
rect 24108 40236 24164 40292
rect 21532 39900 21588 39956
rect 22540 39954 22596 39956
rect 22540 39902 22542 39954
rect 22542 39902 22594 39954
rect 22594 39902 22596 39954
rect 22540 39900 22596 39902
rect 20188 38556 20244 38612
rect 19836 38330 19892 38332
rect 19836 38278 19838 38330
rect 19838 38278 19890 38330
rect 19890 38278 19892 38330
rect 19836 38276 19892 38278
rect 19940 38330 19996 38332
rect 19940 38278 19942 38330
rect 19942 38278 19994 38330
rect 19994 38278 19996 38330
rect 19940 38276 19996 38278
rect 20044 38330 20100 38332
rect 20044 38278 20046 38330
rect 20046 38278 20098 38330
rect 20098 38278 20100 38330
rect 20044 38276 20100 38278
rect 20188 37100 20244 37156
rect 20636 38556 20692 38612
rect 20860 38556 20916 38612
rect 20188 36930 20244 36932
rect 20188 36878 20190 36930
rect 20190 36878 20242 36930
rect 20242 36878 20244 36930
rect 20188 36876 20244 36878
rect 19516 36652 19572 36708
rect 20748 36764 20804 36820
rect 18396 36092 18452 36148
rect 18620 35644 18676 35700
rect 19836 36314 19892 36316
rect 19836 36262 19838 36314
rect 19838 36262 19890 36314
rect 19890 36262 19892 36314
rect 19836 36260 19892 36262
rect 19940 36314 19996 36316
rect 19940 36262 19942 36314
rect 19942 36262 19994 36314
rect 19994 36262 19996 36314
rect 19940 36260 19996 36262
rect 20044 36314 20100 36316
rect 20044 36262 20046 36314
rect 20046 36262 20098 36314
rect 20098 36262 20100 36314
rect 20044 36260 20100 36262
rect 19180 36146 19236 36148
rect 19180 36094 19182 36146
rect 19182 36094 19234 36146
rect 19234 36094 19236 36146
rect 19180 36092 19236 36094
rect 19628 36092 19684 36148
rect 18844 35980 18900 36036
rect 20636 36092 20692 36148
rect 23660 38780 23716 38836
rect 23772 40012 23828 40068
rect 21644 37996 21700 38052
rect 23100 38050 23156 38052
rect 23100 37998 23102 38050
rect 23102 37998 23154 38050
rect 23154 37998 23156 38050
rect 23100 37996 23156 37998
rect 23772 38050 23828 38052
rect 23772 37998 23774 38050
rect 23774 37998 23826 38050
rect 23826 37998 23828 38050
rect 23772 37996 23828 37998
rect 20860 36652 20916 36708
rect 21196 36594 21252 36596
rect 21196 36542 21198 36594
rect 21198 36542 21250 36594
rect 21250 36542 21252 36594
rect 21196 36540 21252 36542
rect 19852 35980 19908 36036
rect 18172 33852 18228 33908
rect 18844 33906 18900 33908
rect 18844 33854 18846 33906
rect 18846 33854 18898 33906
rect 18898 33854 18900 33906
rect 18844 33852 18900 33854
rect 17948 33628 18004 33684
rect 19180 33740 19236 33796
rect 18956 33682 19012 33684
rect 18956 33630 18958 33682
rect 18958 33630 19010 33682
rect 19010 33630 19012 33682
rect 18956 33628 19012 33630
rect 17724 31948 17780 32004
rect 17612 28924 17668 28980
rect 19068 31612 19124 31668
rect 18620 30770 18676 30772
rect 18620 30718 18622 30770
rect 18622 30718 18674 30770
rect 18674 30718 18676 30770
rect 18620 30716 18676 30718
rect 18060 29650 18116 29652
rect 18060 29598 18062 29650
rect 18062 29598 18114 29650
rect 18114 29598 18116 29650
rect 18060 29596 18116 29598
rect 17724 28812 17780 28868
rect 18396 28700 18452 28756
rect 18508 28924 18564 28980
rect 17948 28028 18004 28084
rect 18956 28364 19012 28420
rect 18956 27858 19012 27860
rect 18956 27806 18958 27858
rect 18958 27806 19010 27858
rect 19010 27806 19012 27858
rect 18956 27804 19012 27806
rect 17500 24668 17556 24724
rect 17836 25564 17892 25620
rect 17612 24780 17668 24836
rect 17948 24668 18004 24724
rect 17500 23660 17556 23716
rect 19180 29148 19236 29204
rect 19180 28476 19236 28532
rect 19068 24722 19124 24724
rect 19068 24670 19070 24722
rect 19070 24670 19122 24722
rect 19122 24670 19124 24722
rect 19068 24668 19124 24670
rect 19068 23884 19124 23940
rect 18844 23714 18900 23716
rect 18844 23662 18846 23714
rect 18846 23662 18898 23714
rect 18898 23662 18900 23714
rect 18844 23660 18900 23662
rect 18396 23548 18452 23604
rect 18396 22540 18452 22596
rect 17948 21868 18004 21924
rect 18284 21922 18340 21924
rect 18284 21870 18286 21922
rect 18286 21870 18338 21922
rect 18338 21870 18340 21922
rect 18284 21868 18340 21870
rect 18620 21810 18676 21812
rect 18620 21758 18622 21810
rect 18622 21758 18674 21810
rect 18674 21758 18676 21810
rect 18620 21756 18676 21758
rect 17948 21420 18004 21476
rect 4476 17162 4532 17164
rect 4476 17110 4478 17162
rect 4478 17110 4530 17162
rect 4530 17110 4532 17162
rect 4476 17108 4532 17110
rect 4580 17162 4636 17164
rect 4580 17110 4582 17162
rect 4582 17110 4634 17162
rect 4634 17110 4636 17162
rect 4580 17108 4636 17110
rect 4684 17162 4740 17164
rect 4684 17110 4686 17162
rect 4686 17110 4738 17162
rect 4738 17110 4740 17162
rect 4684 17108 4740 17110
rect 4476 15146 4532 15148
rect 4476 15094 4478 15146
rect 4478 15094 4530 15146
rect 4530 15094 4532 15146
rect 4476 15092 4532 15094
rect 4580 15146 4636 15148
rect 4580 15094 4582 15146
rect 4582 15094 4634 15146
rect 4634 15094 4636 15146
rect 4580 15092 4636 15094
rect 4684 15146 4740 15148
rect 4684 15094 4686 15146
rect 4686 15094 4738 15146
rect 4738 15094 4740 15146
rect 4684 15092 4740 15094
rect 18172 19852 18228 19908
rect 19180 21756 19236 21812
rect 19180 20412 19236 20468
rect 18620 19346 18676 19348
rect 18620 19294 18622 19346
rect 18622 19294 18674 19346
rect 18674 19294 18676 19346
rect 18620 19292 18676 19294
rect 17724 15650 17780 15652
rect 17724 15598 17726 15650
rect 17726 15598 17778 15650
rect 17778 15598 17780 15650
rect 17724 15596 17780 15598
rect 20748 35980 20804 36036
rect 20188 35084 20244 35140
rect 19628 34690 19684 34692
rect 19628 34638 19630 34690
rect 19630 34638 19682 34690
rect 19682 34638 19684 34690
rect 19628 34636 19684 34638
rect 19836 34298 19892 34300
rect 19836 34246 19838 34298
rect 19838 34246 19890 34298
rect 19890 34246 19892 34298
rect 19836 34244 19892 34246
rect 19940 34298 19996 34300
rect 19940 34246 19942 34298
rect 19942 34246 19994 34298
rect 19994 34246 19996 34298
rect 19940 34244 19996 34246
rect 20044 34298 20100 34300
rect 20044 34246 20046 34298
rect 20046 34246 20098 34298
rect 20098 34246 20100 34298
rect 20044 34244 20100 34246
rect 21420 35644 21476 35700
rect 21644 36876 21700 36932
rect 21868 36818 21924 36820
rect 21868 36766 21870 36818
rect 21870 36766 21922 36818
rect 21922 36766 21924 36818
rect 21868 36764 21924 36766
rect 23100 36930 23156 36932
rect 23100 36878 23102 36930
rect 23102 36878 23154 36930
rect 23154 36878 23156 36930
rect 23100 36876 23156 36878
rect 24220 37714 24276 37716
rect 24220 37662 24222 37714
rect 24222 37662 24274 37714
rect 24274 37662 24276 37714
rect 24220 37660 24276 37662
rect 24220 36930 24276 36932
rect 24220 36878 24222 36930
rect 24222 36878 24274 36930
rect 24274 36878 24276 36930
rect 24220 36876 24276 36878
rect 21868 36540 21924 36596
rect 20412 34802 20468 34804
rect 20412 34750 20414 34802
rect 20414 34750 20466 34802
rect 20466 34750 20468 34802
rect 20412 34748 20468 34750
rect 20188 33964 20244 34020
rect 20188 33794 20244 33796
rect 20188 33742 20190 33794
rect 20190 33742 20242 33794
rect 20242 33742 20244 33794
rect 20188 33740 20244 33742
rect 19740 33628 19796 33684
rect 19516 32956 19572 33012
rect 19836 32282 19892 32284
rect 19836 32230 19838 32282
rect 19838 32230 19890 32282
rect 19890 32230 19892 32282
rect 19836 32228 19892 32230
rect 19940 32282 19996 32284
rect 19940 32230 19942 32282
rect 19942 32230 19994 32282
rect 19994 32230 19996 32282
rect 19940 32228 19996 32230
rect 20044 32282 20100 32284
rect 20044 32230 20046 32282
rect 20046 32230 20098 32282
rect 20098 32230 20100 32282
rect 20044 32228 20100 32230
rect 20300 32674 20356 32676
rect 20300 32622 20302 32674
rect 20302 32622 20354 32674
rect 20354 32622 20356 32674
rect 20300 32620 20356 32622
rect 21308 34636 21364 34692
rect 20860 34018 20916 34020
rect 20860 33966 20862 34018
rect 20862 33966 20914 34018
rect 20914 33966 20916 34018
rect 20860 33964 20916 33966
rect 20972 33906 21028 33908
rect 20972 33854 20974 33906
rect 20974 33854 21026 33906
rect 21026 33854 21028 33906
rect 20972 33852 21028 33854
rect 21532 34802 21588 34804
rect 21532 34750 21534 34802
rect 21534 34750 21586 34802
rect 21586 34750 21588 34802
rect 21532 34748 21588 34750
rect 21644 34860 21700 34916
rect 21980 34860 22036 34916
rect 21756 33964 21812 34020
rect 21420 33628 21476 33684
rect 20636 32786 20692 32788
rect 20636 32734 20638 32786
rect 20638 32734 20690 32786
rect 20690 32734 20692 32786
rect 20636 32732 20692 32734
rect 20188 31948 20244 32004
rect 19516 31836 19572 31892
rect 20188 31666 20244 31668
rect 20188 31614 20190 31666
rect 20190 31614 20242 31666
rect 20242 31614 20244 31666
rect 20188 31612 20244 31614
rect 20412 30546 20468 30548
rect 20412 30494 20414 30546
rect 20414 30494 20466 30546
rect 20466 30494 20468 30546
rect 20412 30492 20468 30494
rect 19836 30266 19892 30268
rect 19836 30214 19838 30266
rect 19838 30214 19890 30266
rect 19890 30214 19892 30266
rect 19836 30212 19892 30214
rect 19940 30266 19996 30268
rect 19940 30214 19942 30266
rect 19942 30214 19994 30266
rect 19994 30214 19996 30266
rect 19940 30212 19996 30214
rect 20044 30266 20100 30268
rect 20044 30214 20046 30266
rect 20046 30214 20098 30266
rect 20098 30214 20100 30266
rect 20044 30212 20100 30214
rect 19628 30044 19684 30100
rect 19628 29148 19684 29204
rect 19516 28700 19572 28756
rect 19404 28028 19460 28084
rect 19852 28924 19908 28980
rect 21644 33570 21700 33572
rect 21644 33518 21646 33570
rect 21646 33518 21698 33570
rect 21698 33518 21700 33570
rect 21644 33516 21700 33518
rect 23548 36594 23604 36596
rect 23548 36542 23550 36594
rect 23550 36542 23602 36594
rect 23602 36542 23604 36594
rect 23548 36540 23604 36542
rect 23996 36540 24052 36596
rect 22876 34802 22932 34804
rect 22876 34750 22878 34802
rect 22878 34750 22930 34802
rect 22930 34750 22932 34802
rect 22876 34748 22932 34750
rect 23324 34802 23380 34804
rect 23324 34750 23326 34802
rect 23326 34750 23378 34802
rect 23378 34750 23380 34802
rect 23324 34748 23380 34750
rect 22428 34690 22484 34692
rect 22428 34638 22430 34690
rect 22430 34638 22482 34690
rect 22482 34638 22484 34690
rect 22428 34636 22484 34638
rect 22316 34300 22372 34356
rect 23212 34076 23268 34132
rect 22652 33906 22708 33908
rect 22652 33854 22654 33906
rect 22654 33854 22706 33906
rect 22706 33854 22708 33906
rect 22652 33852 22708 33854
rect 22092 32956 22148 33012
rect 22204 32732 22260 32788
rect 23772 34690 23828 34692
rect 23772 34638 23774 34690
rect 23774 34638 23826 34690
rect 23826 34638 23828 34690
rect 23772 34636 23828 34638
rect 23660 33852 23716 33908
rect 22428 32508 22484 32564
rect 22876 31836 22932 31892
rect 21308 31388 21364 31444
rect 22204 31388 22260 31444
rect 23548 33628 23604 33684
rect 24556 43596 24612 43652
rect 24668 43372 24724 43428
rect 25676 43708 25732 43764
rect 28140 47964 28196 48020
rect 27356 46172 27412 46228
rect 27020 43820 27076 43876
rect 25116 41804 25172 41860
rect 24556 40236 24612 40292
rect 24668 41746 24724 41748
rect 24668 41694 24670 41746
rect 24670 41694 24722 41746
rect 24722 41694 24724 41746
rect 24668 41692 24724 41694
rect 24668 39900 24724 39956
rect 24444 39676 24500 39732
rect 24780 40348 24836 40404
rect 26124 43762 26180 43764
rect 26124 43710 26126 43762
rect 26126 43710 26178 43762
rect 26178 43710 26180 43762
rect 26124 43708 26180 43710
rect 27244 45724 27300 45780
rect 27692 46172 27748 46228
rect 28476 48018 28532 48020
rect 28476 47966 28478 48018
rect 28478 47966 28530 48018
rect 28530 47966 28532 48018
rect 28476 47964 28532 47966
rect 28588 46844 28644 46900
rect 29372 46898 29428 46900
rect 29372 46846 29374 46898
rect 29374 46846 29426 46898
rect 29426 46846 29428 46898
rect 29372 46844 29428 46846
rect 28252 46732 28308 46788
rect 29820 46732 29876 46788
rect 30604 46172 30660 46228
rect 27804 44604 27860 44660
rect 32060 46956 32116 47012
rect 32060 46620 32116 46676
rect 32284 46226 32340 46228
rect 32284 46174 32286 46226
rect 32286 46174 32338 46226
rect 32338 46174 32340 46226
rect 32284 46172 32340 46174
rect 31052 45948 31108 46004
rect 31948 46060 32004 46116
rect 31500 45890 31556 45892
rect 31500 45838 31502 45890
rect 31502 45838 31554 45890
rect 31554 45838 31556 45890
rect 31500 45836 31556 45838
rect 27244 43596 27300 43652
rect 27244 42978 27300 42980
rect 27244 42926 27246 42978
rect 27246 42926 27298 42978
rect 27298 42926 27300 42978
rect 27244 42924 27300 42926
rect 28028 42812 28084 42868
rect 26796 42140 26852 42196
rect 27468 41970 27524 41972
rect 27468 41918 27470 41970
rect 27470 41918 27522 41970
rect 27522 41918 27524 41970
rect 27468 41916 27524 41918
rect 25676 41692 25732 41748
rect 27132 41804 27188 41860
rect 26796 41692 26852 41748
rect 25564 41580 25620 41636
rect 25452 41020 25508 41076
rect 25788 40850 25844 40852
rect 25788 40798 25790 40850
rect 25790 40798 25842 40850
rect 25842 40798 25844 40850
rect 25788 40796 25844 40798
rect 26348 39954 26404 39956
rect 26348 39902 26350 39954
rect 26350 39902 26402 39954
rect 26402 39902 26404 39954
rect 26348 39900 26404 39902
rect 25452 39730 25508 39732
rect 25452 39678 25454 39730
rect 25454 39678 25506 39730
rect 25506 39678 25508 39730
rect 25452 39676 25508 39678
rect 25900 38834 25956 38836
rect 25900 38782 25902 38834
rect 25902 38782 25954 38834
rect 25954 38782 25956 38834
rect 25900 38780 25956 38782
rect 25340 38722 25396 38724
rect 25340 38670 25342 38722
rect 25342 38670 25394 38722
rect 25394 38670 25396 38722
rect 25340 38668 25396 38670
rect 25228 37996 25284 38052
rect 24444 36652 24500 36708
rect 25564 37660 25620 37716
rect 26012 36706 26068 36708
rect 26012 36654 26014 36706
rect 26014 36654 26066 36706
rect 26066 36654 26068 36706
rect 26012 36652 26068 36654
rect 24668 36540 24724 36596
rect 25900 36540 25956 36596
rect 26460 36428 26516 36484
rect 24556 35810 24612 35812
rect 24556 35758 24558 35810
rect 24558 35758 24610 35810
rect 24610 35758 24612 35810
rect 24556 35756 24612 35758
rect 26348 35756 26404 35812
rect 24668 34578 24724 34580
rect 24668 34526 24670 34578
rect 24670 34526 24722 34578
rect 24722 34526 24724 34578
rect 24668 34524 24724 34526
rect 24108 34076 24164 34132
rect 24108 33628 24164 33684
rect 24332 32786 24388 32788
rect 24332 32734 24334 32786
rect 24334 32734 24386 32786
rect 24386 32734 24388 32786
rect 24332 32732 24388 32734
rect 24668 34076 24724 34132
rect 25676 35196 25732 35252
rect 24892 33964 24948 34020
rect 25116 33628 25172 33684
rect 22988 31388 23044 31444
rect 21420 30492 21476 30548
rect 21420 30098 21476 30100
rect 21420 30046 21422 30098
rect 21422 30046 21474 30098
rect 21474 30046 21476 30098
rect 21420 30044 21476 30046
rect 21084 29596 21140 29652
rect 21196 29708 21252 29764
rect 20636 28978 20692 28980
rect 20636 28926 20638 28978
rect 20638 28926 20690 28978
rect 20690 28926 20692 28978
rect 20636 28924 20692 28926
rect 21196 29036 21252 29092
rect 20300 28754 20356 28756
rect 20300 28702 20302 28754
rect 20302 28702 20354 28754
rect 20354 28702 20356 28754
rect 20300 28700 20356 28702
rect 21868 29874 21924 29876
rect 21868 29822 21870 29874
rect 21870 29822 21922 29874
rect 21922 29822 21924 29874
rect 21868 29820 21924 29822
rect 21756 29372 21812 29428
rect 21532 28924 21588 28980
rect 22092 28924 22148 28980
rect 22316 28812 22372 28868
rect 23100 29762 23156 29764
rect 23100 29710 23102 29762
rect 23102 29710 23154 29762
rect 23154 29710 23156 29762
rect 23100 29708 23156 29710
rect 22988 28700 23044 28756
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 22316 28252 22372 28308
rect 20044 28196 20100 28198
rect 19516 27356 19572 27412
rect 22204 26572 22260 26628
rect 19836 26234 19892 26236
rect 19836 26182 19838 26234
rect 19838 26182 19890 26234
rect 19890 26182 19892 26234
rect 19836 26180 19892 26182
rect 19940 26234 19996 26236
rect 19940 26182 19942 26234
rect 19942 26182 19994 26234
rect 19994 26182 19996 26234
rect 19940 26180 19996 26182
rect 20044 26234 20100 26236
rect 20044 26182 20046 26234
rect 20046 26182 20098 26234
rect 20098 26182 20100 26234
rect 20044 26180 20100 26182
rect 19964 25730 20020 25732
rect 19964 25678 19966 25730
rect 19966 25678 20018 25730
rect 20018 25678 20020 25730
rect 19964 25676 20020 25678
rect 20524 25228 20580 25284
rect 19404 24834 19460 24836
rect 19404 24782 19406 24834
rect 19406 24782 19458 24834
rect 19458 24782 19460 24834
rect 19404 24780 19460 24782
rect 19964 24780 20020 24836
rect 19836 24218 19892 24220
rect 19836 24166 19838 24218
rect 19838 24166 19890 24218
rect 19890 24166 19892 24218
rect 19836 24164 19892 24166
rect 19940 24218 19996 24220
rect 19940 24166 19942 24218
rect 19942 24166 19994 24218
rect 19994 24166 19996 24218
rect 19940 24164 19996 24166
rect 20044 24218 20100 24220
rect 20044 24166 20046 24218
rect 20046 24166 20098 24218
rect 20098 24166 20100 24218
rect 20044 24164 20100 24166
rect 20300 23660 20356 23716
rect 20188 22540 20244 22596
rect 19836 22202 19892 22204
rect 19836 22150 19838 22202
rect 19838 22150 19890 22202
rect 19890 22150 19892 22202
rect 19836 22148 19892 22150
rect 19940 22202 19996 22204
rect 19940 22150 19942 22202
rect 19942 22150 19994 22202
rect 19994 22150 19996 22202
rect 19940 22148 19996 22150
rect 20044 22202 20100 22204
rect 20044 22150 20046 22202
rect 20046 22150 20098 22202
rect 20098 22150 20100 22202
rect 20044 22148 20100 22150
rect 19852 20802 19908 20804
rect 19852 20750 19854 20802
rect 19854 20750 19906 20802
rect 19906 20750 19908 20802
rect 19852 20748 19908 20750
rect 21868 26124 21924 26180
rect 21420 25676 21476 25732
rect 21420 25340 21476 25396
rect 21420 24892 21476 24948
rect 20636 22540 20692 22596
rect 21868 25340 21924 25396
rect 24668 32562 24724 32564
rect 24668 32510 24670 32562
rect 24670 32510 24722 32562
rect 24722 32510 24724 32562
rect 24668 32508 24724 32510
rect 24220 31890 24276 31892
rect 24220 31838 24222 31890
rect 24222 31838 24274 31890
rect 24274 31838 24276 31890
rect 24220 31836 24276 31838
rect 24668 31778 24724 31780
rect 24668 31726 24670 31778
rect 24670 31726 24722 31778
rect 24722 31726 24724 31778
rect 24668 31724 24724 31726
rect 24220 30380 24276 30436
rect 24556 30156 24612 30212
rect 24444 29932 24500 29988
rect 24668 29820 24724 29876
rect 24108 28588 24164 28644
rect 24332 28530 24388 28532
rect 24332 28478 24334 28530
rect 24334 28478 24386 28530
rect 24386 28478 24388 28530
rect 24332 28476 24388 28478
rect 24556 27692 24612 27748
rect 23436 27244 23492 27300
rect 24668 27468 24724 27524
rect 23324 26124 23380 26180
rect 21980 24892 22036 24948
rect 22764 25564 22820 25620
rect 21980 24722 22036 24724
rect 21980 24670 21982 24722
rect 21982 24670 22034 24722
rect 22034 24670 22036 24722
rect 21980 24668 22036 24670
rect 22316 24444 22372 24500
rect 22092 23938 22148 23940
rect 22092 23886 22094 23938
rect 22094 23886 22146 23938
rect 22146 23886 22148 23938
rect 22092 23884 22148 23886
rect 21756 22652 21812 22708
rect 22540 23602 22596 23604
rect 22540 23550 22542 23602
rect 22542 23550 22594 23602
rect 22594 23550 22596 23602
rect 22540 23548 22596 23550
rect 23324 25228 23380 25284
rect 22988 24892 23044 24948
rect 24108 26626 24164 26628
rect 24108 26574 24110 26626
rect 24110 26574 24162 26626
rect 24162 26574 24164 26626
rect 24108 26572 24164 26574
rect 24892 32562 24948 32564
rect 24892 32510 24894 32562
rect 24894 32510 24946 32562
rect 24946 32510 24948 32562
rect 24892 32508 24948 32510
rect 25340 34300 25396 34356
rect 25788 33906 25844 33908
rect 25788 33854 25790 33906
rect 25790 33854 25842 33906
rect 25842 33854 25844 33906
rect 25788 33852 25844 33854
rect 26124 34524 26180 34580
rect 25340 32786 25396 32788
rect 25340 32734 25342 32786
rect 25342 32734 25394 32786
rect 25394 32734 25396 32786
rect 25340 32732 25396 32734
rect 26236 33964 26292 34020
rect 25564 32732 25620 32788
rect 25900 32844 25956 32900
rect 25900 32674 25956 32676
rect 25900 32622 25902 32674
rect 25902 32622 25954 32674
rect 25954 32622 25956 32674
rect 25900 32620 25956 32622
rect 26012 32508 26068 32564
rect 25228 32060 25284 32116
rect 25228 31836 25284 31892
rect 26012 31724 26068 31780
rect 25116 31052 25172 31108
rect 26012 30994 26068 30996
rect 26012 30942 26014 30994
rect 26014 30942 26066 30994
rect 26066 30942 26068 30994
rect 26012 30940 26068 30942
rect 25788 30268 25844 30324
rect 25676 29820 25732 29876
rect 25228 29426 25284 29428
rect 25228 29374 25230 29426
rect 25230 29374 25282 29426
rect 25282 29374 25284 29426
rect 25228 29372 25284 29374
rect 25452 28700 25508 28756
rect 24892 28028 24948 28084
rect 24780 25340 24836 25396
rect 24556 25116 24612 25172
rect 23548 24444 23604 24500
rect 24108 24444 24164 24500
rect 23212 23884 23268 23940
rect 20748 21644 20804 21700
rect 20300 20524 20356 20580
rect 20188 20412 20244 20468
rect 19836 20186 19892 20188
rect 19836 20134 19838 20186
rect 19838 20134 19890 20186
rect 19890 20134 19892 20186
rect 19836 20132 19892 20134
rect 19940 20186 19996 20188
rect 19940 20134 19942 20186
rect 19942 20134 19994 20186
rect 19994 20134 19996 20186
rect 19940 20132 19996 20134
rect 20044 20186 20100 20188
rect 20044 20134 20046 20186
rect 20046 20134 20098 20186
rect 20098 20134 20100 20186
rect 20044 20132 20100 20134
rect 19628 19794 19684 19796
rect 19628 19742 19630 19794
rect 19630 19742 19682 19794
rect 19682 19742 19684 19794
rect 19628 19740 19684 19742
rect 19292 19682 19348 19684
rect 19292 19630 19294 19682
rect 19294 19630 19346 19682
rect 19346 19630 19348 19682
rect 19292 19628 19348 19630
rect 21196 21698 21252 21700
rect 21196 21646 21198 21698
rect 21198 21646 21250 21698
rect 21250 21646 21252 21698
rect 21196 21644 21252 21646
rect 21420 20690 21476 20692
rect 21420 20638 21422 20690
rect 21422 20638 21474 20690
rect 21474 20638 21476 20690
rect 21420 20636 21476 20638
rect 22540 20636 22596 20692
rect 20748 20412 20804 20468
rect 21644 20578 21700 20580
rect 21644 20526 21646 20578
rect 21646 20526 21698 20578
rect 21698 20526 21700 20578
rect 21644 20524 21700 20526
rect 20300 19740 20356 19796
rect 19836 18170 19892 18172
rect 19836 18118 19838 18170
rect 19838 18118 19890 18170
rect 19890 18118 19892 18170
rect 19836 18116 19892 18118
rect 19940 18170 19996 18172
rect 19940 18118 19942 18170
rect 19942 18118 19994 18170
rect 19994 18118 19996 18170
rect 19940 18116 19996 18118
rect 20044 18170 20100 18172
rect 20044 18118 20046 18170
rect 20046 18118 20098 18170
rect 20098 18118 20100 18170
rect 20044 18116 20100 18118
rect 18732 16828 18788 16884
rect 19516 16828 19572 16884
rect 17500 14588 17556 14644
rect 16828 13746 16884 13748
rect 16828 13694 16830 13746
rect 16830 13694 16882 13746
rect 16882 13694 16884 13746
rect 16828 13692 16884 13694
rect 17836 14700 17892 14756
rect 4476 13130 4532 13132
rect 4476 13078 4478 13130
rect 4478 13078 4530 13130
rect 4530 13078 4532 13130
rect 4476 13076 4532 13078
rect 4580 13130 4636 13132
rect 4580 13078 4582 13130
rect 4582 13078 4634 13130
rect 4634 13078 4636 13130
rect 4580 13076 4636 13078
rect 4684 13130 4740 13132
rect 4684 13078 4686 13130
rect 4686 13078 4738 13130
rect 4738 13078 4740 13130
rect 4684 13076 4740 13078
rect 19180 14754 19236 14756
rect 19180 14702 19182 14754
rect 19182 14702 19234 14754
rect 19234 14702 19236 14754
rect 19180 14700 19236 14702
rect 18396 14364 18452 14420
rect 18284 13692 18340 13748
rect 22540 19964 22596 20020
rect 22092 19516 22148 19572
rect 21868 16716 21924 16772
rect 22092 16604 22148 16660
rect 19836 16154 19892 16156
rect 19836 16102 19838 16154
rect 19838 16102 19890 16154
rect 19890 16102 19892 16154
rect 19836 16100 19892 16102
rect 19940 16154 19996 16156
rect 19940 16102 19942 16154
rect 19942 16102 19994 16154
rect 19994 16102 19996 16154
rect 19940 16100 19996 16102
rect 20044 16154 20100 16156
rect 20044 16102 20046 16154
rect 20046 16102 20098 16154
rect 20098 16102 20100 16154
rect 20044 16100 20100 16102
rect 19740 15762 19796 15764
rect 19740 15710 19742 15762
rect 19742 15710 19794 15762
rect 19794 15710 19796 15762
rect 19740 15708 19796 15710
rect 19852 15596 19908 15652
rect 19628 14642 19684 14644
rect 19628 14590 19630 14642
rect 19630 14590 19682 14642
rect 19682 14590 19684 14642
rect 19628 14588 19684 14590
rect 23436 23602 23492 23604
rect 23436 23550 23438 23602
rect 23438 23550 23490 23602
rect 23490 23550 23492 23602
rect 23436 23548 23492 23550
rect 22764 21644 22820 21700
rect 23212 20636 23268 20692
rect 23660 20690 23716 20692
rect 23660 20638 23662 20690
rect 23662 20638 23714 20690
rect 23714 20638 23716 20690
rect 23660 20636 23716 20638
rect 22764 19570 22820 19572
rect 22764 19518 22766 19570
rect 22766 19518 22818 19570
rect 22818 19518 22820 19570
rect 22764 19516 22820 19518
rect 22988 16770 23044 16772
rect 22988 16718 22990 16770
rect 22990 16718 23042 16770
rect 23042 16718 23044 16770
rect 22988 16716 23044 16718
rect 23212 16716 23268 16772
rect 22540 16492 22596 16548
rect 23660 16716 23716 16772
rect 23436 16546 23492 16548
rect 23436 16494 23438 16546
rect 23438 16494 23490 16546
rect 23490 16494 23492 16546
rect 23436 16492 23492 16494
rect 22092 15596 22148 15652
rect 20188 14866 20244 14868
rect 20188 14814 20190 14866
rect 20190 14814 20242 14866
rect 20242 14814 20244 14866
rect 20188 14812 20244 14814
rect 20748 15036 20804 15092
rect 19964 14364 20020 14420
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18620 11564 18676 11620
rect 4476 11114 4532 11116
rect 4476 11062 4478 11114
rect 4478 11062 4530 11114
rect 4530 11062 4532 11114
rect 4476 11060 4532 11062
rect 4580 11114 4636 11116
rect 4580 11062 4582 11114
rect 4582 11062 4634 11114
rect 4634 11062 4636 11114
rect 4580 11060 4636 11062
rect 4684 11114 4740 11116
rect 4684 11062 4686 11114
rect 4686 11062 4738 11114
rect 4738 11062 4740 11114
rect 4684 11060 4740 11062
rect 18172 9826 18228 9828
rect 18172 9774 18174 9826
rect 18174 9774 18226 9826
rect 18226 9774 18228 9826
rect 18172 9772 18228 9774
rect 19836 12122 19892 12124
rect 19836 12070 19838 12122
rect 19838 12070 19890 12122
rect 19890 12070 19892 12122
rect 19836 12068 19892 12070
rect 19940 12122 19996 12124
rect 19940 12070 19942 12122
rect 19942 12070 19994 12122
rect 19994 12070 19996 12122
rect 19940 12068 19996 12070
rect 20044 12122 20100 12124
rect 20044 12070 20046 12122
rect 20046 12070 20098 12122
rect 20098 12070 20100 12122
rect 20044 12068 20100 12070
rect 19740 11618 19796 11620
rect 19740 11566 19742 11618
rect 19742 11566 19794 11618
rect 19794 11566 19796 11618
rect 19740 11564 19796 11566
rect 18956 10668 19012 10724
rect 19404 11506 19460 11508
rect 19404 11454 19406 11506
rect 19406 11454 19458 11506
rect 19458 11454 19460 11506
rect 19404 11452 19460 11454
rect 20524 11452 20580 11508
rect 19836 10106 19892 10108
rect 19836 10054 19838 10106
rect 19838 10054 19890 10106
rect 19890 10054 19892 10106
rect 19836 10052 19892 10054
rect 19940 10106 19996 10108
rect 19940 10054 19942 10106
rect 19942 10054 19994 10106
rect 19994 10054 19996 10106
rect 19940 10052 19996 10054
rect 20044 10106 20100 10108
rect 20044 10054 20046 10106
rect 20046 10054 20098 10106
rect 20098 10054 20100 10106
rect 20044 10052 20100 10054
rect 21420 15036 21476 15092
rect 21420 14530 21476 14532
rect 21420 14478 21422 14530
rect 21422 14478 21474 14530
rect 21474 14478 21476 14530
rect 21420 14476 21476 14478
rect 21756 14364 21812 14420
rect 22540 14418 22596 14420
rect 22540 14366 22542 14418
rect 22542 14366 22594 14418
rect 22594 14366 22596 14418
rect 22540 14364 22596 14366
rect 20972 13634 21028 13636
rect 20972 13582 20974 13634
rect 20974 13582 21026 13634
rect 21026 13582 21028 13634
rect 20972 13580 21028 13582
rect 21756 13580 21812 13636
rect 23660 15874 23716 15876
rect 23660 15822 23662 15874
rect 23662 15822 23714 15874
rect 23714 15822 23716 15874
rect 23660 15820 23716 15822
rect 25340 28418 25396 28420
rect 25340 28366 25342 28418
rect 25342 28366 25394 28418
rect 25394 28366 25396 28418
rect 25340 28364 25396 28366
rect 25340 28082 25396 28084
rect 25340 28030 25342 28082
rect 25342 28030 25394 28082
rect 25394 28030 25396 28082
rect 25340 28028 25396 28030
rect 29148 44940 29204 44996
rect 28252 44658 28308 44660
rect 28252 44606 28254 44658
rect 28254 44606 28306 44658
rect 28306 44606 28308 44658
rect 28252 44604 28308 44606
rect 28700 44604 28756 44660
rect 29036 43986 29092 43988
rect 29036 43934 29038 43986
rect 29038 43934 29090 43986
rect 29090 43934 29092 43986
rect 29036 43932 29092 43934
rect 32620 46956 32676 47012
rect 33068 46844 33124 46900
rect 32508 46732 32564 46788
rect 33180 46674 33236 46676
rect 33180 46622 33182 46674
rect 33182 46622 33234 46674
rect 33234 46622 33236 46674
rect 33180 46620 33236 46622
rect 32508 46060 32564 46116
rect 36988 48860 37044 48916
rect 35196 47402 35252 47404
rect 35196 47350 35198 47402
rect 35198 47350 35250 47402
rect 35250 47350 35252 47402
rect 35196 47348 35252 47350
rect 35300 47402 35356 47404
rect 35300 47350 35302 47402
rect 35302 47350 35354 47402
rect 35354 47350 35356 47402
rect 35300 47348 35356 47350
rect 35404 47402 35460 47404
rect 35404 47350 35406 47402
rect 35406 47350 35458 47402
rect 35458 47350 35460 47402
rect 35404 47348 35460 47350
rect 34188 46956 34244 47012
rect 34076 46898 34132 46900
rect 34076 46846 34078 46898
rect 34078 46846 34130 46898
rect 34130 46846 34132 46898
rect 34076 46844 34132 46846
rect 33068 46002 33124 46004
rect 33068 45950 33070 46002
rect 33070 45950 33122 46002
rect 33122 45950 33124 46002
rect 33068 45948 33124 45950
rect 32396 44940 32452 44996
rect 32620 45052 32676 45108
rect 28140 43596 28196 43652
rect 28140 42754 28196 42756
rect 28140 42702 28142 42754
rect 28142 42702 28194 42754
rect 28194 42702 28196 42754
rect 28140 42700 28196 42702
rect 30268 43932 30324 43988
rect 29036 42924 29092 42980
rect 31724 43932 31780 43988
rect 32172 43986 32228 43988
rect 32172 43934 32174 43986
rect 32174 43934 32226 43986
rect 32226 43934 32228 43986
rect 32172 43932 32228 43934
rect 32060 43708 32116 43764
rect 29596 42754 29652 42756
rect 29596 42702 29598 42754
rect 29598 42702 29650 42754
rect 29650 42702 29652 42754
rect 29596 42700 29652 42702
rect 29372 42140 29428 42196
rect 29708 42028 29764 42084
rect 30268 41970 30324 41972
rect 30268 41918 30270 41970
rect 30270 41918 30322 41970
rect 30322 41918 30324 41970
rect 30268 41916 30324 41918
rect 28476 41804 28532 41860
rect 28140 41746 28196 41748
rect 28140 41694 28142 41746
rect 28142 41694 28194 41746
rect 28194 41694 28196 41746
rect 28140 41692 28196 41694
rect 28812 41746 28868 41748
rect 28812 41694 28814 41746
rect 28814 41694 28866 41746
rect 28866 41694 28868 41746
rect 28812 41692 28868 41694
rect 28028 41020 28084 41076
rect 27916 40348 27972 40404
rect 27356 38722 27412 38724
rect 27356 38670 27358 38722
rect 27358 38670 27410 38722
rect 27410 38670 27412 38722
rect 27356 38668 27412 38670
rect 27356 36594 27412 36596
rect 27356 36542 27358 36594
rect 27358 36542 27410 36594
rect 27410 36542 27412 36594
rect 27356 36540 27412 36542
rect 27916 36482 27972 36484
rect 27916 36430 27918 36482
rect 27918 36430 27970 36482
rect 27970 36430 27972 36482
rect 27916 36428 27972 36430
rect 27020 35810 27076 35812
rect 27020 35758 27022 35810
rect 27022 35758 27074 35810
rect 27074 35758 27076 35810
rect 27020 35756 27076 35758
rect 26908 35196 26964 35252
rect 28364 36540 28420 36596
rect 29260 36594 29316 36596
rect 29260 36542 29262 36594
rect 29262 36542 29314 36594
rect 29314 36542 29316 36594
rect 29260 36540 29316 36542
rect 27580 35196 27636 35252
rect 26684 34802 26740 34804
rect 26684 34750 26686 34802
rect 26686 34750 26738 34802
rect 26738 34750 26740 34802
rect 26684 34748 26740 34750
rect 26684 33964 26740 34020
rect 27356 33906 27412 33908
rect 27356 33854 27358 33906
rect 27358 33854 27410 33906
rect 27410 33854 27412 33906
rect 27356 33852 27412 33854
rect 29484 35532 29540 35588
rect 28028 34802 28084 34804
rect 28028 34750 28030 34802
rect 28030 34750 28082 34802
rect 28082 34750 28084 34802
rect 28028 34748 28084 34750
rect 28364 34524 28420 34580
rect 29260 34748 29316 34804
rect 27916 33852 27972 33908
rect 26460 32060 26516 32116
rect 26348 31836 26404 31892
rect 25900 29932 25956 29988
rect 26460 30156 26516 30212
rect 26124 29762 26180 29764
rect 26124 29710 26126 29762
rect 26126 29710 26178 29762
rect 26178 29710 26180 29762
rect 26124 29708 26180 29710
rect 26348 29762 26404 29764
rect 26348 29710 26350 29762
rect 26350 29710 26402 29762
rect 26402 29710 26404 29762
rect 26348 29708 26404 29710
rect 26348 29090 26404 29092
rect 26348 29038 26350 29090
rect 26350 29038 26402 29090
rect 26402 29038 26404 29090
rect 26348 29036 26404 29038
rect 27020 30828 27076 30884
rect 28588 32956 28644 33012
rect 27916 31052 27972 31108
rect 26684 30380 26740 30436
rect 27020 30044 27076 30100
rect 25564 27916 25620 27972
rect 26012 28252 26068 28308
rect 25676 27746 25732 27748
rect 25676 27694 25678 27746
rect 25678 27694 25730 27746
rect 25730 27694 25732 27746
rect 25676 27692 25732 27694
rect 25900 27858 25956 27860
rect 25900 27806 25902 27858
rect 25902 27806 25954 27858
rect 25954 27806 25956 27858
rect 25900 27804 25956 27806
rect 25788 27132 25844 27188
rect 25676 26796 25732 26852
rect 25564 26124 25620 26180
rect 25452 25228 25508 25284
rect 25564 25340 25620 25396
rect 24892 24610 24948 24612
rect 24892 24558 24894 24610
rect 24894 24558 24946 24610
rect 24946 24558 24948 24610
rect 24892 24556 24948 24558
rect 25004 24444 25060 24500
rect 24556 23938 24612 23940
rect 24556 23886 24558 23938
rect 24558 23886 24610 23938
rect 24610 23886 24612 23938
rect 24556 23884 24612 23886
rect 24780 23772 24836 23828
rect 24108 23602 24164 23604
rect 24108 23550 24110 23602
rect 24110 23550 24162 23602
rect 24162 23550 24164 23602
rect 24108 23548 24164 23550
rect 23884 23436 23940 23492
rect 23884 22652 23940 22708
rect 25116 23714 25172 23716
rect 25116 23662 25118 23714
rect 25118 23662 25170 23714
rect 25170 23662 25172 23714
rect 25116 23660 25172 23662
rect 24892 23436 24948 23492
rect 25564 24780 25620 24836
rect 25452 24444 25508 24500
rect 25228 22594 25284 22596
rect 25228 22542 25230 22594
rect 25230 22542 25282 22594
rect 25282 22542 25284 22594
rect 25228 22540 25284 22542
rect 24556 21644 24612 21700
rect 24220 21586 24276 21588
rect 24220 21534 24222 21586
rect 24222 21534 24274 21586
rect 24274 21534 24276 21586
rect 24220 21532 24276 21534
rect 24780 20636 24836 20692
rect 24220 20524 24276 20580
rect 24332 19628 24388 19684
rect 24220 16716 24276 16772
rect 23996 16492 24052 16548
rect 24108 16604 24164 16660
rect 24108 15484 24164 15540
rect 23324 14476 23380 14532
rect 23548 14364 23604 14420
rect 23660 13356 23716 13412
rect 26236 27804 26292 27860
rect 26236 27356 26292 27412
rect 26124 27132 26180 27188
rect 26124 26908 26180 26964
rect 26460 27020 26516 27076
rect 26348 26514 26404 26516
rect 26348 26462 26350 26514
rect 26350 26462 26402 26514
rect 26402 26462 26404 26514
rect 26348 26460 26404 26462
rect 26236 25452 26292 25508
rect 26124 24444 26180 24500
rect 25900 23884 25956 23940
rect 25452 23660 25508 23716
rect 27132 29874 27188 29876
rect 27132 29822 27134 29874
rect 27134 29822 27186 29874
rect 27186 29822 27188 29874
rect 27132 29820 27188 29822
rect 27132 29148 27188 29204
rect 27468 30380 27524 30436
rect 27132 28476 27188 28532
rect 27244 28588 27300 28644
rect 27132 28140 27188 28196
rect 26908 27970 26964 27972
rect 26908 27918 26910 27970
rect 26910 27918 26962 27970
rect 26962 27918 26964 27970
rect 26908 27916 26964 27918
rect 27020 27804 27076 27860
rect 26796 27356 26852 27412
rect 26796 26908 26852 26964
rect 26796 26460 26852 26516
rect 27020 27580 27076 27636
rect 27580 28418 27636 28420
rect 27580 28366 27582 28418
rect 27582 28366 27634 28418
rect 27634 28366 27636 28418
rect 27580 28364 27636 28366
rect 28140 30940 28196 30996
rect 28140 30380 28196 30436
rect 28476 31106 28532 31108
rect 28476 31054 28478 31106
rect 28478 31054 28530 31106
rect 28530 31054 28532 31106
rect 28476 31052 28532 31054
rect 29148 30380 29204 30436
rect 28364 29708 28420 29764
rect 28028 28812 28084 28868
rect 28140 28700 28196 28756
rect 28812 29708 28868 29764
rect 28476 29372 28532 29428
rect 28812 29372 28868 29428
rect 28252 28642 28308 28644
rect 28252 28590 28254 28642
rect 28254 28590 28306 28642
rect 28306 28590 28308 28642
rect 28252 28588 28308 28590
rect 27916 28252 27972 28308
rect 28476 27970 28532 27972
rect 28476 27918 28478 27970
rect 28478 27918 28530 27970
rect 28530 27918 28532 27970
rect 28476 27916 28532 27918
rect 28140 27858 28196 27860
rect 28140 27806 28142 27858
rect 28142 27806 28194 27858
rect 28194 27806 28196 27858
rect 28140 27804 28196 27806
rect 28140 27468 28196 27524
rect 27356 26796 27412 26852
rect 29148 28700 29204 28756
rect 30380 40236 30436 40292
rect 30940 41746 30996 41748
rect 30940 41694 30942 41746
rect 30942 41694 30994 41746
rect 30994 41694 30996 41746
rect 30940 41692 30996 41694
rect 30716 39676 30772 39732
rect 29932 38668 29988 38724
rect 29820 35810 29876 35812
rect 29820 35758 29822 35810
rect 29822 35758 29874 35810
rect 29874 35758 29876 35810
rect 29820 35756 29876 35758
rect 29708 35196 29764 35252
rect 29372 34578 29428 34580
rect 29372 34526 29374 34578
rect 29374 34526 29426 34578
rect 29426 34526 29428 34578
rect 29372 34524 29428 34526
rect 29484 32956 29540 33012
rect 29820 32844 29876 32900
rect 30268 37660 30324 37716
rect 30604 35644 30660 35700
rect 31836 40236 31892 40292
rect 31164 39730 31220 39732
rect 31164 39678 31166 39730
rect 31166 39678 31218 39730
rect 31218 39678 31220 39730
rect 31164 39676 31220 39678
rect 31052 37714 31108 37716
rect 31052 37662 31054 37714
rect 31054 37662 31106 37714
rect 31106 37662 31108 37714
rect 31052 37660 31108 37662
rect 31388 35644 31444 35700
rect 33740 45890 33796 45892
rect 33740 45838 33742 45890
rect 33742 45838 33794 45890
rect 33794 45838 33796 45890
rect 33740 45836 33796 45838
rect 33404 43932 33460 43988
rect 33628 44044 33684 44100
rect 33292 43036 33348 43092
rect 32956 42866 33012 42868
rect 32956 42814 32958 42866
rect 32958 42814 33010 42866
rect 33010 42814 33012 42866
rect 32956 42812 33012 42814
rect 33404 42140 33460 42196
rect 34076 44994 34132 44996
rect 34076 44942 34078 44994
rect 34078 44942 34130 44994
rect 34130 44942 34132 44994
rect 34076 44940 34132 44942
rect 34860 46956 34916 47012
rect 35196 46620 35252 46676
rect 34524 46172 34580 46228
rect 35196 45386 35252 45388
rect 35196 45334 35198 45386
rect 35198 45334 35250 45386
rect 35250 45334 35252 45386
rect 35196 45332 35252 45334
rect 35300 45386 35356 45388
rect 35300 45334 35302 45386
rect 35302 45334 35354 45386
rect 35354 45334 35356 45386
rect 35300 45332 35356 45334
rect 35404 45386 35460 45388
rect 35404 45334 35406 45386
rect 35406 45334 35458 45386
rect 35458 45334 35460 45386
rect 35404 45332 35460 45334
rect 39228 48914 39284 48916
rect 39228 48862 39230 48914
rect 39230 48862 39282 48914
rect 39282 48862 39284 48914
rect 39228 48860 39284 48862
rect 38780 48802 38836 48804
rect 38780 48750 38782 48802
rect 38782 48750 38834 48802
rect 38834 48750 38836 48802
rect 38780 48748 38836 48750
rect 40684 48802 40740 48804
rect 40684 48750 40686 48802
rect 40686 48750 40738 48802
rect 40738 48750 40740 48802
rect 40684 48748 40740 48750
rect 38332 48690 38388 48692
rect 38332 48638 38334 48690
rect 38334 48638 38386 48690
rect 38386 48638 38388 48690
rect 38332 48636 38388 48638
rect 39004 48636 39060 48692
rect 36988 46844 37044 46900
rect 37548 46898 37604 46900
rect 37548 46846 37550 46898
rect 37550 46846 37602 46898
rect 37602 46846 37604 46898
rect 37548 46844 37604 46846
rect 36988 45276 37044 45332
rect 35308 45106 35364 45108
rect 35308 45054 35310 45106
rect 35310 45054 35362 45106
rect 35362 45054 35364 45106
rect 35308 45052 35364 45054
rect 34188 44828 34244 44884
rect 34524 44940 34580 44996
rect 34188 44098 34244 44100
rect 34188 44046 34190 44098
rect 34190 44046 34242 44098
rect 34242 44046 34244 44098
rect 34188 44044 34244 44046
rect 33964 43090 34020 43092
rect 33964 43038 33966 43090
rect 33966 43038 34018 43090
rect 34018 43038 34020 43090
rect 33964 43036 34020 43038
rect 34636 42812 34692 42868
rect 33852 41916 33908 41972
rect 34412 41970 34468 41972
rect 34412 41918 34414 41970
rect 34414 41918 34466 41970
rect 34466 41918 34468 41970
rect 34412 41916 34468 41918
rect 33964 41858 34020 41860
rect 33964 41806 33966 41858
rect 33966 41806 34018 41858
rect 34018 41806 34020 41858
rect 33964 41804 34020 41806
rect 34748 41468 34804 41524
rect 33516 39900 33572 39956
rect 32172 37996 32228 38052
rect 31836 35810 31892 35812
rect 31836 35758 31838 35810
rect 31838 35758 31890 35810
rect 31890 35758 31892 35810
rect 31836 35756 31892 35758
rect 30716 33794 30772 33796
rect 30716 33742 30718 33794
rect 30718 33742 30770 33794
rect 30770 33742 30772 33794
rect 30716 33740 30772 33742
rect 30268 32732 30324 32788
rect 29372 31890 29428 31892
rect 29372 31838 29374 31890
rect 29374 31838 29426 31890
rect 29426 31838 29428 31890
rect 29372 31836 29428 31838
rect 29484 30604 29540 30660
rect 30492 32674 30548 32676
rect 30492 32622 30494 32674
rect 30494 32622 30546 32674
rect 30546 32622 30548 32674
rect 30492 32620 30548 32622
rect 30156 30764 30212 30772
rect 30156 30716 30158 30764
rect 30158 30716 30210 30764
rect 30210 30716 30212 30764
rect 29932 30658 29988 30660
rect 29932 30606 29934 30658
rect 29934 30606 29986 30658
rect 29986 30606 29988 30658
rect 29932 30604 29988 30606
rect 30044 30434 30100 30436
rect 30044 30382 30046 30434
rect 30046 30382 30098 30434
rect 30098 30382 30100 30434
rect 30044 30380 30100 30382
rect 29484 29036 29540 29092
rect 29932 28924 29988 28980
rect 28812 27858 28868 27860
rect 28812 27806 28814 27858
rect 28814 27806 28866 27858
rect 28866 27806 28868 27858
rect 28812 27804 28868 27806
rect 29260 28476 29316 28532
rect 29260 27468 29316 27524
rect 28700 27020 28756 27076
rect 27356 26626 27412 26628
rect 27356 26574 27358 26626
rect 27358 26574 27410 26626
rect 27410 26574 27412 26626
rect 27356 26572 27412 26574
rect 27468 26514 27524 26516
rect 27468 26462 27470 26514
rect 27470 26462 27522 26514
rect 27522 26462 27524 26514
rect 27468 26460 27524 26462
rect 26348 24108 26404 24164
rect 27020 26124 27076 26180
rect 26572 24498 26628 24500
rect 26572 24446 26574 24498
rect 26574 24446 26626 24498
rect 26626 24446 26628 24498
rect 26572 24444 26628 24446
rect 27804 25676 27860 25732
rect 27468 25564 27524 25620
rect 26908 25506 26964 25508
rect 26908 25454 26910 25506
rect 26910 25454 26962 25506
rect 26962 25454 26964 25506
rect 26908 25452 26964 25454
rect 27020 24834 27076 24836
rect 27020 24782 27022 24834
rect 27022 24782 27074 24834
rect 27074 24782 27076 24834
rect 27020 24780 27076 24782
rect 26684 23938 26740 23940
rect 26684 23886 26686 23938
rect 26686 23886 26738 23938
rect 26738 23886 26740 23938
rect 26684 23884 26740 23886
rect 27244 24556 27300 24612
rect 26348 23826 26404 23828
rect 26348 23774 26350 23826
rect 26350 23774 26402 23826
rect 26402 23774 26404 23826
rect 26348 23772 26404 23774
rect 25788 23548 25844 23604
rect 25676 22540 25732 22596
rect 26124 22316 26180 22372
rect 26348 23548 26404 23604
rect 25564 21698 25620 21700
rect 25564 21646 25566 21698
rect 25566 21646 25618 21698
rect 25618 21646 25620 21698
rect 25564 21644 25620 21646
rect 26124 21532 26180 21588
rect 26236 21420 26292 21476
rect 24892 19292 24948 19348
rect 25340 20076 25396 20132
rect 25564 20188 25620 20244
rect 26796 21420 26852 21476
rect 25900 20076 25956 20132
rect 28476 26738 28532 26740
rect 28476 26686 28478 26738
rect 28478 26686 28530 26738
rect 28530 26686 28532 26738
rect 28476 26684 28532 26686
rect 28252 26460 28308 26516
rect 28476 25676 28532 25732
rect 27580 23772 27636 23828
rect 27804 23602 27860 23604
rect 27804 23550 27806 23602
rect 27806 23550 27858 23602
rect 27858 23550 27860 23602
rect 27804 23548 27860 23550
rect 27468 20300 27524 20356
rect 26236 19964 26292 20020
rect 26460 20076 26516 20132
rect 26236 19682 26292 19684
rect 26236 19630 26238 19682
rect 26238 19630 26290 19682
rect 26290 19630 26292 19682
rect 26236 19628 26292 19630
rect 25564 19516 25620 19572
rect 24444 16658 24500 16660
rect 24444 16606 24446 16658
rect 24446 16606 24498 16658
rect 24498 16606 24500 16658
rect 24444 16604 24500 16606
rect 24780 16658 24836 16660
rect 24780 16606 24782 16658
rect 24782 16606 24834 16658
rect 24834 16606 24836 16658
rect 24780 16604 24836 16606
rect 26012 18562 26068 18564
rect 26012 18510 26014 18562
rect 26014 18510 26066 18562
rect 26066 18510 26068 18562
rect 26012 18508 26068 18510
rect 26796 17836 26852 17892
rect 28588 25340 28644 25396
rect 28812 26460 28868 26516
rect 28924 26348 28980 26404
rect 28140 25116 28196 25172
rect 28140 24556 28196 24612
rect 28252 24668 28308 24724
rect 28252 23660 28308 23716
rect 28364 24444 28420 24500
rect 28700 23826 28756 23828
rect 28700 23774 28702 23826
rect 28702 23774 28754 23826
rect 28754 23774 28756 23826
rect 28700 23772 28756 23774
rect 29708 27580 29764 27636
rect 29596 26348 29652 26404
rect 30492 31052 30548 31108
rect 30492 30716 30548 30772
rect 30940 30716 30996 30772
rect 30604 30658 30660 30660
rect 30604 30606 30606 30658
rect 30606 30606 30658 30658
rect 30658 30606 30660 30658
rect 30604 30604 30660 30606
rect 30716 29932 30772 29988
rect 30716 29036 30772 29092
rect 30156 27356 30212 27412
rect 31276 33740 31332 33796
rect 31164 32844 31220 32900
rect 31276 32620 31332 32676
rect 31836 33906 31892 33908
rect 31836 33854 31838 33906
rect 31838 33854 31890 33906
rect 31890 33854 31892 33906
rect 31836 33852 31892 33854
rect 32396 33628 32452 33684
rect 33516 38556 33572 38612
rect 33180 38050 33236 38052
rect 33180 37998 33182 38050
rect 33182 37998 33234 38050
rect 33234 37998 33236 38050
rect 33180 37996 33236 37998
rect 34076 39730 34132 39732
rect 34076 39678 34078 39730
rect 34078 39678 34130 39730
rect 34130 39678 34132 39730
rect 34076 39676 34132 39678
rect 34412 38556 34468 38612
rect 33180 35698 33236 35700
rect 33180 35646 33182 35698
rect 33182 35646 33234 35698
rect 33234 35646 33236 35698
rect 33180 35644 33236 35646
rect 32732 35308 32788 35364
rect 31164 30882 31220 30884
rect 31164 30830 31166 30882
rect 31166 30830 31218 30882
rect 31218 30830 31220 30882
rect 31164 30828 31220 30830
rect 31276 30658 31332 30660
rect 31276 30606 31278 30658
rect 31278 30606 31330 30658
rect 31330 30606 31332 30658
rect 31276 30604 31332 30606
rect 31164 29036 31220 29092
rect 30044 26684 30100 26740
rect 29372 25340 29428 25396
rect 30044 26514 30100 26516
rect 30044 26462 30046 26514
rect 30046 26462 30098 26514
rect 30098 26462 30100 26514
rect 30044 26460 30100 26462
rect 30492 26236 30548 26292
rect 30940 26348 30996 26404
rect 30716 25900 30772 25956
rect 30380 25564 30436 25620
rect 32060 30882 32116 30884
rect 32060 30830 32062 30882
rect 32062 30830 32114 30882
rect 32114 30830 32116 30882
rect 32060 30828 32116 30830
rect 31836 30380 31892 30436
rect 31612 29484 31668 29540
rect 31500 27858 31556 27860
rect 31500 27806 31502 27858
rect 31502 27806 31554 27858
rect 31554 27806 31556 27858
rect 31500 27804 31556 27806
rect 32060 28530 32116 28532
rect 32060 28478 32062 28530
rect 32062 28478 32114 28530
rect 32114 28478 32116 28530
rect 32060 28476 32116 28478
rect 32508 30716 32564 30772
rect 32620 31164 32676 31220
rect 32732 30828 32788 30884
rect 32396 30268 32452 30324
rect 32396 27804 32452 27860
rect 31836 27634 31892 27636
rect 31836 27582 31838 27634
rect 31838 27582 31890 27634
rect 31890 27582 31892 27634
rect 31836 27580 31892 27582
rect 31612 26908 31668 26964
rect 31276 26236 31332 26292
rect 31388 26572 31444 26628
rect 31164 25730 31220 25732
rect 31164 25678 31166 25730
rect 31166 25678 31218 25730
rect 31218 25678 31220 25730
rect 31164 25676 31220 25678
rect 31052 25116 31108 25172
rect 30268 24892 30324 24948
rect 30044 24780 30100 24836
rect 29820 24722 29876 24724
rect 29820 24670 29822 24722
rect 29822 24670 29874 24722
rect 29874 24670 29876 24722
rect 29820 24668 29876 24670
rect 29260 24498 29316 24500
rect 29260 24446 29262 24498
rect 29262 24446 29314 24498
rect 29314 24446 29316 24498
rect 29260 24444 29316 24446
rect 29036 23714 29092 23716
rect 29036 23662 29038 23714
rect 29038 23662 29090 23714
rect 29090 23662 29092 23714
rect 29036 23660 29092 23662
rect 28924 23548 28980 23604
rect 28924 21420 28980 21476
rect 28476 20300 28532 20356
rect 27468 20076 27524 20132
rect 25228 15484 25284 15540
rect 25004 14812 25060 14868
rect 24444 13858 24500 13860
rect 24444 13806 24446 13858
rect 24446 13806 24498 13858
rect 24498 13806 24500 13858
rect 24444 13804 24500 13806
rect 25340 14700 25396 14756
rect 26012 16716 26068 16772
rect 25676 13804 25732 13860
rect 26796 16604 26852 16660
rect 26684 14700 26740 14756
rect 25900 14476 25956 14532
rect 25340 13692 25396 13748
rect 24892 13468 24948 13524
rect 21756 11452 21812 11508
rect 21420 10722 21476 10724
rect 21420 10670 21422 10722
rect 21422 10670 21474 10722
rect 21474 10670 21476 10722
rect 21420 10668 21476 10670
rect 20748 10498 20804 10500
rect 20748 10446 20750 10498
rect 20750 10446 20802 10498
rect 20802 10446 20804 10498
rect 20748 10444 20804 10446
rect 20300 9996 20356 10052
rect 19068 9772 19124 9828
rect 22988 11506 23044 11508
rect 22988 11454 22990 11506
rect 22990 11454 23042 11506
rect 23042 11454 23044 11506
rect 22988 11452 23044 11454
rect 22876 10892 22932 10948
rect 22316 10498 22372 10500
rect 22316 10446 22318 10498
rect 22318 10446 22370 10498
rect 22370 10446 22372 10498
rect 22316 10444 22372 10446
rect 21644 9996 21700 10052
rect 4476 9098 4532 9100
rect 4476 9046 4478 9098
rect 4478 9046 4530 9098
rect 4530 9046 4532 9098
rect 4476 9044 4532 9046
rect 4580 9098 4636 9100
rect 4580 9046 4582 9098
rect 4582 9046 4634 9098
rect 4634 9046 4636 9098
rect 4580 9044 4636 9046
rect 4684 9098 4740 9100
rect 4684 9046 4686 9098
rect 4686 9046 4738 9098
rect 4738 9046 4740 9098
rect 4684 9044 4740 9046
rect 19836 8090 19892 8092
rect 19836 8038 19838 8090
rect 19838 8038 19890 8090
rect 19890 8038 19892 8090
rect 19836 8036 19892 8038
rect 19940 8090 19996 8092
rect 19940 8038 19942 8090
rect 19942 8038 19994 8090
rect 19994 8038 19996 8090
rect 19940 8036 19996 8038
rect 20044 8090 20100 8092
rect 20044 8038 20046 8090
rect 20046 8038 20098 8090
rect 20098 8038 20100 8090
rect 20044 8036 20100 8038
rect 22092 8706 22148 8708
rect 22092 8654 22094 8706
rect 22094 8654 22146 8706
rect 22146 8654 22148 8706
rect 22092 8652 22148 8654
rect 23996 10892 24052 10948
rect 24444 11564 24500 11620
rect 23436 9772 23492 9828
rect 23772 9772 23828 9828
rect 22540 8706 22596 8708
rect 22540 8654 22542 8706
rect 22542 8654 22594 8706
rect 22594 8654 22596 8706
rect 22540 8652 22596 8654
rect 25228 11676 25284 11732
rect 23772 8652 23828 8708
rect 22988 8540 23044 8596
rect 23660 8594 23716 8596
rect 23660 8542 23662 8594
rect 23662 8542 23714 8594
rect 23714 8542 23716 8594
rect 23660 8540 23716 8542
rect 23996 9660 24052 9716
rect 22876 8428 22932 8484
rect 24668 9714 24724 9716
rect 24668 9662 24670 9714
rect 24670 9662 24722 9714
rect 24722 9662 24724 9714
rect 24668 9660 24724 9662
rect 23996 8482 24052 8484
rect 23996 8430 23998 8482
rect 23998 8430 24050 8482
rect 24050 8430 24052 8482
rect 23996 8428 24052 8430
rect 27132 18732 27188 18788
rect 27804 17890 27860 17892
rect 27804 17838 27806 17890
rect 27806 17838 27858 17890
rect 27858 17838 27860 17890
rect 27804 17836 27860 17838
rect 27020 15932 27076 15988
rect 27132 14754 27188 14756
rect 27132 14702 27134 14754
rect 27134 14702 27186 14754
rect 27186 14702 27188 14754
rect 27132 14700 27188 14702
rect 26684 14530 26740 14532
rect 26684 14478 26686 14530
rect 26686 14478 26738 14530
rect 26738 14478 26740 14530
rect 26684 14476 26740 14478
rect 26236 13522 26292 13524
rect 26236 13470 26238 13522
rect 26238 13470 26290 13522
rect 26290 13470 26292 13522
rect 26236 13468 26292 13470
rect 27020 13468 27076 13524
rect 27804 16546 27860 16548
rect 27804 16494 27806 16546
rect 27806 16494 27858 16546
rect 27858 16494 27860 16546
rect 27804 16492 27860 16494
rect 30940 23826 30996 23828
rect 30940 23774 30942 23826
rect 30942 23774 30994 23826
rect 30994 23774 30996 23826
rect 30940 23772 30996 23774
rect 32396 27020 32452 27076
rect 31612 26460 31668 26516
rect 31612 26236 31668 26292
rect 31388 25004 31444 25060
rect 32172 25730 32228 25732
rect 32172 25678 32174 25730
rect 32174 25678 32226 25730
rect 32226 25678 32228 25730
rect 32172 25676 32228 25678
rect 32508 28476 32564 28532
rect 33516 35644 33572 35700
rect 34076 35698 34132 35700
rect 34076 35646 34078 35698
rect 34078 35646 34130 35698
rect 34130 35646 34132 35698
rect 34076 35644 34132 35646
rect 33740 34802 33796 34804
rect 33740 34750 33742 34802
rect 33742 34750 33794 34802
rect 33794 34750 33796 34802
rect 33740 34748 33796 34750
rect 36092 44882 36148 44884
rect 36092 44830 36094 44882
rect 36094 44830 36146 44882
rect 36146 44830 36148 44882
rect 36092 44828 36148 44830
rect 37548 44994 37604 44996
rect 37548 44942 37550 44994
rect 37550 44942 37602 44994
rect 37602 44942 37604 44994
rect 37548 44940 37604 44942
rect 37884 45276 37940 45332
rect 36876 44828 36932 44884
rect 35196 43370 35252 43372
rect 35196 43318 35198 43370
rect 35198 43318 35250 43370
rect 35250 43318 35252 43370
rect 35196 43316 35252 43318
rect 35300 43370 35356 43372
rect 35300 43318 35302 43370
rect 35302 43318 35354 43370
rect 35354 43318 35356 43370
rect 35300 43316 35356 43318
rect 35404 43370 35460 43372
rect 35404 43318 35406 43370
rect 35406 43318 35458 43370
rect 35458 43318 35460 43370
rect 35404 43316 35460 43318
rect 37996 44940 38052 44996
rect 37996 43820 38052 43876
rect 36876 42924 36932 42980
rect 34972 40796 35028 40852
rect 35756 41916 35812 41972
rect 35532 41804 35588 41860
rect 35196 41354 35252 41356
rect 35196 41302 35198 41354
rect 35198 41302 35250 41354
rect 35250 41302 35252 41354
rect 35196 41300 35252 41302
rect 35300 41354 35356 41356
rect 35300 41302 35302 41354
rect 35302 41302 35354 41354
rect 35354 41302 35356 41354
rect 35300 41300 35356 41302
rect 35404 41354 35460 41356
rect 35404 41302 35406 41354
rect 35406 41302 35458 41354
rect 35458 41302 35460 41354
rect 35404 41300 35460 41302
rect 35196 40236 35252 40292
rect 34860 40124 34916 40180
rect 35084 40066 35140 40068
rect 35084 40014 35086 40066
rect 35086 40014 35138 40066
rect 35138 40014 35140 40066
rect 35084 40012 35140 40014
rect 36316 41916 36372 41972
rect 36428 41858 36484 41860
rect 36428 41806 36430 41858
rect 36430 41806 36482 41858
rect 36482 41806 36484 41858
rect 36428 41804 36484 41806
rect 36428 40850 36484 40852
rect 36428 40798 36430 40850
rect 36430 40798 36482 40850
rect 36482 40798 36484 40850
rect 36428 40796 36484 40798
rect 35980 40738 36036 40740
rect 35980 40686 35982 40738
rect 35982 40686 36034 40738
rect 36034 40686 36036 40738
rect 35980 40684 36036 40686
rect 37100 40460 37156 40516
rect 35980 40124 36036 40180
rect 36988 40236 37044 40292
rect 36540 39954 36596 39956
rect 36540 39902 36542 39954
rect 36542 39902 36594 39954
rect 36594 39902 36596 39954
rect 36540 39900 36596 39902
rect 35196 39338 35252 39340
rect 35196 39286 35198 39338
rect 35198 39286 35250 39338
rect 35250 39286 35252 39338
rect 35196 39284 35252 39286
rect 35300 39338 35356 39340
rect 35300 39286 35302 39338
rect 35302 39286 35354 39338
rect 35354 39286 35356 39338
rect 35300 39284 35356 39286
rect 35404 39338 35460 39340
rect 35404 39286 35406 39338
rect 35406 39286 35458 39338
rect 35458 39286 35460 39338
rect 35404 39284 35460 39286
rect 35532 38556 35588 38612
rect 36316 38556 36372 38612
rect 36316 37660 36372 37716
rect 35196 37322 35252 37324
rect 35196 37270 35198 37322
rect 35198 37270 35250 37322
rect 35250 37270 35252 37322
rect 35196 37268 35252 37270
rect 35300 37322 35356 37324
rect 35300 37270 35302 37322
rect 35302 37270 35354 37322
rect 35354 37270 35356 37322
rect 35300 37268 35356 37270
rect 35404 37322 35460 37324
rect 35404 37270 35406 37322
rect 35406 37270 35458 37322
rect 35458 37270 35460 37322
rect 35404 37268 35460 37270
rect 37772 42812 37828 42868
rect 38108 43762 38164 43764
rect 38108 43710 38110 43762
rect 38110 43710 38162 43762
rect 38162 43710 38164 43762
rect 38108 43708 38164 43710
rect 37772 41858 37828 41860
rect 37772 41806 37774 41858
rect 37774 41806 37826 41858
rect 37826 41806 37828 41858
rect 37772 41804 37828 41806
rect 37884 40738 37940 40740
rect 37884 40686 37886 40738
rect 37886 40686 37938 40738
rect 37938 40686 37940 40738
rect 37884 40684 37940 40686
rect 37324 39900 37380 39956
rect 37212 38780 37268 38836
rect 37324 39676 37380 39732
rect 37324 39004 37380 39060
rect 40124 46002 40180 46004
rect 40124 45950 40126 46002
rect 40126 45950 40178 46002
rect 40178 45950 40180 46002
rect 40124 45948 40180 45950
rect 39564 45500 39620 45556
rect 41020 46844 41076 46900
rect 42588 48802 42644 48804
rect 42588 48750 42590 48802
rect 42590 48750 42642 48802
rect 42642 48750 42644 48802
rect 42588 48748 42644 48750
rect 41356 48636 41412 48692
rect 43596 48748 43652 48804
rect 40348 45948 40404 46004
rect 40684 46786 40740 46788
rect 40684 46734 40686 46786
rect 40686 46734 40738 46786
rect 40738 46734 40740 46786
rect 40684 46732 40740 46734
rect 40236 45276 40292 45332
rect 41132 46002 41188 46004
rect 41132 45950 41134 46002
rect 41134 45950 41186 46002
rect 41186 45950 41188 46002
rect 41132 45948 41188 45950
rect 39452 43874 39508 43876
rect 39452 43822 39454 43874
rect 39454 43822 39506 43874
rect 39506 43822 39508 43874
rect 39452 43820 39508 43822
rect 39228 42924 39284 42980
rect 39564 43708 39620 43764
rect 40124 43484 40180 43540
rect 39676 42812 39732 42868
rect 39228 42754 39284 42756
rect 39228 42702 39230 42754
rect 39230 42702 39282 42754
rect 39282 42702 39284 42754
rect 39228 42700 39284 42702
rect 38892 41916 38948 41972
rect 38444 40850 38500 40852
rect 38444 40798 38446 40850
rect 38446 40798 38498 40850
rect 38498 40798 38500 40850
rect 38444 40796 38500 40798
rect 38780 40796 38836 40852
rect 37996 40460 38052 40516
rect 38444 40012 38500 40068
rect 37996 39842 38052 39844
rect 37996 39790 37998 39842
rect 37998 39790 38050 39842
rect 38050 39790 38052 39842
rect 37996 39788 38052 39790
rect 37660 37714 37716 37716
rect 37660 37662 37662 37714
rect 37662 37662 37714 37714
rect 37714 37662 37716 37714
rect 37660 37660 37716 37662
rect 37100 37548 37156 37604
rect 38220 37660 38276 37716
rect 36204 36034 36260 36036
rect 36204 35982 36206 36034
rect 36206 35982 36258 36034
rect 36258 35982 36260 36034
rect 36204 35980 36260 35982
rect 34748 35308 34804 35364
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35308 35138 35364 35140
rect 35308 35086 35310 35138
rect 35310 35086 35362 35138
rect 35362 35086 35364 35138
rect 35308 35084 35364 35086
rect 35644 35084 35700 35140
rect 35196 34802 35252 34804
rect 35196 34750 35198 34802
rect 35198 34750 35250 34802
rect 35250 34750 35252 34802
rect 35196 34748 35252 34750
rect 34860 34690 34916 34692
rect 34860 34638 34862 34690
rect 34862 34638 34914 34690
rect 34914 34638 34916 34690
rect 34860 34636 34916 34638
rect 35532 34636 35588 34692
rect 34300 33682 34356 33684
rect 34300 33630 34302 33682
rect 34302 33630 34354 33682
rect 34354 33630 34356 33682
rect 34300 33628 34356 33630
rect 34076 32620 34132 32676
rect 33516 31724 33572 31780
rect 33516 30604 33572 30660
rect 32844 30492 32900 30548
rect 32732 27244 32788 27300
rect 32508 26908 32564 26964
rect 32508 26460 32564 26516
rect 31612 23772 31668 23828
rect 31836 25452 31892 25508
rect 31276 22428 31332 22484
rect 29372 21420 29428 21476
rect 30380 21586 30436 21588
rect 30380 21534 30382 21586
rect 30382 21534 30434 21586
rect 30434 21534 30436 21586
rect 30380 21532 30436 21534
rect 30156 20300 30212 20356
rect 29708 20188 29764 20244
rect 28588 18562 28644 18564
rect 28588 18510 28590 18562
rect 28590 18510 28642 18562
rect 28642 18510 28644 18562
rect 28588 18508 28644 18510
rect 28364 17836 28420 17892
rect 28476 17724 28532 17780
rect 29596 17778 29652 17780
rect 29596 17726 29598 17778
rect 29598 17726 29650 17778
rect 29650 17726 29652 17778
rect 29596 17724 29652 17726
rect 28252 15708 28308 15764
rect 28924 16268 28980 16324
rect 29260 16492 29316 16548
rect 28364 15036 28420 15092
rect 27580 14700 27636 14756
rect 28252 14530 28308 14532
rect 28252 14478 28254 14530
rect 28254 14478 28306 14530
rect 28306 14478 28308 14530
rect 28252 14476 28308 14478
rect 29148 15820 29204 15876
rect 30268 20076 30324 20132
rect 31388 21532 31444 21588
rect 31724 20076 31780 20132
rect 30156 18786 30212 18788
rect 30156 18734 30158 18786
rect 30158 18734 30210 18786
rect 30210 18734 30212 18786
rect 30156 18732 30212 18734
rect 31724 19682 31780 19684
rect 31724 19630 31726 19682
rect 31726 19630 31778 19682
rect 31778 19630 31780 19682
rect 31724 19628 31780 19630
rect 31052 18620 31108 18676
rect 30044 18508 30100 18564
rect 30380 16322 30436 16324
rect 30380 16270 30382 16322
rect 30382 16270 30434 16322
rect 30434 16270 30436 16322
rect 30380 16268 30436 16270
rect 29708 15820 29764 15876
rect 29708 14418 29764 14420
rect 29708 14366 29710 14418
rect 29710 14366 29762 14418
rect 29762 14366 29764 14418
rect 29708 14364 29764 14366
rect 28588 13746 28644 13748
rect 28588 13694 28590 13746
rect 28590 13694 28642 13746
rect 28642 13694 28644 13746
rect 28588 13692 28644 13694
rect 29708 13692 29764 13748
rect 27244 13356 27300 13412
rect 27020 12738 27076 12740
rect 27020 12686 27022 12738
rect 27022 12686 27074 12738
rect 27074 12686 27076 12738
rect 27020 12684 27076 12686
rect 25900 11730 25956 11732
rect 25900 11678 25902 11730
rect 25902 11678 25954 11730
rect 25954 11678 25956 11730
rect 25900 11676 25956 11678
rect 25452 11618 25508 11620
rect 25452 11566 25454 11618
rect 25454 11566 25506 11618
rect 25506 11566 25508 11618
rect 25452 11564 25508 11566
rect 26012 9996 26068 10052
rect 25676 9826 25732 9828
rect 25676 9774 25678 9826
rect 25678 9774 25730 9826
rect 25730 9774 25732 9826
rect 25676 9772 25732 9774
rect 25228 9660 25284 9716
rect 27132 11676 27188 11732
rect 28812 11564 28868 11620
rect 26796 9996 26852 10052
rect 26572 9660 26628 9716
rect 28140 9660 28196 9716
rect 28140 8706 28196 8708
rect 28140 8654 28142 8706
rect 28142 8654 28194 8706
rect 28194 8654 28196 8706
rect 28140 8652 28196 8654
rect 31500 18508 31556 18564
rect 30828 16546 30884 16548
rect 30828 16494 30830 16546
rect 30830 16494 30882 16546
rect 30882 16494 30884 16546
rect 30828 16492 30884 16494
rect 31500 16716 31556 16772
rect 30604 15372 30660 15428
rect 31276 15986 31332 15988
rect 31276 15934 31278 15986
rect 31278 15934 31330 15986
rect 31330 15934 31332 15986
rect 31276 15932 31332 15934
rect 30940 15484 30996 15540
rect 30492 14364 30548 14420
rect 31276 15372 31332 15428
rect 31500 15036 31556 15092
rect 30940 14418 30996 14420
rect 30940 14366 30942 14418
rect 30942 14366 30994 14418
rect 30994 14366 30996 14418
rect 30940 14364 30996 14366
rect 30380 13356 30436 13412
rect 29820 11618 29876 11620
rect 29820 11566 29822 11618
rect 29822 11566 29874 11618
rect 29874 11566 29876 11618
rect 29820 11564 29876 11566
rect 29484 11340 29540 11396
rect 21308 7756 21364 7812
rect 22316 7810 22372 7812
rect 22316 7758 22318 7810
rect 22318 7758 22370 7810
rect 22370 7758 22372 7810
rect 22316 7756 22372 7758
rect 28588 8594 28644 8596
rect 28588 8542 28590 8594
rect 28590 8542 28642 8594
rect 28642 8542 28644 8594
rect 28588 8540 28644 8542
rect 27692 8482 27748 8484
rect 27692 8430 27694 8482
rect 27694 8430 27746 8482
rect 27746 8430 27748 8482
rect 27692 8428 27748 8430
rect 28700 8428 28756 8484
rect 29708 9996 29764 10052
rect 29148 8652 29204 8708
rect 24892 7756 24948 7812
rect 28252 7810 28308 7812
rect 28252 7758 28254 7810
rect 28254 7758 28306 7810
rect 28306 7758 28308 7810
rect 28252 7756 28308 7758
rect 29596 8652 29652 8708
rect 29260 8594 29316 8596
rect 29260 8542 29262 8594
rect 29262 8542 29314 8594
rect 29314 8542 29316 8594
rect 29260 8540 29316 8542
rect 30828 11676 30884 11732
rect 30380 11564 30436 11620
rect 30380 10722 30436 10724
rect 30380 10670 30382 10722
rect 30382 10670 30434 10722
rect 30434 10670 30436 10722
rect 30380 10668 30436 10670
rect 31612 12684 31668 12740
rect 32508 25058 32564 25060
rect 32508 25006 32510 25058
rect 32510 25006 32562 25058
rect 32562 25006 32564 25058
rect 32508 25004 32564 25006
rect 31948 24780 32004 24836
rect 32620 24722 32676 24724
rect 32620 24670 32622 24722
rect 32622 24670 32674 24722
rect 32674 24670 32676 24722
rect 32620 24668 32676 24670
rect 35308 33628 35364 33684
rect 35196 33290 35252 33292
rect 35196 33238 35198 33290
rect 35198 33238 35250 33290
rect 35250 33238 35252 33290
rect 35196 33236 35252 33238
rect 35300 33290 35356 33292
rect 35300 33238 35302 33290
rect 35302 33238 35354 33290
rect 35354 33238 35356 33290
rect 35300 33236 35356 33238
rect 35404 33290 35460 33292
rect 35404 33238 35406 33290
rect 35406 33238 35458 33290
rect 35458 33238 35460 33290
rect 35404 33236 35460 33238
rect 35532 32674 35588 32676
rect 35532 32622 35534 32674
rect 35534 32622 35586 32674
rect 35586 32622 35588 32674
rect 35532 32620 35588 32622
rect 34636 31836 34692 31892
rect 33852 31164 33908 31220
rect 33740 30882 33796 30884
rect 33740 30830 33742 30882
rect 33742 30830 33794 30882
rect 33794 30830 33796 30882
rect 33740 30828 33796 30830
rect 33628 30492 33684 30548
rect 36204 34748 36260 34804
rect 37100 35922 37156 35924
rect 37100 35870 37102 35922
rect 37102 35870 37154 35922
rect 37154 35870 37156 35922
rect 37100 35868 37156 35870
rect 37772 36706 37828 36708
rect 37772 36654 37774 36706
rect 37774 36654 37826 36706
rect 37826 36654 37828 36706
rect 37772 36652 37828 36654
rect 37772 35980 37828 36036
rect 38332 35868 38388 35924
rect 37212 34802 37268 34804
rect 37212 34750 37214 34802
rect 37214 34750 37266 34802
rect 37266 34750 37268 34802
rect 37212 34748 37268 34750
rect 35644 31836 35700 31892
rect 35756 32956 35812 33012
rect 33964 30156 34020 30212
rect 34188 30492 34244 30548
rect 33852 29874 33908 29876
rect 33852 29822 33854 29874
rect 33854 29822 33906 29874
rect 33906 29822 33908 29874
rect 33852 29820 33908 29822
rect 33628 29708 33684 29764
rect 34300 30268 34356 30324
rect 34748 30268 34804 30324
rect 35644 31500 35700 31556
rect 35196 31274 35252 31276
rect 35196 31222 35198 31274
rect 35198 31222 35250 31274
rect 35250 31222 35252 31274
rect 35196 31220 35252 31222
rect 35300 31274 35356 31276
rect 35300 31222 35302 31274
rect 35302 31222 35354 31274
rect 35354 31222 35356 31274
rect 35300 31220 35356 31222
rect 35404 31274 35460 31276
rect 35404 31222 35406 31274
rect 35406 31222 35458 31274
rect 35458 31222 35460 31274
rect 35404 31220 35460 31222
rect 34972 30828 35028 30884
rect 35084 30546 35140 30548
rect 35084 30494 35086 30546
rect 35086 30494 35138 30546
rect 35138 30494 35140 30546
rect 35084 30492 35140 30494
rect 34748 29708 34804 29764
rect 34972 30380 35028 30436
rect 33852 29650 33908 29652
rect 33852 29598 33854 29650
rect 33854 29598 33906 29650
rect 33906 29598 33908 29650
rect 33852 29596 33908 29598
rect 35084 30268 35140 30324
rect 33180 29484 33236 29540
rect 32956 28700 33012 28756
rect 33292 28476 33348 28532
rect 33516 28588 33572 28644
rect 33404 27858 33460 27860
rect 33404 27806 33406 27858
rect 33406 27806 33458 27858
rect 33458 27806 33460 27858
rect 33404 27804 33460 27806
rect 33404 27356 33460 27412
rect 33292 27020 33348 27076
rect 33068 26738 33124 26740
rect 33068 26686 33070 26738
rect 33070 26686 33122 26738
rect 33122 26686 33124 26738
rect 33068 26684 33124 26686
rect 32060 23548 32116 23604
rect 32620 23548 32676 23604
rect 32508 22482 32564 22484
rect 32508 22430 32510 22482
rect 32510 22430 32562 22482
rect 32562 22430 32564 22482
rect 32508 22428 32564 22430
rect 32060 20076 32116 20132
rect 32172 19570 32228 19572
rect 32172 19518 32174 19570
rect 32174 19518 32226 19570
rect 32226 19518 32228 19570
rect 32172 19516 32228 19518
rect 31948 16716 32004 16772
rect 32956 23772 33012 23828
rect 33292 23660 33348 23716
rect 33292 22428 33348 22484
rect 33740 27580 33796 27636
rect 38108 34802 38164 34804
rect 38108 34750 38110 34802
rect 38110 34750 38162 34802
rect 38162 34750 38164 34802
rect 38108 34748 38164 34750
rect 37660 34524 37716 34580
rect 37212 33852 37268 33908
rect 37100 32674 37156 32676
rect 37100 32622 37102 32674
rect 37102 32622 37154 32674
rect 37154 32622 37156 32674
rect 37100 32620 37156 32622
rect 37324 32508 37380 32564
rect 36652 31778 36708 31780
rect 36652 31726 36654 31778
rect 36654 31726 36706 31778
rect 36706 31726 36708 31778
rect 36652 31724 36708 31726
rect 35756 31052 35812 31108
rect 36988 31554 37044 31556
rect 36988 31502 36990 31554
rect 36990 31502 37042 31554
rect 37042 31502 37044 31554
rect 36988 31500 37044 31502
rect 36652 30940 36708 30996
rect 36428 30716 36484 30772
rect 35420 30156 35476 30212
rect 36092 29932 36148 29988
rect 36204 30380 36260 30436
rect 35196 29258 35252 29260
rect 35196 29206 35198 29258
rect 35198 29206 35250 29258
rect 35250 29206 35252 29258
rect 35196 29204 35252 29206
rect 35300 29258 35356 29260
rect 35300 29206 35302 29258
rect 35302 29206 35354 29258
rect 35354 29206 35356 29258
rect 35300 29204 35356 29206
rect 35404 29258 35460 29260
rect 35404 29206 35406 29258
rect 35406 29206 35458 29258
rect 35458 29206 35460 29258
rect 35404 29204 35460 29206
rect 34748 28924 34804 28980
rect 34300 28754 34356 28756
rect 34300 28702 34302 28754
rect 34302 28702 34354 28754
rect 34354 28702 34356 28754
rect 34300 28700 34356 28702
rect 34524 28588 34580 28644
rect 33740 26738 33796 26740
rect 33740 26686 33742 26738
rect 33742 26686 33794 26738
rect 33794 26686 33796 26738
rect 33740 26684 33796 26686
rect 33628 25506 33684 25508
rect 33628 25454 33630 25506
rect 33630 25454 33682 25506
rect 33682 25454 33684 25506
rect 33628 25452 33684 25454
rect 33852 25340 33908 25396
rect 34412 27580 34468 27636
rect 35532 28140 35588 28196
rect 35644 28028 35700 28084
rect 35980 29708 36036 29764
rect 37324 30940 37380 30996
rect 36988 30882 37044 30884
rect 36988 30830 36990 30882
rect 36990 30830 37042 30882
rect 37042 30830 37044 30882
rect 36988 30828 37044 30830
rect 36652 30268 36708 30324
rect 37324 30268 37380 30324
rect 37100 29932 37156 29988
rect 35980 29372 36036 29428
rect 36204 29260 36260 29316
rect 36764 29650 36820 29652
rect 36764 29598 36766 29650
rect 36766 29598 36818 29650
rect 36818 29598 36820 29650
rect 36764 29596 36820 29598
rect 37772 31666 37828 31668
rect 37772 31614 37774 31666
rect 37774 31614 37826 31666
rect 37826 31614 37828 31666
rect 37772 31612 37828 31614
rect 38332 35532 38388 35588
rect 38332 33964 38388 34020
rect 39788 41916 39844 41972
rect 39564 40796 39620 40852
rect 39228 40012 39284 40068
rect 38780 39564 38836 39620
rect 39676 40460 39732 40516
rect 39788 39900 39844 39956
rect 39788 39730 39844 39732
rect 39788 39678 39790 39730
rect 39790 39678 39842 39730
rect 39842 39678 39844 39730
rect 39788 39676 39844 39678
rect 39452 39004 39508 39060
rect 38556 38892 38612 38948
rect 39116 38834 39172 38836
rect 39116 38782 39118 38834
rect 39118 38782 39170 38834
rect 39170 38782 39172 38834
rect 39116 38780 39172 38782
rect 39452 38780 39508 38836
rect 38556 37884 38612 37940
rect 38892 37938 38948 37940
rect 38892 37886 38894 37938
rect 38894 37886 38946 37938
rect 38946 37886 38948 37938
rect 38892 37884 38948 37886
rect 38556 37548 38612 37604
rect 40348 43762 40404 43764
rect 40348 43710 40350 43762
rect 40350 43710 40402 43762
rect 40402 43710 40404 43762
rect 40348 43708 40404 43710
rect 50556 48410 50612 48412
rect 50556 48358 50558 48410
rect 50558 48358 50610 48410
rect 50610 48358 50612 48410
rect 50556 48356 50612 48358
rect 50660 48410 50716 48412
rect 50660 48358 50662 48410
rect 50662 48358 50714 48410
rect 50714 48358 50716 48410
rect 50660 48356 50716 48358
rect 50764 48410 50820 48412
rect 50764 48358 50766 48410
rect 50766 48358 50818 48410
rect 50818 48358 50820 48410
rect 50764 48356 50820 48358
rect 43372 46620 43428 46676
rect 42812 45948 42868 46004
rect 42140 45388 42196 45444
rect 41020 43762 41076 43764
rect 41020 43710 41022 43762
rect 41022 43710 41074 43762
rect 41074 43710 41076 43762
rect 41020 43708 41076 43710
rect 41468 43762 41524 43764
rect 41468 43710 41470 43762
rect 41470 43710 41522 43762
rect 41522 43710 41524 43762
rect 41468 43708 41524 43710
rect 40796 43484 40852 43540
rect 40236 42700 40292 42756
rect 41020 42812 41076 42868
rect 40348 40684 40404 40740
rect 40236 40012 40292 40068
rect 40236 39004 40292 39060
rect 40236 38668 40292 38724
rect 38556 36652 38612 36708
rect 38892 36428 38948 36484
rect 38668 34802 38724 34804
rect 38668 34750 38670 34802
rect 38670 34750 38722 34802
rect 38722 34750 38724 34802
rect 38668 34748 38724 34750
rect 40124 35532 40180 35588
rect 39788 32786 39844 32788
rect 39788 32734 39790 32786
rect 39790 32734 39842 32786
rect 39842 32734 39844 32786
rect 39788 32732 39844 32734
rect 38220 31612 38276 31668
rect 38892 32620 38948 32676
rect 37548 30546 37604 30548
rect 37548 30494 37550 30546
rect 37550 30494 37602 30546
rect 37602 30494 37604 30546
rect 37548 30492 37604 30494
rect 37996 30716 38052 30772
rect 37772 30268 37828 30324
rect 36652 29260 36708 29316
rect 36428 28924 36484 28980
rect 35980 28642 36036 28644
rect 35980 28590 35982 28642
rect 35982 28590 36034 28642
rect 36034 28590 36036 28642
rect 35980 28588 36036 28590
rect 37548 29932 37604 29988
rect 37100 28866 37156 28868
rect 37100 28814 37102 28866
rect 37102 28814 37154 28866
rect 37154 28814 37156 28866
rect 37100 28812 37156 28814
rect 36540 28364 36596 28420
rect 36316 27858 36372 27860
rect 36316 27806 36318 27858
rect 36318 27806 36370 27858
rect 36370 27806 36372 27858
rect 36316 27804 36372 27806
rect 34188 26572 34244 26628
rect 35644 27356 35700 27412
rect 35196 27242 35252 27244
rect 35196 27190 35198 27242
rect 35198 27190 35250 27242
rect 35250 27190 35252 27242
rect 35196 27188 35252 27190
rect 35300 27242 35356 27244
rect 35300 27190 35302 27242
rect 35302 27190 35354 27242
rect 35354 27190 35356 27242
rect 35300 27188 35356 27190
rect 35404 27242 35460 27244
rect 35404 27190 35406 27242
rect 35406 27190 35458 27242
rect 35458 27190 35460 27242
rect 35404 27188 35460 27190
rect 34748 26572 34804 26628
rect 35980 27580 36036 27636
rect 36540 27356 36596 27412
rect 33964 24780 34020 24836
rect 33740 23714 33796 23716
rect 33740 23662 33742 23714
rect 33742 23662 33794 23714
rect 33794 23662 33796 23714
rect 33740 23660 33796 23662
rect 35532 25842 35588 25844
rect 35532 25790 35534 25842
rect 35534 25790 35586 25842
rect 35586 25790 35588 25842
rect 35532 25788 35588 25790
rect 34524 25004 34580 25060
rect 34860 25340 34916 25396
rect 34524 24498 34580 24500
rect 34524 24446 34526 24498
rect 34526 24446 34578 24498
rect 34578 24446 34580 24498
rect 34524 24444 34580 24446
rect 34076 23548 34132 23604
rect 35196 25226 35252 25228
rect 35196 25174 35198 25226
rect 35198 25174 35250 25226
rect 35250 25174 35252 25226
rect 35196 25172 35252 25174
rect 35300 25226 35356 25228
rect 35300 25174 35302 25226
rect 35302 25174 35354 25226
rect 35354 25174 35356 25226
rect 35300 25172 35356 25174
rect 35404 25226 35460 25228
rect 35404 25174 35406 25226
rect 35406 25174 35458 25226
rect 35458 25174 35460 25226
rect 35404 25172 35460 25174
rect 35196 25004 35252 25060
rect 35644 24780 35700 24836
rect 35980 26012 36036 26068
rect 35420 24444 35476 24500
rect 35868 24108 35924 24164
rect 35196 23660 35252 23716
rect 35196 23210 35252 23212
rect 35196 23158 35198 23210
rect 35198 23158 35250 23210
rect 35250 23158 35252 23210
rect 35196 23156 35252 23158
rect 35300 23210 35356 23212
rect 35300 23158 35302 23210
rect 35302 23158 35354 23210
rect 35354 23158 35356 23210
rect 35300 23156 35356 23158
rect 35404 23210 35460 23212
rect 35404 23158 35406 23210
rect 35406 23158 35458 23210
rect 35458 23158 35460 23210
rect 35404 23156 35460 23158
rect 34412 22764 34468 22820
rect 36540 26348 36596 26404
rect 36988 27580 37044 27636
rect 37436 28642 37492 28644
rect 37436 28590 37438 28642
rect 37438 28590 37490 28642
rect 37490 28590 37492 28642
rect 37436 28588 37492 28590
rect 38444 31724 38500 31780
rect 38556 31666 38612 31668
rect 38556 31614 38558 31666
rect 38558 31614 38610 31666
rect 38610 31614 38612 31666
rect 38556 31612 38612 31614
rect 38556 30940 38612 30996
rect 38108 30434 38164 30436
rect 38108 30382 38110 30434
rect 38110 30382 38162 30434
rect 38162 30382 38164 30434
rect 38108 30380 38164 30382
rect 37884 29932 37940 29988
rect 38332 29874 38388 29876
rect 38332 29822 38334 29874
rect 38334 29822 38386 29874
rect 38386 29822 38388 29874
rect 38332 29820 38388 29822
rect 37884 29762 37940 29764
rect 37884 29710 37886 29762
rect 37886 29710 37938 29762
rect 37938 29710 37940 29762
rect 37884 29708 37940 29710
rect 38556 30492 38612 30548
rect 39004 31836 39060 31892
rect 39900 31612 39956 31668
rect 39004 30828 39060 30884
rect 37996 28530 38052 28532
rect 37996 28478 37998 28530
rect 37998 28478 38050 28530
rect 38050 28478 38052 28530
rect 37996 28476 38052 28478
rect 37884 28028 37940 28084
rect 36764 26012 36820 26068
rect 37212 26796 37268 26852
rect 37100 26738 37156 26740
rect 37100 26686 37102 26738
rect 37102 26686 37154 26738
rect 37154 26686 37156 26738
rect 37100 26684 37156 26686
rect 36204 24892 36260 24948
rect 36540 24780 36596 24836
rect 36988 25228 37044 25284
rect 36764 24892 36820 24948
rect 37212 24332 37268 24388
rect 36764 24108 36820 24164
rect 37548 26460 37604 26516
rect 37772 27356 37828 27412
rect 37772 26012 37828 26068
rect 38444 27634 38500 27636
rect 38444 27582 38446 27634
rect 38446 27582 38498 27634
rect 38498 27582 38500 27634
rect 38444 27580 38500 27582
rect 38668 28364 38724 28420
rect 38556 27356 38612 27412
rect 38668 27804 38724 27860
rect 38892 27692 38948 27748
rect 39452 30658 39508 30660
rect 39452 30606 39454 30658
rect 39454 30606 39506 30658
rect 39506 30606 39508 30658
rect 39452 30604 39508 30606
rect 39228 30492 39284 30548
rect 39788 30156 39844 30212
rect 39676 29596 39732 29652
rect 39788 29036 39844 29092
rect 39452 28476 39508 28532
rect 40460 39676 40516 39732
rect 41244 42812 41300 42868
rect 41244 41916 41300 41972
rect 41692 41916 41748 41972
rect 42588 45276 42644 45332
rect 43820 46732 43876 46788
rect 44044 46674 44100 46676
rect 44044 46622 44046 46674
rect 44046 46622 44098 46674
rect 44098 46622 44100 46674
rect 44044 46620 44100 46622
rect 43708 46172 43764 46228
rect 43932 46060 43988 46116
rect 43372 45500 43428 45556
rect 42700 44044 42756 44100
rect 42588 42866 42644 42868
rect 42588 42814 42590 42866
rect 42590 42814 42642 42866
rect 42642 42814 42644 42866
rect 42588 42812 42644 42814
rect 43260 43708 43316 43764
rect 42812 43036 42868 43092
rect 43036 43260 43092 43316
rect 41916 42642 41972 42644
rect 41916 42590 41918 42642
rect 41918 42590 41970 42642
rect 41970 42590 41972 42642
rect 41916 42588 41972 42590
rect 42700 42588 42756 42644
rect 42364 42476 42420 42532
rect 41356 41746 41412 41748
rect 41356 41694 41358 41746
rect 41358 41694 41410 41746
rect 41410 41694 41412 41746
rect 41356 41692 41412 41694
rect 41468 41522 41524 41524
rect 41468 41470 41470 41522
rect 41470 41470 41522 41522
rect 41522 41470 41524 41522
rect 41468 41468 41524 41470
rect 43260 42812 43316 42868
rect 43148 42588 43204 42644
rect 42140 41692 42196 41748
rect 41356 40684 41412 40740
rect 44044 46172 44100 46228
rect 43708 44882 43764 44884
rect 43708 44830 43710 44882
rect 43710 44830 43762 44882
rect 43762 44830 43764 44882
rect 43708 44828 43764 44830
rect 43484 44268 43540 44324
rect 43484 44098 43540 44100
rect 43484 44046 43486 44098
rect 43486 44046 43538 44098
rect 43538 44046 43540 44098
rect 43484 44044 43540 44046
rect 43596 43148 43652 43204
rect 43596 42866 43652 42868
rect 43596 42814 43598 42866
rect 43598 42814 43650 42866
rect 43650 42814 43652 42866
rect 43596 42812 43652 42814
rect 45164 46172 45220 46228
rect 46172 46114 46228 46116
rect 46172 46062 46174 46114
rect 46174 46062 46226 46114
rect 46226 46062 46228 46114
rect 46172 46060 46228 46062
rect 44044 44828 44100 44884
rect 43932 44268 43988 44324
rect 48076 45836 48132 45892
rect 44716 44828 44772 44884
rect 44156 44716 44212 44772
rect 45052 44770 45108 44772
rect 45052 44718 45054 44770
rect 45054 44718 45106 44770
rect 45106 44718 45108 44770
rect 45052 44716 45108 44718
rect 44156 44044 44212 44100
rect 43932 43596 43988 43652
rect 46620 44716 46676 44772
rect 45164 43596 45220 43652
rect 44940 43260 44996 43316
rect 45164 43148 45220 43204
rect 44716 42530 44772 42532
rect 44716 42478 44718 42530
rect 44718 42478 44770 42530
rect 44770 42478 44772 42530
rect 44716 42476 44772 42478
rect 45388 43036 45444 43092
rect 44604 41858 44660 41860
rect 44604 41806 44606 41858
rect 44606 41806 44658 41858
rect 44658 41806 44660 41858
rect 44604 41804 44660 41806
rect 41916 40012 41972 40068
rect 42028 40460 42084 40516
rect 41020 39788 41076 39844
rect 41468 39842 41524 39844
rect 41468 39790 41470 39842
rect 41470 39790 41522 39842
rect 41522 39790 41524 39842
rect 41468 39788 41524 39790
rect 42140 39788 42196 39844
rect 40572 38892 40628 38948
rect 40460 37884 40516 37940
rect 40348 35810 40404 35812
rect 40348 35758 40350 35810
rect 40350 35758 40402 35810
rect 40402 35758 40404 35810
rect 40348 35756 40404 35758
rect 40348 34018 40404 34020
rect 40348 33966 40350 34018
rect 40350 33966 40402 34018
rect 40402 33966 40404 34018
rect 40348 33964 40404 33966
rect 40796 38780 40852 38836
rect 41132 38722 41188 38724
rect 41132 38670 41134 38722
rect 41134 38670 41186 38722
rect 41186 38670 41188 38722
rect 41132 38668 41188 38670
rect 41244 36988 41300 37044
rect 41356 37548 41412 37604
rect 41244 36706 41300 36708
rect 41244 36654 41246 36706
rect 41246 36654 41298 36706
rect 41298 36654 41300 36706
rect 41244 36652 41300 36654
rect 41244 35810 41300 35812
rect 41244 35758 41246 35810
rect 41246 35758 41298 35810
rect 41298 35758 41300 35810
rect 41244 35756 41300 35758
rect 41580 37996 41636 38052
rect 42140 39564 42196 39620
rect 41916 38892 41972 38948
rect 42476 39676 42532 39732
rect 42364 38892 42420 38948
rect 41468 36428 41524 36484
rect 41692 35698 41748 35700
rect 41692 35646 41694 35698
rect 41694 35646 41746 35698
rect 41746 35646 41748 35698
rect 41692 35644 41748 35646
rect 41020 33852 41076 33908
rect 40572 32620 40628 32676
rect 40460 32562 40516 32564
rect 40460 32510 40462 32562
rect 40462 32510 40514 32562
rect 40514 32510 40516 32562
rect 40460 32508 40516 32510
rect 41356 33628 41412 33684
rect 41020 32674 41076 32676
rect 41020 32622 41022 32674
rect 41022 32622 41074 32674
rect 41074 32622 41076 32674
rect 41020 32620 41076 32622
rect 41244 31836 41300 31892
rect 40908 31612 40964 31668
rect 40572 30716 40628 30772
rect 41132 30716 41188 30772
rect 40236 30156 40292 30212
rect 40908 29874 40964 29876
rect 40908 29822 40910 29874
rect 40910 29822 40962 29874
rect 40962 29822 40964 29874
rect 40908 29820 40964 29822
rect 40348 29650 40404 29652
rect 40348 29598 40350 29650
rect 40350 29598 40402 29650
rect 40402 29598 40404 29650
rect 40348 29596 40404 29598
rect 42364 35644 42420 35700
rect 42588 38722 42644 38724
rect 42588 38670 42590 38722
rect 42590 38670 42642 38722
rect 42642 38670 42644 38722
rect 42588 38668 42644 38670
rect 41804 35196 41860 35252
rect 41804 34578 41860 34580
rect 41804 34526 41806 34578
rect 41806 34526 41858 34578
rect 41858 34526 41860 34578
rect 41804 34524 41860 34526
rect 42252 33852 42308 33908
rect 42364 33740 42420 33796
rect 42028 32508 42084 32564
rect 43596 40460 43652 40516
rect 43596 40124 43652 40180
rect 43932 40236 43988 40292
rect 42700 37548 42756 37604
rect 43036 37996 43092 38052
rect 42588 36876 42644 36932
rect 43260 37938 43316 37940
rect 43260 37886 43262 37938
rect 43262 37886 43314 37938
rect 43314 37886 43316 37938
rect 43260 37884 43316 37886
rect 42700 35756 42756 35812
rect 45612 42754 45668 42756
rect 45612 42702 45614 42754
rect 45614 42702 45666 42754
rect 45666 42702 45668 42754
rect 45612 42700 45668 42702
rect 47404 43596 47460 43652
rect 46396 42866 46452 42868
rect 46396 42814 46398 42866
rect 46398 42814 46450 42866
rect 46450 42814 46452 42866
rect 46396 42812 46452 42814
rect 46844 42642 46900 42644
rect 46844 42590 46846 42642
rect 46846 42590 46898 42642
rect 46898 42590 46900 42642
rect 46844 42588 46900 42590
rect 47628 42812 47684 42868
rect 47404 42588 47460 42644
rect 49420 45890 49476 45892
rect 49420 45838 49422 45890
rect 49422 45838 49474 45890
rect 49474 45838 49476 45890
rect 49420 45836 49476 45838
rect 49756 45388 49812 45444
rect 50092 45388 50148 45444
rect 49084 45276 49140 45332
rect 49644 44604 49700 44660
rect 48636 43708 48692 43764
rect 49532 43762 49588 43764
rect 49532 43710 49534 43762
rect 49534 43710 49586 43762
rect 49586 43710 49588 43762
rect 49532 43708 49588 43710
rect 48188 42642 48244 42644
rect 48188 42590 48190 42642
rect 48190 42590 48242 42642
rect 48242 42590 48244 42642
rect 48188 42588 48244 42590
rect 49756 42812 49812 42868
rect 49084 42028 49140 42084
rect 49420 42588 49476 42644
rect 46620 41858 46676 41860
rect 46620 41806 46622 41858
rect 46622 41806 46674 41858
rect 46674 41806 46676 41858
rect 46620 41804 46676 41806
rect 47964 40850 48020 40852
rect 47964 40798 47966 40850
rect 47966 40798 48018 40850
rect 48018 40798 48020 40850
rect 47964 40796 48020 40798
rect 49420 40796 49476 40852
rect 47068 40738 47124 40740
rect 47068 40686 47070 40738
rect 47070 40686 47122 40738
rect 47122 40686 47124 40738
rect 47068 40684 47124 40686
rect 47740 40738 47796 40740
rect 47740 40686 47742 40738
rect 47742 40686 47794 40738
rect 47794 40686 47796 40738
rect 47740 40684 47796 40686
rect 45500 40236 45556 40292
rect 44940 40124 44996 40180
rect 44492 40066 44548 40068
rect 44492 40014 44494 40066
rect 44494 40014 44546 40066
rect 44546 40014 44548 40066
rect 44492 40012 44548 40014
rect 44044 39730 44100 39732
rect 44044 39678 44046 39730
rect 44046 39678 44098 39730
rect 44098 39678 44100 39730
rect 44044 39676 44100 39678
rect 45276 40124 45332 40180
rect 44604 38780 44660 38836
rect 46396 40124 46452 40180
rect 45388 40066 45444 40068
rect 45388 40014 45390 40066
rect 45390 40014 45442 40066
rect 45442 40014 45444 40066
rect 45388 40012 45444 40014
rect 44940 38722 44996 38724
rect 44940 38670 44942 38722
rect 44942 38670 44994 38722
rect 44994 38670 44996 38722
rect 44940 38668 44996 38670
rect 46396 37996 46452 38052
rect 46508 40012 46564 40068
rect 46508 38668 46564 38724
rect 46732 39676 46788 39732
rect 43708 35308 43764 35364
rect 42924 34524 42980 34580
rect 42588 32508 42644 32564
rect 41132 29484 41188 29540
rect 41132 28812 41188 28868
rect 39788 27746 39844 27748
rect 39788 27694 39790 27746
rect 39790 27694 39842 27746
rect 39842 27694 39844 27746
rect 39788 27692 39844 27694
rect 39116 26796 39172 26852
rect 38780 26684 38836 26740
rect 38332 26348 38388 26404
rect 38444 26460 38500 26516
rect 37996 26012 38052 26068
rect 37548 25340 37604 25396
rect 36204 23660 36260 23716
rect 35756 22876 35812 22932
rect 35084 22594 35140 22596
rect 35084 22542 35086 22594
rect 35086 22542 35138 22594
rect 35138 22542 35140 22594
rect 35084 22540 35140 22542
rect 33180 21586 33236 21588
rect 33180 21534 33182 21586
rect 33182 21534 33234 21586
rect 33234 21534 33236 21586
rect 33180 21532 33236 21534
rect 33180 19964 33236 20020
rect 32508 18620 32564 18676
rect 32172 17612 32228 17668
rect 32508 17500 32564 17556
rect 32284 16492 32340 16548
rect 31948 15260 32004 15316
rect 32060 15596 32116 15652
rect 32956 15650 33012 15652
rect 32956 15598 32958 15650
rect 32958 15598 33010 15650
rect 33010 15598 33012 15650
rect 32956 15596 33012 15598
rect 33628 21922 33684 21924
rect 33628 21870 33630 21922
rect 33630 21870 33682 21922
rect 33682 21870 33684 21922
rect 33628 21868 33684 21870
rect 34748 21868 34804 21924
rect 33404 19852 33460 19908
rect 32396 15260 32452 15316
rect 33180 15484 33236 15540
rect 32396 14700 32452 14756
rect 32508 15036 32564 15092
rect 33180 14924 33236 14980
rect 33292 14700 33348 14756
rect 35532 21868 35588 21924
rect 34860 21532 34916 21588
rect 38332 25788 38388 25844
rect 38108 24332 38164 24388
rect 38668 25900 38724 25956
rect 39004 26460 39060 26516
rect 38892 26348 38948 26404
rect 40012 27858 40068 27860
rect 40012 27806 40014 27858
rect 40014 27806 40066 27858
rect 40066 27806 40068 27858
rect 40012 27804 40068 27806
rect 41692 28588 41748 28644
rect 43148 34578 43204 34580
rect 43148 34526 43150 34578
rect 43150 34526 43202 34578
rect 43202 34526 43204 34578
rect 43148 34524 43204 34526
rect 43484 33740 43540 33796
rect 44044 35308 44100 35364
rect 45164 36706 45220 36708
rect 45164 36654 45166 36706
rect 45166 36654 45218 36706
rect 45218 36654 45220 36706
rect 45164 36652 45220 36654
rect 46732 36540 46788 36596
rect 44492 35698 44548 35700
rect 44492 35646 44494 35698
rect 44494 35646 44546 35698
rect 44546 35646 44548 35698
rect 44492 35644 44548 35646
rect 44940 35308 44996 35364
rect 44380 35196 44436 35252
rect 44268 35084 44324 35140
rect 44828 35084 44884 35140
rect 44044 34914 44100 34916
rect 44044 34862 44046 34914
rect 44046 34862 44098 34914
rect 44098 34862 44100 34914
rect 44044 34860 44100 34862
rect 44716 34860 44772 34916
rect 44492 34636 44548 34692
rect 44268 33794 44324 33796
rect 44268 33742 44270 33794
rect 44270 33742 44322 33794
rect 44322 33742 44324 33794
rect 44268 33740 44324 33742
rect 43708 33628 43764 33684
rect 42140 31836 42196 31892
rect 43932 32732 43988 32788
rect 44716 34018 44772 34020
rect 44716 33966 44718 34018
rect 44718 33966 44770 34018
rect 44770 33966 44772 34018
rect 44716 33964 44772 33966
rect 44940 34914 44996 34916
rect 44940 34862 44942 34914
rect 44942 34862 44994 34914
rect 44994 34862 44996 34914
rect 44940 34860 44996 34862
rect 45836 35308 45892 35364
rect 45724 33794 45780 33796
rect 45724 33742 45726 33794
rect 45726 33742 45778 33794
rect 45778 33742 45780 33794
rect 45724 33740 45780 33742
rect 45164 33628 45220 33684
rect 43036 31836 43092 31892
rect 42140 29372 42196 29428
rect 42028 28476 42084 28532
rect 41692 27916 41748 27972
rect 39900 26684 39956 26740
rect 40012 26796 40068 26852
rect 39116 25900 39172 25956
rect 39228 26012 39284 26068
rect 39564 26460 39620 26516
rect 39564 25116 39620 25172
rect 40348 27634 40404 27636
rect 40348 27582 40350 27634
rect 40350 27582 40402 27634
rect 40402 27582 40404 27634
rect 40348 27580 40404 27582
rect 40348 26572 40404 26628
rect 37884 23714 37940 23716
rect 37884 23662 37886 23714
rect 37886 23662 37938 23714
rect 37938 23662 37940 23714
rect 37884 23660 37940 23662
rect 36988 22930 37044 22932
rect 36988 22878 36990 22930
rect 36990 22878 37042 22930
rect 37042 22878 37044 22930
rect 36988 22876 37044 22878
rect 36092 22594 36148 22596
rect 36092 22542 36094 22594
rect 36094 22542 36146 22594
rect 36146 22542 36148 22594
rect 36092 22540 36148 22542
rect 35644 21644 35700 21700
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34188 19964 34244 20020
rect 34524 19906 34580 19908
rect 34524 19854 34526 19906
rect 34526 19854 34578 19906
rect 34578 19854 34580 19906
rect 34524 19852 34580 19854
rect 34188 19794 34244 19796
rect 34188 19742 34190 19794
rect 34190 19742 34242 19794
rect 34242 19742 34244 19794
rect 34188 19740 34244 19742
rect 33628 18732 33684 18788
rect 34524 18786 34580 18788
rect 34524 18734 34526 18786
rect 34526 18734 34578 18786
rect 34578 18734 34580 18786
rect 34524 18732 34580 18734
rect 34076 18562 34132 18564
rect 34076 18510 34078 18562
rect 34078 18510 34130 18562
rect 34130 18510 34132 18562
rect 34076 18508 34132 18510
rect 36204 21644 36260 21700
rect 37548 22764 37604 22820
rect 37100 21644 37156 21700
rect 36428 20690 36484 20692
rect 36428 20638 36430 20690
rect 36430 20638 36482 20690
rect 36482 20638 36484 20690
rect 36428 20636 36484 20638
rect 35868 19964 35924 20020
rect 35196 19178 35252 19180
rect 35196 19126 35198 19178
rect 35198 19126 35250 19178
rect 35250 19126 35252 19178
rect 35196 19124 35252 19126
rect 35300 19178 35356 19180
rect 35300 19126 35302 19178
rect 35302 19126 35354 19178
rect 35354 19126 35356 19178
rect 35300 19124 35356 19126
rect 35404 19178 35460 19180
rect 35404 19126 35406 19178
rect 35406 19126 35458 19178
rect 35458 19126 35460 19178
rect 35404 19124 35460 19126
rect 36316 20132 36372 20188
rect 37100 20524 37156 20580
rect 36652 19964 36708 20020
rect 36092 19682 36148 19684
rect 36092 19630 36094 19682
rect 36094 19630 36146 19682
rect 36146 19630 36148 19682
rect 36092 19628 36148 19630
rect 38220 22764 38276 22820
rect 37884 21810 37940 21812
rect 37884 21758 37886 21810
rect 37886 21758 37938 21810
rect 37938 21758 37940 21810
rect 37884 21756 37940 21758
rect 37660 20524 37716 20580
rect 37100 19628 37156 19684
rect 37660 20076 37716 20132
rect 38220 21756 38276 21812
rect 38780 20860 38836 20916
rect 38556 20690 38612 20692
rect 38556 20638 38558 20690
rect 38558 20638 38610 20690
rect 38610 20638 38612 20690
rect 38556 20636 38612 20638
rect 37772 19964 37828 20020
rect 39340 23938 39396 23940
rect 39340 23886 39342 23938
rect 39342 23886 39394 23938
rect 39394 23886 39396 23938
rect 39340 23884 39396 23886
rect 38668 19964 38724 20020
rect 36204 18732 36260 18788
rect 36652 18732 36708 18788
rect 34972 18674 35028 18676
rect 34972 18622 34974 18674
rect 34974 18622 35026 18674
rect 35026 18622 35028 18674
rect 34972 18620 35028 18622
rect 34748 18508 34804 18564
rect 36316 18562 36372 18564
rect 36316 18510 36318 18562
rect 36318 18510 36370 18562
rect 36370 18510 36372 18562
rect 36316 18508 36372 18510
rect 34636 17836 34692 17892
rect 33516 17500 33572 17556
rect 33628 15372 33684 15428
rect 33740 15036 33796 15092
rect 34188 17666 34244 17668
rect 34188 17614 34190 17666
rect 34190 17614 34242 17666
rect 34242 17614 34244 17666
rect 34188 17612 34244 17614
rect 34748 17276 34804 17332
rect 35644 17500 35700 17556
rect 35196 17162 35252 17164
rect 35196 17110 35198 17162
rect 35198 17110 35250 17162
rect 35250 17110 35252 17162
rect 35196 17108 35252 17110
rect 35300 17162 35356 17164
rect 35300 17110 35302 17162
rect 35302 17110 35354 17162
rect 35354 17110 35356 17162
rect 35300 17108 35356 17110
rect 35404 17162 35460 17164
rect 35404 17110 35406 17162
rect 35406 17110 35458 17162
rect 35458 17110 35460 17162
rect 35404 17108 35460 17110
rect 34412 15596 34468 15652
rect 34188 15372 34244 15428
rect 35196 15146 35252 15148
rect 35196 15094 35198 15146
rect 35198 15094 35250 15146
rect 35250 15094 35252 15146
rect 35196 15092 35252 15094
rect 35300 15146 35356 15148
rect 35300 15094 35302 15146
rect 35302 15094 35354 15146
rect 35354 15094 35356 15146
rect 35300 15092 35356 15094
rect 35404 15146 35460 15148
rect 35404 15094 35406 15146
rect 35406 15094 35458 15146
rect 35458 15094 35460 15146
rect 35404 15092 35460 15094
rect 33740 14588 33796 14644
rect 35084 14642 35140 14644
rect 35084 14590 35086 14642
rect 35086 14590 35138 14642
rect 35138 14590 35140 14642
rect 35084 14588 35140 14590
rect 35532 14418 35588 14420
rect 35532 14366 35534 14418
rect 35534 14366 35586 14418
rect 35586 14366 35588 14418
rect 35532 14364 35588 14366
rect 35980 15820 36036 15876
rect 36316 15596 36372 15652
rect 37772 18732 37828 18788
rect 38668 18508 38724 18564
rect 40012 25900 40068 25956
rect 40124 24498 40180 24500
rect 40124 24446 40126 24498
rect 40126 24446 40178 24498
rect 40178 24446 40180 24498
rect 40124 24444 40180 24446
rect 40236 24220 40292 24276
rect 40572 26738 40628 26740
rect 40572 26686 40574 26738
rect 40574 26686 40626 26738
rect 40626 26686 40628 26738
rect 40572 26684 40628 26686
rect 42140 27970 42196 27972
rect 42140 27918 42142 27970
rect 42142 27918 42194 27970
rect 42194 27918 42196 27970
rect 42140 27916 42196 27918
rect 41020 27804 41076 27860
rect 41356 27858 41412 27860
rect 41356 27806 41358 27858
rect 41358 27806 41410 27858
rect 41410 27806 41412 27858
rect 41356 27804 41412 27806
rect 41356 27580 41412 27636
rect 42588 28642 42644 28644
rect 42588 28590 42590 28642
rect 42590 28590 42642 28642
rect 42642 28590 42644 28642
rect 42588 28588 42644 28590
rect 42028 27692 42084 27748
rect 40684 26572 40740 26628
rect 41244 26402 41300 26404
rect 41244 26350 41246 26402
rect 41246 26350 41298 26402
rect 41298 26350 41300 26402
rect 41244 26348 41300 26350
rect 40572 25116 40628 25172
rect 40348 23436 40404 23492
rect 40460 24108 40516 24164
rect 39900 21810 39956 21812
rect 39900 21758 39902 21810
rect 39902 21758 39954 21810
rect 39954 21758 39956 21810
rect 39900 21756 39956 21758
rect 40460 21756 40516 21812
rect 40796 24444 40852 24500
rect 42364 27916 42420 27972
rect 42140 26572 42196 26628
rect 42140 25954 42196 25956
rect 42140 25902 42142 25954
rect 42142 25902 42194 25954
rect 42194 25902 42196 25954
rect 42140 25900 42196 25902
rect 42028 25730 42084 25732
rect 42028 25678 42030 25730
rect 42030 25678 42082 25730
rect 42082 25678 42084 25730
rect 42028 25676 42084 25678
rect 41468 24444 41524 24500
rect 42140 24444 42196 24500
rect 41692 24220 41748 24276
rect 41244 23884 41300 23940
rect 41580 24108 41636 24164
rect 41020 22764 41076 22820
rect 41916 23884 41972 23940
rect 44380 29820 44436 29876
rect 45276 32732 45332 32788
rect 46060 34860 46116 34916
rect 47180 34860 47236 34916
rect 45724 32786 45780 32788
rect 45724 32734 45726 32786
rect 45726 32734 45778 32786
rect 45778 32734 45780 32786
rect 45724 32732 45780 32734
rect 46620 33740 46676 33796
rect 46732 33682 46788 33684
rect 46732 33630 46734 33682
rect 46734 33630 46786 33682
rect 46786 33630 46788 33682
rect 46732 33628 46788 33630
rect 46060 31778 46116 31780
rect 46060 31726 46062 31778
rect 46062 31726 46114 31778
rect 46114 31726 46116 31778
rect 46060 31724 46116 31726
rect 45500 30546 45556 30548
rect 45500 30494 45502 30546
rect 45502 30494 45554 30546
rect 45554 30494 45556 30546
rect 45500 30492 45556 30494
rect 46284 30380 46340 30436
rect 45724 29986 45780 29988
rect 45724 29934 45726 29986
rect 45726 29934 45778 29986
rect 45778 29934 45780 29986
rect 45724 29932 45780 29934
rect 45388 29874 45444 29876
rect 45388 29822 45390 29874
rect 45390 29822 45442 29874
rect 45442 29822 45444 29874
rect 45388 29820 45444 29822
rect 43260 29596 43316 29652
rect 43260 28364 43316 28420
rect 43260 27970 43316 27972
rect 43260 27918 43262 27970
rect 43262 27918 43314 27970
rect 43314 27918 43316 27970
rect 43260 27916 43316 27918
rect 44268 29484 44324 29540
rect 42812 27804 42868 27860
rect 43596 27804 43652 27860
rect 44380 29372 44436 29428
rect 44716 28476 44772 28532
rect 45052 28364 45108 28420
rect 45164 27970 45220 27972
rect 45164 27918 45166 27970
rect 45166 27918 45218 27970
rect 45218 27918 45220 27970
rect 45164 27916 45220 27918
rect 44716 26850 44772 26852
rect 44716 26798 44718 26850
rect 44718 26798 44770 26850
rect 44770 26798 44772 26850
rect 44716 26796 44772 26798
rect 44268 26684 44324 26740
rect 42924 26626 42980 26628
rect 42924 26574 42926 26626
rect 42926 26574 42978 26626
rect 42978 26574 42980 26626
rect 42924 26572 42980 26574
rect 43820 25842 43876 25844
rect 43820 25790 43822 25842
rect 43822 25790 43874 25842
rect 43874 25790 43876 25842
rect 43820 25788 43876 25790
rect 42476 25676 42532 25732
rect 45500 28530 45556 28532
rect 45500 28478 45502 28530
rect 45502 28478 45554 28530
rect 45554 28478 45556 28530
rect 45500 28476 45556 28478
rect 46060 27970 46116 27972
rect 46060 27918 46062 27970
rect 46062 27918 46114 27970
rect 46114 27918 46116 27970
rect 46060 27916 46116 27918
rect 45612 27804 45668 27860
rect 46396 29372 46452 29428
rect 46620 30380 46676 30436
rect 49084 40572 49140 40628
rect 49196 40460 49252 40516
rect 49532 40738 49588 40740
rect 49532 40686 49534 40738
rect 49534 40686 49586 40738
rect 49586 40686 49588 40738
rect 49532 40684 49588 40686
rect 50652 47794 50708 47796
rect 50652 47742 50654 47794
rect 50654 47742 50706 47794
rect 50706 47742 50708 47794
rect 50652 47740 50708 47742
rect 50556 46394 50612 46396
rect 50556 46342 50558 46394
rect 50558 46342 50610 46394
rect 50610 46342 50612 46394
rect 50556 46340 50612 46342
rect 50660 46394 50716 46396
rect 50660 46342 50662 46394
rect 50662 46342 50714 46394
rect 50714 46342 50716 46394
rect 50660 46340 50716 46342
rect 50764 46394 50820 46396
rect 50764 46342 50766 46394
rect 50766 46342 50818 46394
rect 50818 46342 50820 46394
rect 50764 46340 50820 46342
rect 50316 45388 50372 45444
rect 50204 44828 50260 44884
rect 50988 44882 51044 44884
rect 50988 44830 50990 44882
rect 50990 44830 51042 44882
rect 51042 44830 51044 44882
rect 50988 44828 51044 44830
rect 50652 44604 50708 44660
rect 50876 44716 50932 44772
rect 50556 44378 50612 44380
rect 50556 44326 50558 44378
rect 50558 44326 50610 44378
rect 50610 44326 50612 44378
rect 50556 44324 50612 44326
rect 50660 44378 50716 44380
rect 50660 44326 50662 44378
rect 50662 44326 50714 44378
rect 50714 44326 50716 44378
rect 50660 44324 50716 44326
rect 50764 44378 50820 44380
rect 50764 44326 50766 44378
rect 50766 44326 50818 44378
rect 50818 44326 50820 44378
rect 50764 44324 50820 44326
rect 50204 43708 50260 43764
rect 50876 43874 50932 43876
rect 50876 43822 50878 43874
rect 50878 43822 50930 43874
rect 50930 43822 50932 43874
rect 50876 43820 50932 43822
rect 51212 44770 51268 44772
rect 51212 44718 51214 44770
rect 51214 44718 51266 44770
rect 51266 44718 51268 44770
rect 51212 44716 51268 44718
rect 51436 44658 51492 44660
rect 51436 44606 51438 44658
rect 51438 44606 51490 44658
rect 51490 44606 51492 44658
rect 51436 44604 51492 44606
rect 50204 42866 50260 42868
rect 50204 42814 50206 42866
rect 50206 42814 50258 42866
rect 50258 42814 50260 42866
rect 50204 42812 50260 42814
rect 50092 41804 50148 41860
rect 49756 40460 49812 40516
rect 48188 39842 48244 39844
rect 48188 39790 48190 39842
rect 48190 39790 48242 39842
rect 48242 39790 48244 39842
rect 48188 39788 48244 39790
rect 47516 39618 47572 39620
rect 47516 39566 47518 39618
rect 47518 39566 47570 39618
rect 47570 39566 47572 39618
rect 47516 39564 47572 39566
rect 48188 38892 48244 38948
rect 49420 40236 49476 40292
rect 49980 40012 50036 40068
rect 48636 38780 48692 38836
rect 47628 38668 47684 38724
rect 48188 38722 48244 38724
rect 48188 38670 48190 38722
rect 48190 38670 48242 38722
rect 48242 38670 48244 38722
rect 48188 38668 48244 38670
rect 49308 39564 49364 39620
rect 53452 47794 53508 47796
rect 53452 47742 53454 47794
rect 53454 47742 53506 47794
rect 53506 47742 53508 47794
rect 53452 47740 53508 47742
rect 52556 45388 52612 45444
rect 52668 45276 52724 45332
rect 52332 45164 52388 45220
rect 51884 44770 51940 44772
rect 51884 44718 51886 44770
rect 51886 44718 51938 44770
rect 51938 44718 51940 44770
rect 51884 44716 51940 44718
rect 51884 43986 51940 43988
rect 51884 43934 51886 43986
rect 51886 43934 51938 43986
rect 51938 43934 51940 43986
rect 51884 43932 51940 43934
rect 52668 44770 52724 44772
rect 52668 44718 52670 44770
rect 52670 44718 52722 44770
rect 52722 44718 52724 44770
rect 52668 44716 52724 44718
rect 52332 43820 52388 43876
rect 52892 43874 52948 43876
rect 52892 43822 52894 43874
rect 52894 43822 52946 43874
rect 52946 43822 52948 43874
rect 52892 43820 52948 43822
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50540 42140 50596 42196
rect 50428 41634 50484 41636
rect 50428 41582 50430 41634
rect 50430 41582 50482 41634
rect 50482 41582 50484 41634
rect 50428 41580 50484 41582
rect 50204 40460 50260 40516
rect 50876 42082 50932 42084
rect 50876 42030 50878 42082
rect 50878 42030 50930 42082
rect 50930 42030 50932 42082
rect 50876 42028 50932 42030
rect 50540 40460 50596 40516
rect 50556 40346 50612 40348
rect 50556 40294 50558 40346
rect 50558 40294 50610 40346
rect 50610 40294 50612 40346
rect 50556 40292 50612 40294
rect 50660 40346 50716 40348
rect 50660 40294 50662 40346
rect 50662 40294 50714 40346
rect 50714 40294 50716 40346
rect 50660 40292 50716 40294
rect 50764 40346 50820 40348
rect 50764 40294 50766 40346
rect 50766 40294 50818 40346
rect 50818 40294 50820 40346
rect 50764 40292 50820 40294
rect 50428 38780 50484 38836
rect 50764 39788 50820 39844
rect 49084 38444 49140 38500
rect 47740 38050 47796 38052
rect 47740 37998 47742 38050
rect 47742 37998 47794 38050
rect 47794 37998 47796 38050
rect 47740 37996 47796 37998
rect 48188 37884 48244 37940
rect 49084 37938 49140 37940
rect 49084 37886 49086 37938
rect 49086 37886 49138 37938
rect 49138 37886 49140 37938
rect 49084 37884 49140 37886
rect 47852 36540 47908 36596
rect 49084 37100 49140 37156
rect 49756 38556 49812 38612
rect 49756 38050 49812 38052
rect 49756 37998 49758 38050
rect 49758 37998 49810 38050
rect 49810 37998 49812 38050
rect 49756 37996 49812 37998
rect 51212 42028 51268 42084
rect 51548 42028 51604 42084
rect 51996 42642 52052 42644
rect 51996 42590 51998 42642
rect 51998 42590 52050 42642
rect 52050 42590 52052 42642
rect 51996 42588 52052 42590
rect 51324 41746 51380 41748
rect 51324 41694 51326 41746
rect 51326 41694 51378 41746
rect 51378 41694 51380 41746
rect 51324 41692 51380 41694
rect 52220 41970 52276 41972
rect 52220 41918 52222 41970
rect 52222 41918 52274 41970
rect 52274 41918 52276 41970
rect 52220 41916 52276 41918
rect 51996 41804 52052 41860
rect 52332 41692 52388 41748
rect 53004 40850 53060 40852
rect 53004 40798 53006 40850
rect 53006 40798 53058 40850
rect 53058 40798 53060 40850
rect 53004 40796 53060 40798
rect 53788 46002 53844 46004
rect 53788 45950 53790 46002
rect 53790 45950 53842 46002
rect 53842 45950 53844 46002
rect 53788 45948 53844 45950
rect 53452 45164 53508 45220
rect 53676 44828 53732 44884
rect 53116 44604 53172 44660
rect 53340 43932 53396 43988
rect 53116 42812 53172 42868
rect 50764 38722 50820 38724
rect 50764 38670 50766 38722
rect 50766 38670 50818 38722
rect 50818 38670 50820 38722
rect 50764 38668 50820 38670
rect 51996 39788 52052 39844
rect 51996 38892 52052 38948
rect 52108 38668 52164 38724
rect 51100 38556 51156 38612
rect 50652 38444 50708 38500
rect 49420 35922 49476 35924
rect 49420 35870 49422 35922
rect 49422 35870 49474 35922
rect 49474 35870 49476 35922
rect 49420 35868 49476 35870
rect 48972 35698 49028 35700
rect 48972 35646 48974 35698
rect 48974 35646 49026 35698
rect 49026 35646 49028 35698
rect 48972 35644 49028 35646
rect 48188 34860 48244 34916
rect 49420 34914 49476 34916
rect 49420 34862 49422 34914
rect 49422 34862 49474 34914
rect 49474 34862 49476 34914
rect 49420 34860 49476 34862
rect 48860 34748 48916 34804
rect 47068 32786 47124 32788
rect 47068 32734 47070 32786
rect 47070 32734 47122 32786
rect 47122 32734 47124 32786
rect 47068 32732 47124 32734
rect 47292 32956 47348 33012
rect 49868 34802 49924 34804
rect 49868 34750 49870 34802
rect 49870 34750 49922 34802
rect 49922 34750 49924 34802
rect 49868 34748 49924 34750
rect 50204 36540 50260 36596
rect 50204 35922 50260 35924
rect 50204 35870 50206 35922
rect 50206 35870 50258 35922
rect 50258 35870 50260 35922
rect 50204 35868 50260 35870
rect 50092 35698 50148 35700
rect 50092 35646 50094 35698
rect 50094 35646 50146 35698
rect 50146 35646 50148 35698
rect 50092 35644 50148 35646
rect 49980 34636 50036 34692
rect 48860 33740 48916 33796
rect 46732 30156 46788 30212
rect 47852 31612 47908 31668
rect 49868 33404 49924 33460
rect 47964 31724 48020 31780
rect 48748 31666 48804 31668
rect 48748 31614 48750 31666
rect 48750 31614 48802 31666
rect 48802 31614 48804 31666
rect 48748 31612 48804 31614
rect 47964 30716 48020 30772
rect 48188 30492 48244 30548
rect 47068 29708 47124 29764
rect 47404 29708 47460 29764
rect 46732 29372 46788 29428
rect 46396 28866 46452 28868
rect 46396 28814 46398 28866
rect 46398 28814 46450 28866
rect 46450 28814 46452 28866
rect 46396 28812 46452 28814
rect 46508 27916 46564 27972
rect 47068 28812 47124 28868
rect 45500 26738 45556 26740
rect 45500 26686 45502 26738
rect 45502 26686 45554 26738
rect 45554 26686 45556 26738
rect 45500 26684 45556 26686
rect 45612 26626 45668 26628
rect 45612 26574 45614 26626
rect 45614 26574 45666 26626
rect 45666 26574 45668 26626
rect 45612 26572 45668 26574
rect 45612 25788 45668 25844
rect 44380 25730 44436 25732
rect 44380 25678 44382 25730
rect 44382 25678 44434 25730
rect 44434 25678 44436 25730
rect 44380 25676 44436 25678
rect 43820 25452 43876 25508
rect 42364 24108 42420 24164
rect 42476 23884 42532 23940
rect 41916 22818 41972 22820
rect 41916 22766 41918 22818
rect 41918 22766 41970 22818
rect 41970 22766 41972 22818
rect 41916 22764 41972 22766
rect 41132 21756 41188 21812
rect 40124 20860 40180 20916
rect 40012 20578 40068 20580
rect 40012 20526 40014 20578
rect 40014 20526 40066 20578
rect 40066 20526 40068 20578
rect 40012 20524 40068 20526
rect 39228 19628 39284 19684
rect 39116 18786 39172 18788
rect 39116 18734 39118 18786
rect 39118 18734 39170 18786
rect 39170 18734 39172 18786
rect 39116 18732 39172 18734
rect 39452 19740 39508 19796
rect 38780 18620 38836 18676
rect 39788 18450 39844 18452
rect 39788 18398 39790 18450
rect 39790 18398 39842 18450
rect 39842 18398 39844 18450
rect 39788 18396 39844 18398
rect 40684 20914 40740 20916
rect 40684 20862 40686 20914
rect 40686 20862 40738 20914
rect 40738 20862 40740 20914
rect 40684 20860 40740 20862
rect 41244 21644 41300 21700
rect 38780 17836 38836 17892
rect 39452 17890 39508 17892
rect 39452 17838 39454 17890
rect 39454 17838 39506 17890
rect 39506 17838 39508 17890
rect 39452 17836 39508 17838
rect 36764 17554 36820 17556
rect 36764 17502 36766 17554
rect 36766 17502 36818 17554
rect 36818 17502 36820 17554
rect 36764 17500 36820 17502
rect 39900 17890 39956 17892
rect 39900 17838 39902 17890
rect 39902 17838 39954 17890
rect 39954 17838 39956 17890
rect 39900 17836 39956 17838
rect 39788 17500 39844 17556
rect 36428 14924 36484 14980
rect 36652 14364 36708 14420
rect 36764 17276 36820 17332
rect 39228 16604 39284 16660
rect 39900 16604 39956 16660
rect 38556 16380 38612 16436
rect 37100 15874 37156 15876
rect 37100 15822 37102 15874
rect 37102 15822 37154 15874
rect 37154 15822 37156 15874
rect 37100 15820 37156 15822
rect 37548 15762 37604 15764
rect 37548 15710 37550 15762
rect 37550 15710 37602 15762
rect 37602 15710 37604 15762
rect 37548 15708 37604 15710
rect 37996 15650 38052 15652
rect 37996 15598 37998 15650
rect 37998 15598 38050 15650
rect 38050 15598 38052 15650
rect 37996 15596 38052 15598
rect 37884 14924 37940 14980
rect 37324 14754 37380 14756
rect 37324 14702 37326 14754
rect 37326 14702 37378 14754
rect 37378 14702 37380 14754
rect 37324 14700 37380 14702
rect 38668 14700 38724 14756
rect 38220 14642 38276 14644
rect 38220 14590 38222 14642
rect 38222 14590 38274 14642
rect 38274 14590 38276 14642
rect 38220 14588 38276 14590
rect 37772 14364 37828 14420
rect 35196 13130 35252 13132
rect 35196 13078 35198 13130
rect 35198 13078 35250 13130
rect 35250 13078 35252 13130
rect 35196 13076 35252 13078
rect 35300 13130 35356 13132
rect 35300 13078 35302 13130
rect 35302 13078 35354 13130
rect 35354 13078 35356 13130
rect 35300 13076 35356 13078
rect 35404 13130 35460 13132
rect 35404 13078 35406 13130
rect 35406 13078 35458 13130
rect 35458 13078 35460 13130
rect 35404 13076 35460 13078
rect 33404 12684 33460 12740
rect 33740 12738 33796 12740
rect 33740 12686 33742 12738
rect 33742 12686 33794 12738
rect 33794 12686 33796 12738
rect 33740 12684 33796 12686
rect 31164 11452 31220 11508
rect 31948 11340 32004 11396
rect 31724 10668 31780 10724
rect 31164 10108 31220 10164
rect 32508 10556 32564 10612
rect 32396 10498 32452 10500
rect 32396 10446 32398 10498
rect 32398 10446 32450 10498
rect 32450 10446 32452 10498
rect 32396 10444 32452 10446
rect 35532 12402 35588 12404
rect 35532 12350 35534 12402
rect 35534 12350 35586 12402
rect 35586 12350 35588 12402
rect 35532 12348 35588 12350
rect 33068 11506 33124 11508
rect 33068 11454 33070 11506
rect 33070 11454 33122 11506
rect 33122 11454 33124 11506
rect 33068 11452 33124 11454
rect 35196 11114 35252 11116
rect 35196 11062 35198 11114
rect 35198 11062 35250 11114
rect 35250 11062 35252 11114
rect 35196 11060 35252 11062
rect 35300 11114 35356 11116
rect 35300 11062 35302 11114
rect 35302 11062 35354 11114
rect 35354 11062 35356 11114
rect 35300 11060 35356 11062
rect 35404 11114 35460 11116
rect 35404 11062 35406 11114
rect 35406 11062 35458 11114
rect 35458 11062 35460 11114
rect 35404 11060 35460 11062
rect 35980 12402 36036 12404
rect 35980 12350 35982 12402
rect 35982 12350 36034 12402
rect 36034 12350 36036 12402
rect 35980 12348 36036 12350
rect 35868 11340 35924 11396
rect 35980 10722 36036 10724
rect 35980 10670 35982 10722
rect 35982 10670 36034 10722
rect 36034 10670 36036 10722
rect 35980 10668 36036 10670
rect 37324 12402 37380 12404
rect 37324 12350 37326 12402
rect 37326 12350 37378 12402
rect 37378 12350 37380 12402
rect 37324 12348 37380 12350
rect 34188 10610 34244 10612
rect 34188 10558 34190 10610
rect 34190 10558 34242 10610
rect 34242 10558 34244 10610
rect 34188 10556 34244 10558
rect 36540 10556 36596 10612
rect 33628 10444 33684 10500
rect 33964 9996 34020 10052
rect 35196 9996 35252 10052
rect 36428 9996 36484 10052
rect 35196 9098 35252 9100
rect 35196 9046 35198 9098
rect 35198 9046 35250 9098
rect 35250 9046 35252 9098
rect 35196 9044 35252 9046
rect 35300 9098 35356 9100
rect 35300 9046 35302 9098
rect 35302 9046 35354 9098
rect 35354 9046 35356 9098
rect 35300 9044 35356 9046
rect 35404 9098 35460 9100
rect 35404 9046 35406 9098
rect 35406 9046 35458 9098
rect 35458 9046 35460 9098
rect 35404 9044 35460 9046
rect 37324 10780 37380 10836
rect 37324 10108 37380 10164
rect 39004 13580 39060 13636
rect 37660 12348 37716 12404
rect 38220 12402 38276 12404
rect 38220 12350 38222 12402
rect 38222 12350 38274 12402
rect 38274 12350 38276 12402
rect 38220 12348 38276 12350
rect 37772 11676 37828 11732
rect 37772 10668 37828 10724
rect 38556 11676 38612 11732
rect 39452 13580 39508 13636
rect 40124 18562 40180 18564
rect 40124 18510 40126 18562
rect 40126 18510 40178 18562
rect 40178 18510 40180 18562
rect 40124 18508 40180 18510
rect 40348 17554 40404 17556
rect 40348 17502 40350 17554
rect 40350 17502 40402 17554
rect 40402 17502 40404 17554
rect 40348 17500 40404 17502
rect 41020 19682 41076 19684
rect 41020 19630 41022 19682
rect 41022 19630 41074 19682
rect 41074 19630 41076 19682
rect 41020 19628 41076 19630
rect 41468 21474 41524 21476
rect 41468 21422 41470 21474
rect 41470 21422 41522 21474
rect 41522 21422 41524 21474
rect 41468 21420 41524 21422
rect 41580 21308 41636 21364
rect 43036 22818 43092 22820
rect 43036 22766 43038 22818
rect 43038 22766 43090 22818
rect 43090 22766 43092 22818
rect 43036 22764 43092 22766
rect 43484 22818 43540 22820
rect 43484 22766 43486 22818
rect 43486 22766 43538 22818
rect 43538 22766 43540 22818
rect 43484 22764 43540 22766
rect 41692 21532 41748 21588
rect 43036 21698 43092 21700
rect 43036 21646 43038 21698
rect 43038 21646 43090 21698
rect 43090 21646 43092 21698
rect 43036 21644 43092 21646
rect 42252 21586 42308 21588
rect 42252 21534 42254 21586
rect 42254 21534 42306 21586
rect 42306 21534 42308 21586
rect 42252 21532 42308 21534
rect 42700 21308 42756 21364
rect 41804 20972 41860 21028
rect 43036 21026 43092 21028
rect 43036 20974 43038 21026
rect 43038 20974 43090 21026
rect 43090 20974 43092 21026
rect 43036 20972 43092 20974
rect 43372 20860 43428 20916
rect 41580 20578 41636 20580
rect 41580 20526 41582 20578
rect 41582 20526 41634 20578
rect 41634 20526 41636 20578
rect 41580 20524 41636 20526
rect 41356 19628 41412 19684
rect 41020 18508 41076 18564
rect 42812 20466 42868 20468
rect 42812 20414 42814 20466
rect 42814 20414 42866 20466
rect 42866 20414 42868 20466
rect 42812 20412 42868 20414
rect 41244 18508 41300 18564
rect 41132 18396 41188 18452
rect 40908 17500 40964 17556
rect 41468 17890 41524 17892
rect 41468 17838 41470 17890
rect 41470 17838 41522 17890
rect 41522 17838 41524 17890
rect 41468 17836 41524 17838
rect 41244 17724 41300 17780
rect 40236 15874 40292 15876
rect 40236 15822 40238 15874
rect 40238 15822 40290 15874
rect 40290 15822 40292 15874
rect 40236 15820 40292 15822
rect 40012 13692 40068 13748
rect 38892 12348 38948 12404
rect 38668 10780 38724 10836
rect 38444 10556 38500 10612
rect 41132 16546 41188 16548
rect 41132 16494 41134 16546
rect 41134 16494 41186 16546
rect 41186 16494 41188 16546
rect 41132 16492 41188 16494
rect 40684 16434 40740 16436
rect 40684 16382 40686 16434
rect 40686 16382 40738 16434
rect 40738 16382 40740 16434
rect 40684 16380 40740 16382
rect 41244 15874 41300 15876
rect 41244 15822 41246 15874
rect 41246 15822 41298 15874
rect 41298 15822 41300 15874
rect 41244 15820 41300 15822
rect 41804 19628 41860 19684
rect 44268 23996 44324 24052
rect 44380 23938 44436 23940
rect 44380 23886 44382 23938
rect 44382 23886 44434 23938
rect 44434 23886 44436 23938
rect 44380 23884 44436 23886
rect 45276 24834 45332 24836
rect 45276 24782 45278 24834
rect 45278 24782 45330 24834
rect 45330 24782 45332 24834
rect 45276 24780 45332 24782
rect 46956 27804 47012 27860
rect 46060 25730 46116 25732
rect 46060 25678 46062 25730
rect 46062 25678 46114 25730
rect 46114 25678 46116 25730
rect 46060 25676 46116 25678
rect 45724 24834 45780 24836
rect 45724 24782 45726 24834
rect 45726 24782 45778 24834
rect 45778 24782 45780 24834
rect 45724 24780 45780 24782
rect 46396 24780 46452 24836
rect 45612 23884 45668 23940
rect 46060 23996 46116 24052
rect 45724 23772 45780 23828
rect 44940 22482 44996 22484
rect 44940 22430 44942 22482
rect 44942 22430 44994 22482
rect 44994 22430 44996 22482
rect 44940 22428 44996 22430
rect 43708 20412 43764 20468
rect 43484 18508 43540 18564
rect 42252 17948 42308 18004
rect 42140 17836 42196 17892
rect 41692 17612 41748 17668
rect 41916 17500 41972 17556
rect 43260 17836 43316 17892
rect 42252 17778 42308 17780
rect 42252 17726 42254 17778
rect 42254 17726 42306 17778
rect 42306 17726 42308 17778
rect 42252 17724 42308 17726
rect 44492 17836 44548 17892
rect 43708 17724 43764 17780
rect 42700 17666 42756 17668
rect 42700 17614 42702 17666
rect 42702 17614 42754 17666
rect 42754 17614 42756 17666
rect 42700 17612 42756 17614
rect 41692 14476 41748 14532
rect 41132 13580 41188 13636
rect 43484 14588 43540 14644
rect 43484 13580 43540 13636
rect 39228 10780 39284 10836
rect 41020 10780 41076 10836
rect 41580 10780 41636 10836
rect 42364 10780 42420 10836
rect 42028 10722 42084 10724
rect 42028 10670 42030 10722
rect 42030 10670 42082 10722
rect 42082 10670 42084 10722
rect 42028 10668 42084 10670
rect 45052 20690 45108 20692
rect 45052 20638 45054 20690
rect 45054 20638 45106 20690
rect 45106 20638 45108 20690
rect 45052 20636 45108 20638
rect 46508 21644 46564 21700
rect 48076 28812 48132 28868
rect 47740 28588 47796 28644
rect 49308 32450 49364 32452
rect 49308 32398 49310 32450
rect 49310 32398 49362 32450
rect 49362 32398 49364 32450
rect 49308 32396 49364 32398
rect 50204 32562 50260 32564
rect 50204 32510 50206 32562
rect 50206 32510 50258 32562
rect 50258 32510 50260 32562
rect 50204 32508 50260 32510
rect 50092 31778 50148 31780
rect 50092 31726 50094 31778
rect 50094 31726 50146 31778
rect 50146 31726 50148 31778
rect 50092 31724 50148 31726
rect 49084 30940 49140 30996
rect 48972 30604 49028 30660
rect 51772 38444 51828 38500
rect 50556 38330 50612 38332
rect 50556 38278 50558 38330
rect 50558 38278 50610 38330
rect 50610 38278 50612 38330
rect 50556 38276 50612 38278
rect 50660 38330 50716 38332
rect 50660 38278 50662 38330
rect 50662 38278 50714 38330
rect 50714 38278 50716 38330
rect 50660 38276 50716 38278
rect 50764 38330 50820 38332
rect 50764 38278 50766 38330
rect 50766 38278 50818 38330
rect 50818 38278 50820 38330
rect 50764 38276 50820 38278
rect 51548 37826 51604 37828
rect 51548 37774 51550 37826
rect 51550 37774 51602 37826
rect 51602 37774 51604 37826
rect 51548 37772 51604 37774
rect 52780 38946 52836 38948
rect 52780 38894 52782 38946
rect 52782 38894 52834 38946
rect 52834 38894 52836 38946
rect 52780 38892 52836 38894
rect 53452 42588 53508 42644
rect 54908 46002 54964 46004
rect 54908 45950 54910 46002
rect 54910 45950 54962 46002
rect 54962 45950 54964 46002
rect 54908 45948 54964 45950
rect 54124 45388 54180 45444
rect 54796 44882 54852 44884
rect 54796 44830 54798 44882
rect 54798 44830 54850 44882
rect 54850 44830 54852 44882
rect 54796 44828 54852 44830
rect 54012 43932 54068 43988
rect 54684 43986 54740 43988
rect 54684 43934 54686 43986
rect 54686 43934 54738 43986
rect 54738 43934 54740 43986
rect 54684 43932 54740 43934
rect 55356 46002 55412 46004
rect 55356 45950 55358 46002
rect 55358 45950 55410 46002
rect 55410 45950 55412 46002
rect 55356 45948 55412 45950
rect 56700 43986 56756 43988
rect 56700 43934 56702 43986
rect 56702 43934 56754 43986
rect 56754 43934 56756 43986
rect 56700 43932 56756 43934
rect 57148 43986 57204 43988
rect 57148 43934 57150 43986
rect 57150 43934 57202 43986
rect 57202 43934 57204 43986
rect 57148 43932 57204 43934
rect 53676 42140 53732 42196
rect 53564 41916 53620 41972
rect 54460 42812 54516 42868
rect 54236 42754 54292 42756
rect 54236 42702 54238 42754
rect 54238 42702 54290 42754
rect 54290 42702 54292 42754
rect 54236 42700 54292 42702
rect 56140 42924 56196 42980
rect 55132 42812 55188 42868
rect 55020 42700 55076 42756
rect 54348 42028 54404 42084
rect 53788 41580 53844 41636
rect 53676 40626 53732 40628
rect 53676 40574 53678 40626
rect 53678 40574 53730 40626
rect 53730 40574 53732 40626
rect 53676 40572 53732 40574
rect 50876 36652 50932 36708
rect 51212 36540 51268 36596
rect 50556 36314 50612 36316
rect 50556 36262 50558 36314
rect 50558 36262 50610 36314
rect 50610 36262 50612 36314
rect 50556 36260 50612 36262
rect 50660 36314 50716 36316
rect 50660 36262 50662 36314
rect 50662 36262 50714 36314
rect 50714 36262 50716 36314
rect 50660 36260 50716 36262
rect 50764 36314 50820 36316
rect 50764 36262 50766 36314
rect 50766 36262 50818 36314
rect 50818 36262 50820 36314
rect 50764 36260 50820 36262
rect 50652 34748 50708 34804
rect 50556 34298 50612 34300
rect 50556 34246 50558 34298
rect 50558 34246 50610 34298
rect 50610 34246 50612 34298
rect 50556 34244 50612 34246
rect 50660 34298 50716 34300
rect 50660 34246 50662 34298
rect 50662 34246 50714 34298
rect 50714 34246 50716 34298
rect 50660 34244 50716 34246
rect 50764 34298 50820 34300
rect 50764 34246 50766 34298
rect 50766 34246 50818 34298
rect 50818 34246 50820 34298
rect 50764 34244 50820 34246
rect 51212 34914 51268 34916
rect 51212 34862 51214 34914
rect 51214 34862 51266 34914
rect 51266 34862 51268 34914
rect 51212 34860 51268 34862
rect 51324 34748 51380 34804
rect 51436 35644 51492 35700
rect 51884 35196 51940 35252
rect 51548 34690 51604 34692
rect 51548 34638 51550 34690
rect 51550 34638 51602 34690
rect 51602 34638 51604 34690
rect 51548 34636 51604 34638
rect 51548 34018 51604 34020
rect 51548 33966 51550 34018
rect 51550 33966 51602 34018
rect 51602 33966 51604 34018
rect 51548 33964 51604 33966
rect 50988 32620 51044 32676
rect 50556 32282 50612 32284
rect 50556 32230 50558 32282
rect 50558 32230 50610 32282
rect 50610 32230 50612 32282
rect 50556 32228 50612 32230
rect 50660 32282 50716 32284
rect 50660 32230 50662 32282
rect 50662 32230 50714 32282
rect 50714 32230 50716 32282
rect 50660 32228 50716 32230
rect 50764 32282 50820 32284
rect 50764 32230 50766 32282
rect 50766 32230 50818 32282
rect 50818 32230 50820 32282
rect 50764 32228 50820 32230
rect 50988 32396 51044 32452
rect 50316 31500 50372 31556
rect 51100 32508 51156 32564
rect 49420 30268 49476 30324
rect 48748 30156 48804 30212
rect 48300 28754 48356 28756
rect 48300 28702 48302 28754
rect 48302 28702 48354 28754
rect 48354 28702 48356 28754
rect 48300 28700 48356 28702
rect 50652 30434 50708 30436
rect 50652 30382 50654 30434
rect 50654 30382 50706 30434
rect 50706 30382 50708 30434
rect 50652 30380 50708 30382
rect 50556 30266 50612 30268
rect 50316 30156 50372 30212
rect 50556 30214 50558 30266
rect 50558 30214 50610 30266
rect 50610 30214 50612 30266
rect 50556 30212 50612 30214
rect 50660 30266 50716 30268
rect 50660 30214 50662 30266
rect 50662 30214 50714 30266
rect 50714 30214 50716 30266
rect 50660 30212 50716 30214
rect 50764 30266 50820 30268
rect 50764 30214 50766 30266
rect 50766 30214 50818 30266
rect 50818 30214 50820 30266
rect 50764 30212 50820 30214
rect 49756 28700 49812 28756
rect 50204 28812 50260 28868
rect 48972 28588 49028 28644
rect 48188 26796 48244 26852
rect 48524 27468 48580 27524
rect 47852 26460 47908 26516
rect 47628 25788 47684 25844
rect 48076 25676 48132 25732
rect 47740 21698 47796 21700
rect 47740 21646 47742 21698
rect 47742 21646 47794 21698
rect 47794 21646 47796 21698
rect 47740 21644 47796 21646
rect 48412 21644 48468 21700
rect 47404 21308 47460 21364
rect 46172 20636 46228 20692
rect 46732 20802 46788 20804
rect 46732 20750 46734 20802
rect 46734 20750 46786 20802
rect 46786 20750 46788 20802
rect 46732 20748 46788 20750
rect 47628 20802 47684 20804
rect 47628 20750 47630 20802
rect 47630 20750 47682 20802
rect 47682 20750 47684 20802
rect 47628 20748 47684 20750
rect 48076 20636 48132 20692
rect 48188 21308 48244 21364
rect 48412 20748 48468 20804
rect 49308 28476 49364 28532
rect 48636 26460 48692 26516
rect 49756 26738 49812 26740
rect 49756 26686 49758 26738
rect 49758 26686 49810 26738
rect 49810 26686 49812 26738
rect 49756 26684 49812 26686
rect 50540 28866 50596 28868
rect 50540 28814 50542 28866
rect 50542 28814 50594 28866
rect 50594 28814 50596 28866
rect 50540 28812 50596 28814
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 49644 25842 49700 25844
rect 49644 25790 49646 25842
rect 49646 25790 49698 25842
rect 49698 25790 49700 25842
rect 49644 25788 49700 25790
rect 49084 25730 49140 25732
rect 49084 25678 49086 25730
rect 49086 25678 49138 25730
rect 49138 25678 49140 25730
rect 49084 25676 49140 25678
rect 50204 25676 50260 25732
rect 48860 23826 48916 23828
rect 48860 23774 48862 23826
rect 48862 23774 48914 23826
rect 48914 23774 48916 23826
rect 48860 23772 48916 23774
rect 49420 23772 49476 23828
rect 49532 23714 49588 23716
rect 49532 23662 49534 23714
rect 49534 23662 49586 23714
rect 49586 23662 49588 23714
rect 49532 23660 49588 23662
rect 49980 23996 50036 24052
rect 50652 27970 50708 27972
rect 50652 27918 50654 27970
rect 50654 27918 50706 27970
rect 50706 27918 50708 27970
rect 50652 27916 50708 27918
rect 51436 31724 51492 31780
rect 51884 35026 51940 35028
rect 51884 34974 51886 35026
rect 51886 34974 51938 35026
rect 51938 34974 51940 35026
rect 51884 34972 51940 34974
rect 52892 37826 52948 37828
rect 52892 37774 52894 37826
rect 52894 37774 52946 37826
rect 52946 37774 52948 37826
rect 52892 37772 52948 37774
rect 52780 36706 52836 36708
rect 52780 36654 52782 36706
rect 52782 36654 52834 36706
rect 52834 36654 52836 36706
rect 52780 36652 52836 36654
rect 53116 36930 53172 36932
rect 53116 36878 53118 36930
rect 53118 36878 53170 36930
rect 53170 36878 53172 36930
rect 53116 36876 53172 36878
rect 54796 41580 54852 41636
rect 56028 42812 56084 42868
rect 55356 42700 55412 42756
rect 55692 42754 55748 42756
rect 55692 42702 55694 42754
rect 55694 42702 55746 42754
rect 55746 42702 55748 42754
rect 55692 42700 55748 42702
rect 55804 42476 55860 42532
rect 53900 40066 53956 40068
rect 53900 40014 53902 40066
rect 53902 40014 53954 40066
rect 53954 40014 53956 40066
rect 53900 40012 53956 40014
rect 56476 42866 56532 42868
rect 56476 42814 56478 42866
rect 56478 42814 56530 42866
rect 56530 42814 56532 42866
rect 56476 42812 56532 42814
rect 56924 42754 56980 42756
rect 56924 42702 56926 42754
rect 56926 42702 56978 42754
rect 56978 42702 56980 42754
rect 56924 42700 56980 42702
rect 56140 42588 56196 42644
rect 57372 42642 57428 42644
rect 57372 42590 57374 42642
rect 57374 42590 57426 42642
rect 57426 42590 57428 42642
rect 57372 42588 57428 42590
rect 56700 42530 56756 42532
rect 56700 42478 56702 42530
rect 56702 42478 56754 42530
rect 56754 42478 56756 42530
rect 56700 42476 56756 42478
rect 55804 41580 55860 41636
rect 56140 41692 56196 41748
rect 53788 38722 53844 38724
rect 53788 38670 53790 38722
rect 53790 38670 53842 38722
rect 53842 38670 53844 38722
rect 53788 38668 53844 38670
rect 55580 38892 55636 38948
rect 54684 38722 54740 38724
rect 54684 38670 54686 38722
rect 54686 38670 54738 38722
rect 54738 38670 54740 38722
rect 54684 38668 54740 38670
rect 57148 41746 57204 41748
rect 57148 41694 57150 41746
rect 57150 41694 57202 41746
rect 57202 41694 57204 41746
rect 57148 41692 57204 41694
rect 56476 38946 56532 38948
rect 56476 38894 56478 38946
rect 56478 38894 56530 38946
rect 56530 38894 56532 38946
rect 56476 38892 56532 38894
rect 56028 38722 56084 38724
rect 56028 38670 56030 38722
rect 56030 38670 56082 38722
rect 56082 38670 56084 38722
rect 56028 38668 56084 38670
rect 54348 37100 54404 37156
rect 53788 36876 53844 36932
rect 54124 36652 54180 36708
rect 53004 35196 53060 35252
rect 53116 35756 53172 35812
rect 52556 34972 52612 35028
rect 52780 34860 52836 34916
rect 52108 34748 52164 34804
rect 51884 33740 51940 33796
rect 51548 31836 51604 31892
rect 51324 31500 51380 31556
rect 51212 29650 51268 29652
rect 51212 29598 51214 29650
rect 51214 29598 51266 29650
rect 51266 29598 51268 29650
rect 51212 29596 51268 29598
rect 51548 30940 51604 30996
rect 52332 34636 52388 34692
rect 52220 33458 52276 33460
rect 52220 33406 52222 33458
rect 52222 33406 52274 33458
rect 52274 33406 52276 33458
rect 52220 33404 52276 33406
rect 51884 31836 51940 31892
rect 51660 30492 51716 30548
rect 51772 30044 51828 30100
rect 51548 28812 51604 28868
rect 52780 33852 52836 33908
rect 52668 32844 52724 32900
rect 53004 34860 53060 34916
rect 52892 33794 52948 33796
rect 52892 33742 52894 33794
rect 52894 33742 52946 33794
rect 52946 33742 52948 33794
rect 52892 33740 52948 33742
rect 53340 34972 53396 35028
rect 54348 36876 54404 36932
rect 53900 35810 53956 35812
rect 53900 35758 53902 35810
rect 53902 35758 53954 35810
rect 53954 35758 53956 35810
rect 53900 35756 53956 35758
rect 53788 34860 53844 34916
rect 55804 36652 55860 36708
rect 55916 35980 55972 36036
rect 54012 33964 54068 34020
rect 53900 33682 53956 33684
rect 53900 33630 53902 33682
rect 53902 33630 53954 33682
rect 53954 33630 53956 33682
rect 53900 33628 53956 33630
rect 53788 32844 53844 32900
rect 52444 31500 52500 31556
rect 52220 30940 52276 30996
rect 51996 29596 52052 29652
rect 52332 29650 52388 29652
rect 52332 29598 52334 29650
rect 52334 29598 52386 29650
rect 52386 29598 52388 29650
rect 52332 29596 52388 29598
rect 51884 28812 51940 28868
rect 52780 28866 52836 28868
rect 52780 28814 52782 28866
rect 52782 28814 52834 28866
rect 52834 28814 52836 28866
rect 52780 28812 52836 28814
rect 51100 27858 51156 27860
rect 51100 27806 51102 27858
rect 51102 27806 51154 27858
rect 51154 27806 51156 27858
rect 51100 27804 51156 27806
rect 51660 27916 51716 27972
rect 51884 28476 51940 28532
rect 52108 27916 52164 27972
rect 52332 27858 52388 27860
rect 52332 27806 52334 27858
rect 52334 27806 52386 27858
rect 52386 27806 52388 27858
rect 52332 27804 52388 27806
rect 50428 26684 50484 26740
rect 50988 26684 51044 26740
rect 50876 26626 50932 26628
rect 50876 26574 50878 26626
rect 50878 26574 50930 26626
rect 50930 26574 50932 26626
rect 50876 26572 50932 26574
rect 50556 26234 50612 26236
rect 50556 26182 50558 26234
rect 50558 26182 50610 26234
rect 50610 26182 50612 26234
rect 50556 26180 50612 26182
rect 50660 26234 50716 26236
rect 50660 26182 50662 26234
rect 50662 26182 50714 26234
rect 50714 26182 50716 26234
rect 50660 26180 50716 26182
rect 50764 26234 50820 26236
rect 50764 26182 50766 26234
rect 50766 26182 50818 26234
rect 50818 26182 50820 26234
rect 50764 26180 50820 26182
rect 51548 26796 51604 26852
rect 51324 26738 51380 26740
rect 51324 26686 51326 26738
rect 51326 26686 51378 26738
rect 51378 26686 51380 26738
rect 51324 26684 51380 26686
rect 51212 26572 51268 26628
rect 51660 25116 51716 25172
rect 50204 23660 50260 23716
rect 50556 24218 50612 24220
rect 50556 24166 50558 24218
rect 50558 24166 50610 24218
rect 50610 24166 50612 24218
rect 50556 24164 50612 24166
rect 50660 24218 50716 24220
rect 50660 24166 50662 24218
rect 50662 24166 50714 24218
rect 50714 24166 50716 24218
rect 50660 24164 50716 24166
rect 50764 24218 50820 24220
rect 50764 24166 50766 24218
rect 50766 24166 50818 24218
rect 50818 24166 50820 24218
rect 50764 24164 50820 24166
rect 50428 23996 50484 24052
rect 50652 23660 50708 23716
rect 49756 21756 49812 21812
rect 50556 22202 50612 22204
rect 50556 22150 50558 22202
rect 50558 22150 50610 22202
rect 50610 22150 50612 22202
rect 50556 22148 50612 22150
rect 50660 22202 50716 22204
rect 50660 22150 50662 22202
rect 50662 22150 50714 22202
rect 50714 22150 50716 22202
rect 50660 22148 50716 22150
rect 50764 22202 50820 22204
rect 50764 22150 50766 22202
rect 50766 22150 50818 22202
rect 50818 22150 50820 22202
rect 50764 22148 50820 22150
rect 50204 21644 50260 21700
rect 50764 21810 50820 21812
rect 50764 21758 50766 21810
rect 50766 21758 50818 21810
rect 50818 21758 50820 21810
rect 50764 21756 50820 21758
rect 50652 21532 50708 21588
rect 52108 26572 52164 26628
rect 52220 25730 52276 25732
rect 52220 25678 52222 25730
rect 52222 25678 52274 25730
rect 52274 25678 52276 25730
rect 52220 25676 52276 25678
rect 51884 24668 51940 24724
rect 51884 24498 51940 24500
rect 51884 24446 51886 24498
rect 51886 24446 51938 24498
rect 51938 24446 51940 24498
rect 51884 24444 51940 24446
rect 51772 23772 51828 23828
rect 51436 21756 51492 21812
rect 49308 20636 49364 20692
rect 48524 19852 48580 19908
rect 48300 19740 48356 19796
rect 47964 19628 48020 19684
rect 46172 18508 46228 18564
rect 45612 17500 45668 17556
rect 45052 16658 45108 16660
rect 45052 16606 45054 16658
rect 45054 16606 45106 16658
rect 45106 16606 45108 16658
rect 45052 16604 45108 16606
rect 45724 16604 45780 16660
rect 44604 16492 44660 16548
rect 45164 15036 45220 15092
rect 43820 14642 43876 14644
rect 43820 14590 43822 14642
rect 43822 14590 43874 14642
rect 43874 14590 43876 14642
rect 43820 14588 43876 14590
rect 44940 14642 44996 14644
rect 44940 14590 44942 14642
rect 44942 14590 44994 14642
rect 44994 14590 44996 14642
rect 44940 14588 44996 14590
rect 44268 14530 44324 14532
rect 44268 14478 44270 14530
rect 44270 14478 44322 14530
rect 44322 14478 44324 14530
rect 44268 14476 44324 14478
rect 45500 14530 45556 14532
rect 45500 14478 45502 14530
rect 45502 14478 45554 14530
rect 45554 14478 45556 14530
rect 45500 14476 45556 14478
rect 45388 13746 45444 13748
rect 45388 13694 45390 13746
rect 45390 13694 45442 13746
rect 45442 13694 45444 13746
rect 45388 13692 45444 13694
rect 45388 12348 45444 12404
rect 43484 10668 43540 10724
rect 43596 10780 43652 10836
rect 39116 10610 39172 10612
rect 39116 10558 39118 10610
rect 39118 10558 39170 10610
rect 39170 10558 39172 10610
rect 39116 10556 39172 10558
rect 41132 10610 41188 10612
rect 41132 10558 41134 10610
rect 41134 10558 41186 10610
rect 41186 10558 41188 10610
rect 41132 10556 41188 10558
rect 44044 10610 44100 10612
rect 44044 10558 44046 10610
rect 44046 10558 44098 10610
rect 44098 10558 44100 10610
rect 44044 10556 44100 10558
rect 44380 10556 44436 10612
rect 44492 10668 44548 10724
rect 45164 10610 45220 10612
rect 45164 10558 45166 10610
rect 45166 10558 45218 10610
rect 45218 10558 45220 10610
rect 45164 10556 45220 10558
rect 47180 17500 47236 17556
rect 46956 16546 47012 16548
rect 46956 16494 46958 16546
rect 46958 16494 47010 16546
rect 47010 16494 47012 16546
rect 46956 16492 47012 16494
rect 48748 19682 48804 19684
rect 48748 19630 48750 19682
rect 48750 19630 48802 19682
rect 48802 19630 48804 19682
rect 48748 19628 48804 19630
rect 47404 16604 47460 16660
rect 47292 16492 47348 16548
rect 47628 16380 47684 16436
rect 47516 15708 47572 15764
rect 48972 17500 49028 17556
rect 49756 19906 49812 19908
rect 49756 19854 49758 19906
rect 49758 19854 49810 19906
rect 49810 19854 49812 19906
rect 49756 19852 49812 19854
rect 48524 16492 48580 16548
rect 48412 16434 48468 16436
rect 48412 16382 48414 16434
rect 48414 16382 48466 16434
rect 48466 16382 48468 16434
rect 48412 16380 48468 16382
rect 50092 20636 50148 20692
rect 50764 20636 50820 20692
rect 50556 20186 50612 20188
rect 50556 20134 50558 20186
rect 50558 20134 50610 20186
rect 50610 20134 50612 20186
rect 50556 20132 50612 20134
rect 50660 20186 50716 20188
rect 50660 20134 50662 20186
rect 50662 20134 50714 20186
rect 50714 20134 50716 20186
rect 50660 20132 50716 20134
rect 50764 20186 50820 20188
rect 50764 20134 50766 20186
rect 50766 20134 50818 20186
rect 50818 20134 50820 20186
rect 50764 20132 50820 20134
rect 50204 19794 50260 19796
rect 50204 19742 50206 19794
rect 50206 19742 50258 19794
rect 50258 19742 50260 19794
rect 50204 19740 50260 19742
rect 50540 18562 50596 18564
rect 50540 18510 50542 18562
rect 50542 18510 50594 18562
rect 50594 18510 50596 18562
rect 50540 18508 50596 18510
rect 50556 18170 50612 18172
rect 50556 18118 50558 18170
rect 50558 18118 50610 18170
rect 50610 18118 50612 18170
rect 50556 18116 50612 18118
rect 50660 18170 50716 18172
rect 50660 18118 50662 18170
rect 50662 18118 50714 18170
rect 50714 18118 50716 18170
rect 50660 18116 50716 18118
rect 50764 18170 50820 18172
rect 50764 18118 50766 18170
rect 50766 18118 50818 18170
rect 50818 18118 50820 18170
rect 50764 18116 50820 18118
rect 50876 17612 50932 17668
rect 49532 17500 49588 17556
rect 48860 16434 48916 16436
rect 48860 16382 48862 16434
rect 48862 16382 48914 16434
rect 48914 16382 48916 16434
rect 48860 16380 48916 16382
rect 49196 16380 49252 16436
rect 48300 15820 48356 15876
rect 49084 15932 49140 15988
rect 48412 15596 48468 15652
rect 48636 15708 48692 15764
rect 47740 15538 47796 15540
rect 47740 15486 47742 15538
rect 47742 15486 47794 15538
rect 47794 15486 47796 15538
rect 47740 15484 47796 15486
rect 47628 15148 47684 15204
rect 49196 15874 49252 15876
rect 49196 15822 49198 15874
rect 49198 15822 49250 15874
rect 49250 15822 49252 15874
rect 49196 15820 49252 15822
rect 48972 15484 49028 15540
rect 49420 16268 49476 16324
rect 51548 17836 51604 17892
rect 53116 30044 53172 30100
rect 53900 32508 53956 32564
rect 54684 34914 54740 34916
rect 54684 34862 54686 34914
rect 54686 34862 54738 34914
rect 54738 34862 54740 34914
rect 54684 34860 54740 34862
rect 54908 34802 54964 34804
rect 54908 34750 54910 34802
rect 54910 34750 54962 34802
rect 54962 34750 54964 34802
rect 54908 34748 54964 34750
rect 55692 34690 55748 34692
rect 55692 34638 55694 34690
rect 55694 34638 55746 34690
rect 55746 34638 55748 34690
rect 55692 34636 55748 34638
rect 55020 34076 55076 34132
rect 55692 34076 55748 34132
rect 54348 33906 54404 33908
rect 54348 33854 54350 33906
rect 54350 33854 54402 33906
rect 54402 33854 54404 33906
rect 54348 33852 54404 33854
rect 55804 33682 55860 33684
rect 55804 33630 55806 33682
rect 55806 33630 55858 33682
rect 55858 33630 55860 33682
rect 55804 33628 55860 33630
rect 53900 31778 53956 31780
rect 53900 31726 53902 31778
rect 53902 31726 53954 31778
rect 53954 31726 53956 31778
rect 53900 31724 53956 31726
rect 55020 32674 55076 32676
rect 55020 32622 55022 32674
rect 55022 32622 55074 32674
rect 55074 32622 55076 32674
rect 55020 32620 55076 32622
rect 54124 32508 54180 32564
rect 54124 31948 54180 32004
rect 54124 31500 54180 31556
rect 53900 30268 53956 30324
rect 54236 30380 54292 30436
rect 54012 29596 54068 29652
rect 53228 28476 53284 28532
rect 53340 28812 53396 28868
rect 53116 27970 53172 27972
rect 53116 27918 53118 27970
rect 53118 27918 53170 27970
rect 53170 27918 53172 27970
rect 53116 27916 53172 27918
rect 51660 19740 51716 19796
rect 51996 21756 52052 21812
rect 52892 25116 52948 25172
rect 52892 24444 52948 24500
rect 54124 28866 54180 28868
rect 54124 28814 54126 28866
rect 54126 28814 54178 28866
rect 54178 28814 54180 28866
rect 54124 28812 54180 28814
rect 53676 26738 53732 26740
rect 53676 26686 53678 26738
rect 53678 26686 53730 26738
rect 53730 26686 53732 26738
rect 53676 26684 53732 26686
rect 54460 30658 54516 30660
rect 54460 30606 54462 30658
rect 54462 30606 54514 30658
rect 54514 30606 54516 30658
rect 54460 30604 54516 30606
rect 54348 28476 54404 28532
rect 55468 31724 55524 31780
rect 55468 30604 55524 30660
rect 57148 36652 57204 36708
rect 56700 36034 56756 36036
rect 56700 35982 56702 36034
rect 56702 35982 56754 36034
rect 56754 35982 56756 36034
rect 56700 35980 56756 35982
rect 56140 34914 56196 34916
rect 56140 34862 56142 34914
rect 56142 34862 56194 34914
rect 56194 34862 56196 34914
rect 56140 34860 56196 34862
rect 56588 34690 56644 34692
rect 56588 34638 56590 34690
rect 56590 34638 56642 34690
rect 56642 34638 56644 34690
rect 56588 34636 56644 34638
rect 56028 31836 56084 31892
rect 55692 31612 55748 31668
rect 56700 31836 56756 31892
rect 56476 31778 56532 31780
rect 56476 31726 56478 31778
rect 56478 31726 56530 31778
rect 56530 31726 56532 31778
rect 56476 31724 56532 31726
rect 57036 31724 57092 31780
rect 57148 32002 57204 32004
rect 57148 31950 57150 32002
rect 57150 31950 57202 32002
rect 57202 31950 57204 32002
rect 57148 31948 57204 31950
rect 56588 31612 56644 31668
rect 58156 31890 58212 31892
rect 58156 31838 58158 31890
rect 58158 31838 58210 31890
rect 58210 31838 58212 31890
rect 58156 31836 58212 31838
rect 57596 30268 57652 30324
rect 55692 28754 55748 28756
rect 55692 28702 55694 28754
rect 55694 28702 55746 28754
rect 55746 28702 55748 28754
rect 55692 28700 55748 28702
rect 54572 27916 54628 27972
rect 54684 28476 54740 28532
rect 53452 26572 53508 26628
rect 53900 25900 53956 25956
rect 53452 24668 53508 24724
rect 51996 21532 52052 21588
rect 51996 20524 52052 20580
rect 53900 23938 53956 23940
rect 53900 23886 53902 23938
rect 53902 23886 53954 23938
rect 53954 23886 53956 23938
rect 53900 23884 53956 23886
rect 54124 23884 54180 23940
rect 54460 25676 54516 25732
rect 55356 27970 55412 27972
rect 55356 27918 55358 27970
rect 55358 27918 55410 27970
rect 55410 27918 55412 27970
rect 55356 27916 55412 27918
rect 54908 27858 54964 27860
rect 54908 27806 54910 27858
rect 54910 27806 54962 27858
rect 54962 27806 54964 27858
rect 54908 27804 54964 27806
rect 54908 25900 54964 25956
rect 55356 25954 55412 25956
rect 55356 25902 55358 25954
rect 55358 25902 55410 25954
rect 55410 25902 55412 25954
rect 55356 25900 55412 25902
rect 56700 25954 56756 25956
rect 56700 25902 56702 25954
rect 56702 25902 56754 25954
rect 56754 25902 56756 25954
rect 56700 25900 56756 25902
rect 54908 25116 54964 25172
rect 55804 25116 55860 25172
rect 56700 24722 56756 24724
rect 56700 24670 56702 24722
rect 56702 24670 56754 24722
rect 56754 24670 56756 24722
rect 56700 24668 56756 24670
rect 55692 24332 55748 24388
rect 57484 24386 57540 24388
rect 57484 24334 57486 24386
rect 57486 24334 57538 24386
rect 57538 24334 57540 24386
rect 57484 24332 57540 24334
rect 57148 23938 57204 23940
rect 57148 23886 57150 23938
rect 57150 23886 57202 23938
rect 57202 23886 57204 23938
rect 57148 23884 57204 23886
rect 53564 21810 53620 21812
rect 53564 21758 53566 21810
rect 53566 21758 53618 21810
rect 53618 21758 53620 21810
rect 53564 21756 53620 21758
rect 53564 20578 53620 20580
rect 53564 20526 53566 20578
rect 53566 20526 53618 20578
rect 53618 20526 53620 20578
rect 53564 20524 53620 20526
rect 52780 19964 52836 20020
rect 51884 18620 51940 18676
rect 52668 18620 52724 18676
rect 51996 18508 52052 18564
rect 50092 16434 50148 16436
rect 50092 16382 50094 16434
rect 50094 16382 50146 16434
rect 50146 16382 50148 16434
rect 50092 16380 50148 16382
rect 49644 16268 49700 16324
rect 50540 16268 50596 16324
rect 50556 16154 50612 16156
rect 50556 16102 50558 16154
rect 50558 16102 50610 16154
rect 50610 16102 50612 16154
rect 50556 16100 50612 16102
rect 50660 16154 50716 16156
rect 50660 16102 50662 16154
rect 50662 16102 50714 16154
rect 50714 16102 50716 16154
rect 50660 16100 50716 16102
rect 50764 16154 50820 16156
rect 50764 16102 50766 16154
rect 50766 16102 50818 16154
rect 50818 16102 50820 16154
rect 50764 16100 50820 16102
rect 50092 15874 50148 15876
rect 50092 15822 50094 15874
rect 50094 15822 50146 15874
rect 50146 15822 50148 15874
rect 50092 15820 50148 15822
rect 49868 15596 49924 15652
rect 51100 15986 51156 15988
rect 51100 15934 51102 15986
rect 51102 15934 51154 15986
rect 51154 15934 51156 15986
rect 51100 15932 51156 15934
rect 51212 16380 51268 16436
rect 50988 15874 51044 15876
rect 50988 15822 50990 15874
rect 50990 15822 51042 15874
rect 51042 15822 51044 15874
rect 50988 15820 51044 15822
rect 50540 14588 50596 14644
rect 47068 14476 47124 14532
rect 46396 12402 46452 12404
rect 46396 12350 46398 12402
rect 46398 12350 46450 12402
rect 46450 12350 46452 12402
rect 46396 12348 46452 12350
rect 45388 10780 45444 10836
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 54124 20466 54180 20468
rect 54124 20414 54126 20466
rect 54126 20414 54178 20466
rect 54178 20414 54180 20466
rect 54124 20412 54180 20414
rect 53340 19794 53396 19796
rect 53340 19742 53342 19794
rect 53342 19742 53394 19794
rect 53394 19742 53396 19794
rect 53340 19740 53396 19742
rect 52892 18508 52948 18564
rect 53228 18562 53284 18564
rect 53228 18510 53230 18562
rect 53230 18510 53282 18562
rect 53282 18510 53284 18562
rect 53228 18508 53284 18510
rect 54348 18620 54404 18676
rect 56700 23602 56756 23604
rect 56700 23550 56702 23602
rect 56702 23550 56754 23602
rect 56754 23550 56756 23602
rect 56700 23548 56756 23550
rect 57932 24668 57988 24724
rect 57596 23548 57652 23604
rect 55020 22428 55076 22484
rect 56476 22482 56532 22484
rect 56476 22430 56478 22482
rect 56478 22430 56530 22482
rect 56530 22430 56532 22482
rect 56476 22428 56532 22430
rect 56700 21810 56756 21812
rect 56700 21758 56702 21810
rect 56702 21758 56754 21810
rect 56754 21758 56756 21810
rect 56700 21756 56756 21758
rect 54796 20972 54852 21028
rect 54908 20524 54964 20580
rect 54796 19964 54852 20020
rect 54572 19740 54628 19796
rect 54124 18508 54180 18564
rect 53676 17890 53732 17892
rect 53676 17838 53678 17890
rect 53678 17838 53730 17890
rect 53730 17838 53732 17890
rect 53676 17836 53732 17838
rect 51212 15484 51268 15540
rect 51884 15538 51940 15540
rect 51884 15486 51886 15538
rect 51886 15486 51938 15538
rect 51938 15486 51940 15538
rect 51884 15484 51940 15486
rect 51548 14252 51604 14308
rect 52108 16434 52164 16436
rect 52108 16382 52110 16434
rect 52110 16382 52162 16434
rect 52162 16382 52164 16434
rect 52108 16380 52164 16382
rect 52332 16268 52388 16324
rect 52108 15820 52164 15876
rect 51996 14252 52052 14308
rect 53452 17612 53508 17668
rect 53228 16380 53284 16436
rect 53004 15762 53060 15764
rect 53004 15710 53006 15762
rect 53006 15710 53058 15762
rect 53058 15710 53060 15762
rect 53004 15708 53060 15710
rect 54124 16492 54180 16548
rect 53676 16268 53732 16324
rect 53900 16380 53956 16436
rect 52668 14700 52724 14756
rect 52892 14642 52948 14644
rect 52892 14590 52894 14642
rect 52894 14590 52946 14642
rect 52946 14590 52948 14642
rect 52892 14588 52948 14590
rect 52668 14252 52724 14308
rect 52556 13804 52612 13860
rect 55468 20524 55524 20580
rect 56476 21026 56532 21028
rect 56476 20974 56478 21026
rect 56478 20974 56530 21026
rect 56530 20974 56532 21026
rect 56476 20972 56532 20974
rect 57820 23884 57876 23940
rect 57708 21756 57764 21812
rect 55916 20690 55972 20692
rect 55916 20638 55918 20690
rect 55918 20638 55970 20690
rect 55970 20638 55972 20690
rect 55916 20636 55972 20638
rect 56812 20636 56868 20692
rect 55692 20412 55748 20468
rect 56700 20412 56756 20468
rect 55132 19740 55188 19796
rect 54684 18620 54740 18676
rect 56924 18508 56980 18564
rect 57708 18562 57764 18564
rect 57708 18510 57710 18562
rect 57710 18510 57762 18562
rect 57762 18510 57764 18562
rect 57708 18508 57764 18510
rect 54572 16658 54628 16660
rect 54572 16606 54574 16658
rect 54574 16606 54626 16658
rect 54626 16606 54628 16658
rect 54572 16604 54628 16606
rect 54236 15596 54292 15652
rect 54460 16492 54516 16548
rect 54908 16380 54964 16436
rect 55020 16604 55076 16660
rect 54460 15484 54516 15540
rect 54572 13858 54628 13860
rect 54572 13806 54574 13858
rect 54574 13806 54626 13858
rect 54626 13806 54628 13858
rect 54572 13804 54628 13806
rect 55580 16658 55636 16660
rect 55580 16606 55582 16658
rect 55582 16606 55634 16658
rect 55634 16606 55636 16658
rect 55580 16604 55636 16606
rect 56140 16658 56196 16660
rect 56140 16606 56142 16658
rect 56142 16606 56194 16658
rect 56194 16606 56196 16658
rect 56140 16604 56196 16606
rect 55356 16492 55412 16548
rect 56588 16546 56644 16548
rect 56588 16494 56590 16546
rect 56590 16494 56642 16546
rect 56642 16494 56644 16546
rect 56588 16492 56644 16494
rect 55132 16268 55188 16324
rect 48860 12348 48916 12404
rect 50556 12122 50612 12124
rect 50556 12070 50558 12122
rect 50558 12070 50610 12122
rect 50610 12070 50612 12122
rect 50556 12068 50612 12070
rect 50660 12122 50716 12124
rect 50660 12070 50662 12122
rect 50662 12070 50714 12122
rect 50714 12070 50716 12122
rect 50660 12068 50716 12070
rect 50764 12122 50820 12124
rect 50764 12070 50766 12122
rect 50766 12070 50818 12122
rect 50818 12070 50820 12122
rect 50764 12068 50820 12070
rect 52780 12738 52836 12740
rect 52780 12686 52782 12738
rect 52782 12686 52834 12738
rect 52834 12686 52836 12738
rect 52780 12684 52836 12686
rect 51884 11676 51940 11732
rect 53340 11730 53396 11732
rect 53340 11678 53342 11730
rect 53342 11678 53394 11730
rect 53394 11678 53396 11730
rect 53340 11676 53396 11678
rect 48860 11564 48916 11620
rect 52332 11618 52388 11620
rect 52332 11566 52334 11618
rect 52334 11566 52386 11618
rect 52386 11566 52388 11618
rect 52332 11564 52388 11566
rect 53116 11564 53172 11620
rect 56252 14754 56308 14756
rect 56252 14702 56254 14754
rect 56254 14702 56306 14754
rect 56306 14702 56308 14754
rect 56252 14700 56308 14702
rect 57484 16268 57540 16324
rect 56028 13858 56084 13860
rect 56028 13806 56030 13858
rect 56030 13806 56082 13858
rect 56082 13806 56084 13858
rect 56028 13804 56084 13806
rect 55356 12684 55412 12740
rect 53676 11564 53732 11620
rect 50556 10106 50612 10108
rect 50556 10054 50558 10106
rect 50558 10054 50610 10106
rect 50610 10054 50612 10106
rect 50556 10052 50612 10054
rect 50660 10106 50716 10108
rect 50660 10054 50662 10106
rect 50662 10054 50714 10106
rect 50714 10054 50716 10106
rect 50660 10052 50716 10054
rect 50764 10106 50820 10108
rect 50764 10054 50766 10106
rect 50766 10054 50818 10106
rect 50818 10054 50820 10106
rect 50764 10052 50820 10054
rect 31612 7868 31668 7924
rect 29596 7810 29652 7812
rect 29596 7758 29598 7810
rect 29598 7758 29650 7810
rect 29650 7758 29652 7810
rect 29596 7756 29652 7758
rect 30380 7756 30436 7812
rect 29148 7698 29204 7700
rect 29148 7646 29150 7698
rect 29150 7646 29202 7698
rect 29202 7646 29204 7698
rect 29148 7644 29204 7646
rect 30268 7586 30324 7588
rect 30268 7534 30270 7586
rect 30270 7534 30322 7586
rect 30322 7534 30324 7586
rect 30268 7532 30324 7534
rect 30604 7698 30660 7700
rect 30604 7646 30606 7698
rect 30606 7646 30658 7698
rect 30658 7646 30660 7698
rect 30604 7644 30660 7646
rect 31836 7868 31892 7924
rect 50556 8090 50612 8092
rect 50556 8038 50558 8090
rect 50558 8038 50610 8090
rect 50610 8038 50612 8090
rect 50556 8036 50612 8038
rect 50660 8090 50716 8092
rect 50660 8038 50662 8090
rect 50662 8038 50714 8090
rect 50714 8038 50716 8090
rect 50660 8036 50716 8038
rect 50764 8090 50820 8092
rect 50764 8038 50766 8090
rect 50766 8038 50818 8090
rect 50818 8038 50820 8090
rect 50764 8036 50820 8038
rect 31724 7532 31780 7588
rect 4284 7420 4340 7476
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 3836 6748 3892 6804
rect 19836 6074 19892 6076
rect 19836 6022 19838 6074
rect 19838 6022 19890 6074
rect 19890 6022 19892 6074
rect 19836 6020 19892 6022
rect 19940 6074 19996 6076
rect 19940 6022 19942 6074
rect 19942 6022 19994 6074
rect 19994 6022 19996 6074
rect 19940 6020 19996 6022
rect 20044 6074 20100 6076
rect 20044 6022 20046 6074
rect 20046 6022 20098 6074
rect 20098 6022 20100 6074
rect 20044 6020 20100 6022
rect 50556 6074 50612 6076
rect 50556 6022 50558 6074
rect 50558 6022 50610 6074
rect 50610 6022 50612 6074
rect 50556 6020 50612 6022
rect 50660 6074 50716 6076
rect 50660 6022 50662 6074
rect 50662 6022 50714 6074
rect 50714 6022 50716 6074
rect 50660 6020 50716 6022
rect 50764 6074 50820 6076
rect 50764 6022 50766 6074
rect 50766 6022 50818 6074
rect 50818 6022 50820 6074
rect 50764 6020 50820 6022
rect 4476 5066 4532 5068
rect 4476 5014 4478 5066
rect 4478 5014 4530 5066
rect 4530 5014 4532 5066
rect 4476 5012 4532 5014
rect 4580 5066 4636 5068
rect 4580 5014 4582 5066
rect 4582 5014 4634 5066
rect 4634 5014 4636 5066
rect 4580 5012 4636 5014
rect 4684 5066 4740 5068
rect 4684 5014 4686 5066
rect 4686 5014 4738 5066
rect 4738 5014 4740 5066
rect 4684 5012 4740 5014
rect 35196 5066 35252 5068
rect 35196 5014 35198 5066
rect 35198 5014 35250 5066
rect 35250 5014 35252 5066
rect 35196 5012 35252 5014
rect 35300 5066 35356 5068
rect 35300 5014 35302 5066
rect 35302 5014 35354 5066
rect 35354 5014 35356 5066
rect 35300 5012 35356 5014
rect 35404 5066 35460 5068
rect 35404 5014 35406 5066
rect 35406 5014 35458 5066
rect 35458 5014 35460 5066
rect 35404 5012 35460 5014
rect 19836 4058 19892 4060
rect 19836 4006 19838 4058
rect 19838 4006 19890 4058
rect 19890 4006 19892 4058
rect 19836 4004 19892 4006
rect 19940 4058 19996 4060
rect 19940 4006 19942 4058
rect 19942 4006 19994 4058
rect 19994 4006 19996 4058
rect 19940 4004 19996 4006
rect 20044 4058 20100 4060
rect 20044 4006 20046 4058
rect 20046 4006 20098 4058
rect 20098 4006 20100 4058
rect 20044 4004 20100 4006
rect 50556 4058 50612 4060
rect 50556 4006 50558 4058
rect 50558 4006 50610 4058
rect 50610 4006 50612 4058
rect 50556 4004 50612 4006
rect 50660 4058 50716 4060
rect 50660 4006 50662 4058
rect 50662 4006 50714 4058
rect 50714 4006 50716 4058
rect 50660 4004 50716 4006
rect 50764 4058 50820 4060
rect 50764 4006 50766 4058
rect 50766 4006 50818 4058
rect 50818 4006 50820 4058
rect 50764 4004 50820 4006
<< metal3 >>
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4466 55412 4476 55468
rect 4532 55412 4580 55468
rect 4636 55412 4684 55468
rect 4740 55412 4750 55468
rect 35186 55412 35196 55468
rect 35252 55412 35300 55468
rect 35356 55412 35404 55468
rect 35460 55412 35470 55468
rect 19826 54404 19836 54460
rect 19892 54404 19940 54460
rect 19996 54404 20044 54460
rect 20100 54404 20110 54460
rect 50546 54404 50556 54460
rect 50612 54404 50660 54460
rect 50716 54404 50764 54460
rect 50820 54404 50830 54460
rect 0 53844 800 53872
rect 59200 53844 60000 53872
rect 0 53788 3836 53844
rect 3892 53788 3902 53844
rect 56130 53788 56140 53844
rect 56196 53788 60000 53844
rect 0 53760 800 53788
rect 59200 53760 60000 53788
rect 4466 53396 4476 53452
rect 4532 53396 4580 53452
rect 4636 53396 4684 53452
rect 4740 53396 4750 53452
rect 35186 53396 35196 53452
rect 35252 53396 35300 53452
rect 35356 53396 35404 53452
rect 35460 53396 35470 53452
rect 19826 52388 19836 52444
rect 19892 52388 19940 52444
rect 19996 52388 20044 52444
rect 20100 52388 20110 52444
rect 50546 52388 50556 52444
rect 50612 52388 50660 52444
rect 50716 52388 50764 52444
rect 50820 52388 50830 52444
rect 4466 51380 4476 51436
rect 4532 51380 4580 51436
rect 4636 51380 4684 51436
rect 4740 51380 4750 51436
rect 35186 51380 35196 51436
rect 35252 51380 35300 51436
rect 35356 51380 35404 51436
rect 35460 51380 35470 51436
rect 19826 50372 19836 50428
rect 19892 50372 19940 50428
rect 19996 50372 20044 50428
rect 20100 50372 20110 50428
rect 50546 50372 50556 50428
rect 50612 50372 50660 50428
rect 50716 50372 50764 50428
rect 50820 50372 50830 50428
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 36978 48860 36988 48916
rect 37044 48860 39228 48916
rect 39284 48860 39294 48916
rect 23090 48748 23100 48804
rect 23156 48748 24332 48804
rect 24388 48748 24398 48804
rect 25218 48748 25228 48804
rect 25284 48748 31948 48804
rect 32004 48748 32014 48804
rect 38770 48748 38780 48804
rect 38836 48748 40684 48804
rect 40740 48748 40750 48804
rect 41356 48748 42588 48804
rect 42644 48748 43596 48804
rect 43652 48748 43662 48804
rect 41356 48692 41412 48748
rect 38322 48636 38332 48692
rect 38388 48636 39004 48692
rect 39060 48636 41356 48692
rect 41412 48636 41422 48692
rect 19826 48356 19836 48412
rect 19892 48356 19940 48412
rect 19996 48356 20044 48412
rect 20100 48356 20110 48412
rect 50546 48356 50556 48412
rect 50612 48356 50660 48412
rect 50716 48356 50764 48412
rect 50820 48356 50830 48412
rect 26002 47964 26012 48020
rect 26068 47964 28140 48020
rect 28196 47964 28476 48020
rect 28532 47964 28542 48020
rect 19506 47852 19516 47908
rect 19572 47852 20188 47908
rect 20244 47852 20254 47908
rect 50642 47740 50652 47796
rect 50708 47740 53452 47796
rect 53508 47740 53518 47796
rect 4466 47348 4476 47404
rect 4532 47348 4580 47404
rect 4636 47348 4684 47404
rect 4740 47348 4750 47404
rect 35186 47348 35196 47404
rect 35252 47348 35300 47404
rect 35356 47348 35404 47404
rect 35460 47348 35470 47404
rect 20178 47180 20188 47236
rect 20244 47180 21644 47236
rect 21700 47180 21710 47236
rect 20626 47068 20636 47124
rect 20692 47068 23660 47124
rect 23716 47068 23726 47124
rect 21858 46956 21868 47012
rect 21924 46956 22876 47012
rect 22932 46956 22942 47012
rect 23538 46956 23548 47012
rect 23604 46956 26908 47012
rect 26964 46956 32060 47012
rect 32116 46956 32620 47012
rect 32676 46956 34188 47012
rect 34244 46956 34860 47012
rect 34916 46956 34926 47012
rect 22418 46844 22428 46900
rect 22484 46844 23996 46900
rect 24052 46844 24220 46900
rect 24276 46844 24286 46900
rect 28578 46844 28588 46900
rect 28644 46844 29372 46900
rect 29428 46844 29438 46900
rect 32284 46844 33068 46900
rect 33124 46844 34076 46900
rect 34132 46844 36988 46900
rect 37044 46844 37548 46900
rect 37604 46844 41020 46900
rect 41076 46844 41086 46900
rect 32284 46788 32340 46844
rect 28242 46732 28252 46788
rect 28308 46732 29820 46788
rect 29876 46732 32340 46788
rect 32498 46732 32508 46788
rect 32564 46732 40684 46788
rect 40740 46732 43820 46788
rect 43876 46732 43886 46788
rect 31892 46620 32060 46676
rect 32116 46620 32126 46676
rect 33170 46620 33180 46676
rect 33236 46620 35196 46676
rect 35252 46620 35262 46676
rect 43362 46620 43372 46676
rect 43428 46620 44044 46676
rect 44100 46620 44110 46676
rect 19826 46340 19836 46396
rect 19892 46340 19940 46396
rect 19996 46340 20044 46396
rect 20100 46340 20110 46396
rect 31892 46228 31948 46620
rect 50546 46340 50556 46396
rect 50612 46340 50660 46396
rect 50716 46340 50764 46396
rect 50820 46340 50830 46396
rect 24546 46172 24556 46228
rect 24612 46172 25116 46228
rect 25172 46172 26460 46228
rect 26516 46172 27356 46228
rect 27412 46172 27692 46228
rect 27748 46172 30604 46228
rect 30660 46172 31948 46228
rect 32274 46172 32284 46228
rect 32340 46172 34524 46228
rect 34580 46172 34590 46228
rect 43698 46172 43708 46228
rect 43764 46172 44044 46228
rect 44100 46172 45164 46228
rect 45220 46172 45230 46228
rect 20514 46060 20524 46116
rect 20580 46060 22652 46116
rect 22708 46060 23324 46116
rect 23380 46060 23390 46116
rect 24210 46060 24220 46116
rect 24276 46060 25452 46116
rect 25508 46060 25518 46116
rect 31938 46060 31948 46116
rect 32004 46060 32508 46116
rect 32564 46060 32574 46116
rect 43922 46060 43932 46116
rect 43988 46060 46172 46116
rect 46228 46060 46238 46116
rect 31042 45948 31052 46004
rect 31108 45948 33068 46004
rect 33124 45948 33134 46004
rect 40114 45948 40124 46004
rect 40180 45948 40348 46004
rect 40404 45948 41132 46004
rect 41188 45948 42812 46004
rect 42868 45948 42878 46004
rect 53778 45948 53788 46004
rect 53844 45948 54908 46004
rect 54964 45948 55356 46004
rect 55412 45948 55422 46004
rect 31490 45836 31500 45892
rect 31556 45836 33740 45892
rect 33796 45836 33806 45892
rect 48066 45836 48076 45892
rect 48132 45836 49420 45892
rect 49476 45836 49486 45892
rect 25218 45724 25228 45780
rect 25284 45724 27244 45780
rect 27300 45724 27310 45780
rect 39554 45500 39564 45556
rect 39620 45500 43372 45556
rect 43428 45500 43438 45556
rect 42130 45388 42140 45444
rect 42196 45388 49756 45444
rect 49812 45388 49822 45444
rect 50082 45388 50092 45444
rect 50148 45388 50316 45444
rect 50372 45388 52556 45444
rect 52612 45388 54124 45444
rect 54180 45388 54190 45444
rect 4466 45332 4476 45388
rect 4532 45332 4580 45388
rect 4636 45332 4684 45388
rect 4740 45332 4750 45388
rect 35186 45332 35196 45388
rect 35252 45332 35300 45388
rect 35356 45332 35404 45388
rect 35460 45332 35470 45388
rect 17490 45276 17500 45332
rect 17556 45276 17948 45332
rect 18004 45276 20188 45332
rect 20244 45276 21308 45332
rect 21364 45276 21374 45332
rect 36978 45276 36988 45332
rect 37044 45276 37884 45332
rect 37940 45276 37950 45332
rect 40226 45276 40236 45332
rect 40292 45276 42588 45332
rect 42644 45276 42654 45332
rect 49074 45276 49084 45332
rect 49140 45276 52668 45332
rect 52724 45276 52734 45332
rect 52322 45164 52332 45220
rect 52388 45164 53452 45220
rect 53508 45164 53518 45220
rect 32610 45052 32620 45108
rect 32676 45052 35308 45108
rect 35364 45052 35374 45108
rect 29138 44940 29148 44996
rect 29204 44940 32396 44996
rect 32452 44940 34076 44996
rect 34132 44940 34524 44996
rect 34580 44940 34590 44996
rect 37538 44940 37548 44996
rect 37604 44940 37996 44996
rect 38052 44940 38062 44996
rect 17154 44828 17164 44884
rect 17220 44828 17612 44884
rect 17668 44828 18060 44884
rect 18116 44828 18126 44884
rect 34178 44828 34188 44884
rect 34244 44828 36092 44884
rect 36148 44828 36876 44884
rect 36932 44828 36942 44884
rect 43698 44828 43708 44884
rect 43764 44828 44044 44884
rect 44100 44828 44716 44884
rect 44772 44828 44782 44884
rect 50194 44828 50204 44884
rect 50260 44828 50988 44884
rect 51044 44828 51054 44884
rect 53666 44828 53676 44884
rect 53732 44828 54796 44884
rect 54852 44828 54862 44884
rect 44146 44716 44156 44772
rect 44212 44716 45052 44772
rect 45108 44716 46620 44772
rect 46676 44716 46686 44772
rect 50866 44716 50876 44772
rect 50932 44716 51212 44772
rect 51268 44716 51278 44772
rect 51874 44716 51884 44772
rect 51940 44716 52668 44772
rect 52724 44716 52734 44772
rect 21746 44604 21756 44660
rect 21812 44604 23772 44660
rect 23828 44604 23838 44660
rect 27794 44604 27804 44660
rect 27860 44604 28252 44660
rect 28308 44604 28700 44660
rect 28756 44604 28766 44660
rect 49634 44604 49644 44660
rect 49700 44604 50652 44660
rect 50708 44604 50718 44660
rect 51426 44604 51436 44660
rect 51492 44604 53116 44660
rect 53172 44604 53182 44660
rect 19826 44324 19836 44380
rect 19892 44324 19940 44380
rect 19996 44324 20044 44380
rect 20100 44324 20110 44380
rect 50546 44324 50556 44380
rect 50612 44324 50660 44380
rect 50716 44324 50764 44380
rect 50820 44324 50830 44380
rect 43474 44268 43484 44324
rect 43540 44268 43932 44324
rect 43988 44268 43998 44324
rect 33618 44044 33628 44100
rect 33684 44044 34188 44100
rect 34244 44044 34254 44100
rect 42690 44044 42700 44100
rect 42756 44044 43484 44100
rect 43540 44044 44156 44100
rect 44212 44044 44222 44100
rect 29026 43932 29036 43988
rect 29092 43932 30268 43988
rect 30324 43932 31724 43988
rect 31780 43932 32172 43988
rect 32228 43932 33404 43988
rect 33460 43932 33470 43988
rect 51874 43932 51884 43988
rect 51940 43932 53340 43988
rect 53396 43932 53406 43988
rect 54002 43932 54012 43988
rect 54068 43932 54684 43988
rect 54740 43932 56700 43988
rect 56756 43932 57148 43988
rect 57204 43932 57214 43988
rect 19618 43820 19628 43876
rect 19684 43820 24332 43876
rect 24388 43820 27020 43876
rect 27076 43820 27086 43876
rect 37986 43820 37996 43876
rect 38052 43820 39452 43876
rect 39508 43820 39518 43876
rect 50866 43820 50876 43876
rect 50932 43820 52332 43876
rect 52388 43820 52892 43876
rect 52948 43820 52958 43876
rect 18050 43708 18060 43764
rect 18116 43708 21532 43764
rect 21588 43708 21598 43764
rect 25666 43708 25676 43764
rect 25732 43708 26124 43764
rect 26180 43708 26190 43764
rect 30156 43708 32060 43764
rect 32116 43708 32126 43764
rect 38098 43708 38108 43764
rect 38164 43708 39564 43764
rect 39620 43708 39630 43764
rect 40338 43708 40348 43764
rect 40404 43708 41020 43764
rect 41076 43708 41086 43764
rect 41458 43708 41468 43764
rect 41524 43708 43260 43764
rect 43316 43708 43326 43764
rect 48626 43708 48636 43764
rect 48692 43708 49532 43764
rect 49588 43708 50204 43764
rect 50260 43708 50270 43764
rect 23426 43596 23436 43652
rect 23492 43596 24108 43652
rect 24164 43596 24556 43652
rect 24612 43596 24622 43652
rect 27234 43596 27244 43652
rect 27300 43596 28140 43652
rect 28196 43596 28206 43652
rect 30156 43428 30212 43708
rect 43922 43596 43932 43652
rect 43988 43596 45164 43652
rect 45220 43596 47404 43652
rect 47460 43596 47470 43652
rect 40114 43484 40124 43540
rect 40180 43484 40796 43540
rect 40852 43484 40862 43540
rect 24658 43372 24668 43428
rect 24724 43372 30212 43428
rect 4466 43316 4476 43372
rect 4532 43316 4580 43372
rect 4636 43316 4684 43372
rect 4740 43316 4750 43372
rect 35186 43316 35196 43372
rect 35252 43316 35300 43372
rect 35356 43316 35404 43372
rect 35460 43316 35470 43372
rect 43026 43260 43036 43316
rect 43092 43260 44940 43316
rect 44996 43260 45006 43316
rect 43586 43148 43596 43204
rect 43652 43148 45164 43204
rect 45220 43148 45230 43204
rect 33282 43036 33292 43092
rect 33348 43036 33964 43092
rect 34020 43036 34030 43092
rect 42802 43036 42812 43092
rect 42868 43036 45388 43092
rect 45444 43036 45454 43092
rect 27234 42924 27244 42980
rect 27300 42924 29036 42980
rect 29092 42924 29102 42980
rect 36866 42924 36876 42980
rect 36932 42924 39228 42980
rect 39284 42924 39294 42980
rect 53116 42924 56140 42980
rect 56196 42924 56206 42980
rect 53116 42868 53172 42924
rect 20626 42812 20636 42868
rect 20692 42812 23100 42868
rect 23156 42812 23166 42868
rect 28018 42812 28028 42868
rect 28084 42812 32956 42868
rect 33012 42812 34636 42868
rect 34692 42812 37772 42868
rect 37828 42812 38668 42868
rect 39666 42812 39676 42868
rect 39732 42812 41020 42868
rect 41076 42812 41086 42868
rect 41234 42812 41244 42868
rect 41300 42812 42588 42868
rect 42644 42812 42654 42868
rect 43250 42812 43260 42868
rect 43316 42812 43596 42868
rect 43652 42812 46396 42868
rect 46452 42812 47628 42868
rect 47684 42812 49756 42868
rect 49812 42812 50204 42868
rect 50260 42812 53116 42868
rect 53172 42812 53182 42868
rect 54450 42812 54460 42868
rect 54516 42812 55132 42868
rect 55188 42812 55198 42868
rect 55412 42812 56028 42868
rect 56084 42812 56476 42868
rect 56532 42812 56542 42868
rect 38612 42756 38668 42812
rect 28130 42700 28140 42756
rect 28196 42700 29596 42756
rect 29652 42700 29662 42756
rect 38612 42700 39228 42756
rect 39284 42700 39294 42756
rect 40226 42700 40236 42756
rect 40292 42700 45612 42756
rect 45668 42700 45678 42756
rect 54226 42700 54236 42756
rect 54292 42700 55020 42756
rect 55076 42700 55356 42756
rect 55412 42700 55468 42812
rect 55682 42700 55692 42756
rect 55748 42700 56924 42756
rect 56980 42700 56990 42756
rect 55692 42644 55748 42700
rect 9762 42588 9772 42644
rect 9828 42588 10668 42644
rect 10724 42588 10734 42644
rect 41906 42588 41916 42644
rect 41972 42588 42700 42644
rect 42756 42588 43148 42644
rect 43204 42588 43214 42644
rect 46834 42588 46844 42644
rect 46900 42588 47404 42644
rect 47460 42588 48188 42644
rect 48244 42588 49420 42644
rect 49476 42588 49486 42644
rect 51986 42588 51996 42644
rect 52052 42588 53452 42644
rect 53508 42588 55748 42644
rect 56130 42588 56140 42644
rect 56196 42588 57372 42644
rect 57428 42588 57438 42644
rect 42354 42476 42364 42532
rect 42420 42476 44716 42532
rect 44772 42476 44782 42532
rect 55794 42476 55804 42532
rect 55860 42476 56700 42532
rect 56756 42476 56766 42532
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 21970 42140 21980 42196
rect 22036 42140 22764 42196
rect 22820 42140 26796 42196
rect 26852 42140 29372 42196
rect 29428 42140 33404 42196
rect 33460 42140 33470 42196
rect 50530 42140 50540 42196
rect 50596 42140 53676 42196
rect 53732 42140 53742 42196
rect 29698 42028 29708 42084
rect 29764 42028 34468 42084
rect 49074 42028 49084 42084
rect 49140 42028 50876 42084
rect 50932 42028 51212 42084
rect 51268 42028 51548 42084
rect 51604 42028 54348 42084
rect 54404 42028 54414 42084
rect 34412 41972 34468 42028
rect 52220 41972 52276 42028
rect 53564 41972 53620 42028
rect 8082 41916 8092 41972
rect 8148 41916 8988 41972
rect 9044 41916 9660 41972
rect 9716 41916 9726 41972
rect 19282 41916 19292 41972
rect 19348 41916 20468 41972
rect 21634 41916 21644 41972
rect 21700 41916 22092 41972
rect 22148 41916 22158 41972
rect 24098 41916 24108 41972
rect 24164 41916 27468 41972
rect 27524 41916 27534 41972
rect 30258 41916 30268 41972
rect 30324 41916 33852 41972
rect 33908 41916 33918 41972
rect 34402 41916 34412 41972
rect 34468 41916 35756 41972
rect 35812 41916 36316 41972
rect 36372 41916 38892 41972
rect 38948 41916 39788 41972
rect 39844 41916 41244 41972
rect 41300 41916 41692 41972
rect 41748 41916 41758 41972
rect 52210 41916 52220 41972
rect 52276 41916 52286 41972
rect 53554 41916 53564 41972
rect 53620 41916 53630 41972
rect 4610 41804 4620 41860
rect 4676 41804 6188 41860
rect 6244 41804 6254 41860
rect 10994 41804 11004 41860
rect 11060 41804 12124 41860
rect 12180 41804 12190 41860
rect 20412 41748 20468 41916
rect 21858 41804 21868 41860
rect 21924 41804 22316 41860
rect 22372 41804 25116 41860
rect 25172 41804 25182 41860
rect 27122 41804 27132 41860
rect 27188 41804 28476 41860
rect 28532 41804 28542 41860
rect 33954 41804 33964 41860
rect 34020 41804 35532 41860
rect 35588 41804 36428 41860
rect 36484 41804 37772 41860
rect 37828 41804 37838 41860
rect 44594 41804 44604 41860
rect 44660 41804 46620 41860
rect 46676 41804 50092 41860
rect 50148 41804 51996 41860
rect 52052 41804 52062 41860
rect 1810 41692 1820 41748
rect 1876 41692 3724 41748
rect 3780 41692 3790 41748
rect 20402 41692 20412 41748
rect 20468 41692 21980 41748
rect 22036 41692 22046 41748
rect 22764 41692 24668 41748
rect 24724 41692 25676 41748
rect 25732 41692 26796 41748
rect 26852 41692 26862 41748
rect 28130 41692 28140 41748
rect 28196 41692 28812 41748
rect 28868 41692 30940 41748
rect 30996 41692 31006 41748
rect 41346 41692 41356 41748
rect 41412 41692 42140 41748
rect 42196 41692 42206 41748
rect 51314 41692 51324 41748
rect 51380 41692 52332 41748
rect 52388 41692 52398 41748
rect 56130 41692 56140 41748
rect 56196 41692 57148 41748
rect 57204 41692 57214 41748
rect 22764 41636 22820 41692
rect 6290 41580 6300 41636
rect 6356 41580 7196 41636
rect 7252 41580 7262 41636
rect 19506 41580 19516 41636
rect 19572 41580 20748 41636
rect 20804 41580 22764 41636
rect 22820 41580 22830 41636
rect 23874 41580 23884 41636
rect 23940 41580 25564 41636
rect 25620 41580 25630 41636
rect 50418 41580 50428 41636
rect 50484 41580 53788 41636
rect 53844 41580 54796 41636
rect 54852 41580 55804 41636
rect 55860 41580 55870 41636
rect 9538 41468 9548 41524
rect 9604 41468 10892 41524
rect 10948 41468 10958 41524
rect 34738 41468 34748 41524
rect 34804 41468 41468 41524
rect 41524 41468 41534 41524
rect 4466 41300 4476 41356
rect 4532 41300 4580 41356
rect 4636 41300 4684 41356
rect 4740 41300 4750 41356
rect 35186 41300 35196 41356
rect 35252 41300 35300 41356
rect 35356 41300 35404 41356
rect 35460 41300 35470 41356
rect 20402 41020 20412 41076
rect 20468 41020 22092 41076
rect 22148 41020 25452 41076
rect 25508 41020 28028 41076
rect 28084 41020 28094 41076
rect 19842 40908 19852 40964
rect 19908 40908 20188 40964
rect 20244 40908 20254 40964
rect 18274 40796 18284 40852
rect 18340 40796 19292 40852
rect 19348 40796 20300 40852
rect 20356 40796 21308 40852
rect 21364 40796 24220 40852
rect 24276 40796 25788 40852
rect 25844 40796 25854 40852
rect 34962 40796 34972 40852
rect 35028 40796 36428 40852
rect 36484 40796 38444 40852
rect 38500 40796 38510 40852
rect 38770 40796 38780 40852
rect 38836 40796 39564 40852
rect 39620 40796 39630 40852
rect 47068 40796 47964 40852
rect 48020 40796 48030 40852
rect 49410 40796 49420 40852
rect 49476 40796 53004 40852
rect 53060 40796 53070 40852
rect 47068 40740 47124 40796
rect 3714 40684 3724 40740
rect 3780 40684 4620 40740
rect 4676 40684 4686 40740
rect 20738 40684 20748 40740
rect 20804 40684 22316 40740
rect 22372 40684 22382 40740
rect 35970 40684 35980 40740
rect 36036 40684 37884 40740
rect 37940 40684 37950 40740
rect 40338 40684 40348 40740
rect 40404 40684 41356 40740
rect 41412 40684 47068 40740
rect 47124 40684 47134 40740
rect 47730 40684 47740 40740
rect 47796 40684 49532 40740
rect 49588 40684 49598 40740
rect 6850 40572 6860 40628
rect 6916 40572 8652 40628
rect 8708 40572 10220 40628
rect 10276 40572 10286 40628
rect 49074 40572 49084 40628
rect 49140 40572 53676 40628
rect 53732 40572 53742 40628
rect 1810 40460 1820 40516
rect 1876 40460 2716 40516
rect 2772 40460 5628 40516
rect 5684 40460 5694 40516
rect 6290 40460 6300 40516
rect 6356 40460 7532 40516
rect 7588 40460 7868 40516
rect 7924 40460 7934 40516
rect 37090 40460 37100 40516
rect 37156 40460 37996 40516
rect 38052 40460 39676 40516
rect 39732 40460 42028 40516
rect 42084 40460 43596 40516
rect 43652 40460 43662 40516
rect 49186 40460 49196 40516
rect 49252 40460 49756 40516
rect 49812 40460 50204 40516
rect 50260 40460 50270 40516
rect 50428 40460 50540 40516
rect 50596 40460 50606 40516
rect 0 40404 800 40432
rect 0 40348 1708 40404
rect 1764 40348 1774 40404
rect 2370 40348 2380 40404
rect 2436 40348 4060 40404
rect 4116 40348 6076 40404
rect 6132 40348 6142 40404
rect 24770 40348 24780 40404
rect 24836 40348 27916 40404
rect 27972 40348 27982 40404
rect 0 40320 800 40348
rect 19826 40292 19836 40348
rect 19892 40292 19940 40348
rect 19996 40292 20044 40348
rect 20100 40292 20110 40348
rect 50428 40292 50484 40460
rect 50546 40292 50556 40348
rect 50612 40292 50660 40348
rect 50716 40292 50764 40348
rect 50820 40292 50830 40348
rect 24098 40236 24108 40292
rect 24164 40236 24556 40292
rect 24612 40236 30380 40292
rect 30436 40236 30446 40292
rect 31826 40236 31836 40292
rect 31892 40068 31948 40292
rect 35186 40236 35196 40292
rect 35252 40236 36988 40292
rect 37044 40236 37054 40292
rect 43922 40236 43932 40292
rect 43988 40236 45500 40292
rect 45556 40236 49420 40292
rect 49476 40236 50484 40292
rect 34850 40124 34860 40180
rect 34916 40124 35980 40180
rect 36036 40124 36046 40180
rect 43586 40124 43596 40180
rect 43652 40124 44940 40180
rect 44996 40124 45276 40180
rect 45332 40124 46396 40180
rect 46452 40124 46462 40180
rect 7970 40012 7980 40068
rect 8036 40012 8876 40068
rect 8932 40012 8942 40068
rect 11778 40012 11788 40068
rect 11844 40012 12572 40068
rect 12628 40012 12638 40068
rect 20132 39956 20188 40068
rect 20244 40012 20254 40068
rect 21634 40012 21644 40068
rect 21700 40012 23772 40068
rect 23828 40012 23838 40068
rect 31892 40012 35084 40068
rect 35140 40012 35150 40068
rect 38434 40012 38444 40068
rect 38500 40012 39228 40068
rect 39284 40012 40236 40068
rect 40292 40012 40302 40068
rect 41906 40012 41916 40068
rect 41972 40012 44492 40068
rect 44548 40012 45388 40068
rect 45444 40012 46508 40068
rect 46564 40012 46574 40068
rect 49970 40012 49980 40068
rect 50036 40012 53900 40068
rect 53956 40012 53966 40068
rect 17154 39900 17164 39956
rect 17220 39900 20860 39956
rect 20916 39900 21532 39956
rect 21588 39900 22540 39956
rect 22596 39900 22606 39956
rect 24658 39900 24668 39956
rect 24724 39900 26348 39956
rect 26404 39900 26414 39956
rect 33506 39900 33516 39956
rect 33572 39900 36540 39956
rect 36596 39900 37324 39956
rect 37380 39900 39788 39956
rect 39844 39900 39854 39956
rect 37986 39788 37996 39844
rect 38052 39788 41020 39844
rect 41076 39788 41086 39844
rect 41458 39788 41468 39844
rect 41524 39788 42140 39844
rect 42196 39788 42206 39844
rect 48178 39788 48188 39844
rect 48244 39788 50764 39844
rect 50820 39788 51996 39844
rect 52052 39788 52062 39844
rect 24434 39676 24444 39732
rect 24500 39676 25452 39732
rect 25508 39676 25518 39732
rect 30706 39676 30716 39732
rect 30772 39676 31164 39732
rect 31220 39676 31230 39732
rect 34066 39676 34076 39732
rect 34132 39676 37324 39732
rect 37380 39676 37390 39732
rect 39778 39676 39788 39732
rect 39844 39676 40460 39732
rect 40516 39676 42476 39732
rect 42532 39676 42542 39732
rect 44034 39676 44044 39732
rect 44100 39676 46732 39732
rect 46788 39676 46798 39732
rect 44044 39620 44100 39676
rect 4946 39564 4956 39620
rect 5012 39564 6188 39620
rect 6244 39564 6254 39620
rect 9650 39564 9660 39620
rect 9716 39564 10332 39620
rect 10388 39564 13356 39620
rect 13412 39564 13422 39620
rect 38770 39564 38780 39620
rect 38836 39564 42140 39620
rect 42196 39564 44100 39620
rect 47506 39564 47516 39620
rect 47572 39564 49308 39620
rect 49364 39564 49374 39620
rect 4466 39284 4476 39340
rect 4532 39284 4580 39340
rect 4636 39284 4684 39340
rect 4740 39284 4750 39340
rect 35186 39284 35196 39340
rect 35252 39284 35300 39340
rect 35356 39284 35404 39340
rect 35460 39284 35470 39340
rect 37314 39004 37324 39060
rect 37380 39004 39452 39060
rect 39508 39004 39518 39060
rect 40226 39004 40236 39060
rect 40292 39004 42420 39060
rect 42364 38948 42420 39004
rect 2370 38892 2380 38948
rect 2436 38892 5628 38948
rect 5684 38892 5694 38948
rect 10210 38892 10220 38948
rect 10276 38892 13468 38948
rect 13524 38892 13534 38948
rect 38546 38892 38556 38948
rect 38612 38892 40572 38948
rect 40628 38892 41916 38948
rect 41972 38892 41982 38948
rect 42354 38892 42364 38948
rect 42420 38892 48188 38948
rect 48244 38892 48254 38948
rect 51986 38892 51996 38948
rect 52052 38892 52780 38948
rect 52836 38892 52846 38948
rect 55570 38892 55580 38948
rect 55636 38892 56476 38948
rect 56532 38892 56542 38948
rect 23650 38780 23660 38836
rect 23716 38780 25900 38836
rect 25956 38780 25966 38836
rect 37202 38780 37212 38836
rect 37268 38780 39116 38836
rect 39172 38780 39182 38836
rect 39442 38780 39452 38836
rect 39508 38780 40796 38836
rect 40852 38780 40862 38836
rect 44594 38780 44604 38836
rect 44660 38780 48636 38836
rect 48692 38780 48702 38836
rect 50194 38780 50204 38836
rect 50260 38780 50428 38836
rect 50484 38780 50494 38836
rect 4946 38668 4956 38724
rect 5012 38668 5740 38724
rect 5796 38668 5806 38724
rect 6636 38668 8652 38724
rect 8708 38668 8718 38724
rect 12786 38668 12796 38724
rect 12852 38668 13580 38724
rect 13636 38668 13646 38724
rect 16818 38668 16828 38724
rect 16884 38668 17612 38724
rect 17668 38668 19852 38724
rect 19908 38668 20916 38724
rect 25330 38668 25340 38724
rect 25396 38668 27356 38724
rect 27412 38668 29932 38724
rect 29988 38668 29998 38724
rect 40226 38668 40236 38724
rect 40292 38668 41132 38724
rect 41188 38668 41198 38724
rect 42578 38668 42588 38724
rect 42644 38668 44940 38724
rect 44996 38668 45006 38724
rect 46498 38668 46508 38724
rect 46564 38668 47628 38724
rect 47684 38668 47694 38724
rect 48178 38668 48188 38724
rect 48244 38668 50764 38724
rect 50820 38668 50830 38724
rect 52098 38668 52108 38724
rect 52164 38668 53788 38724
rect 53844 38668 54684 38724
rect 54740 38668 56028 38724
rect 56084 38668 56094 38724
rect 6636 38612 6692 38668
rect 20860 38612 20916 38668
rect 6626 38556 6636 38612
rect 6692 38556 6702 38612
rect 20178 38556 20188 38612
rect 20244 38556 20636 38612
rect 20692 38556 20702 38612
rect 20850 38556 20860 38612
rect 20916 38556 20926 38612
rect 33506 38556 33516 38612
rect 33572 38556 34412 38612
rect 34468 38556 34478 38612
rect 35522 38556 35532 38612
rect 35588 38556 36316 38612
rect 36372 38556 36382 38612
rect 49746 38556 49756 38612
rect 49812 38556 51100 38612
rect 51156 38556 51166 38612
rect 49074 38444 49084 38500
rect 49140 38444 50652 38500
rect 50708 38444 51772 38500
rect 51828 38444 51838 38500
rect 19826 38276 19836 38332
rect 19892 38276 19940 38332
rect 19996 38276 20044 38332
rect 20100 38276 20110 38332
rect 50546 38276 50556 38332
rect 50612 38276 50660 38332
rect 50716 38276 50764 38332
rect 50820 38276 50830 38332
rect 4834 37996 4844 38052
rect 4900 37996 5740 38052
rect 5796 37996 6300 38052
rect 6356 37996 6636 38052
rect 6692 37996 6702 38052
rect 21634 37996 21644 38052
rect 21700 37996 23100 38052
rect 23156 37996 23772 38052
rect 23828 37996 25228 38052
rect 25284 37996 25294 38052
rect 32162 37996 32172 38052
rect 32228 37996 33180 38052
rect 33236 37996 33246 38052
rect 38220 37996 41580 38052
rect 41636 37996 43036 38052
rect 43092 37996 43102 38052
rect 46386 37996 46396 38052
rect 46452 37996 47740 38052
rect 47796 37996 49756 38052
rect 49812 37996 49822 38052
rect 38220 37716 38276 37996
rect 38546 37884 38556 37940
rect 38612 37884 38892 37940
rect 38948 37884 38958 37940
rect 40450 37884 40460 37940
rect 40516 37884 43260 37940
rect 43316 37884 43326 37940
rect 48178 37884 48188 37940
rect 48244 37884 49084 37940
rect 49140 37884 49150 37940
rect 51538 37772 51548 37828
rect 51604 37772 52892 37828
rect 52948 37772 52958 37828
rect 24210 37660 24220 37716
rect 24276 37660 25564 37716
rect 25620 37660 25630 37716
rect 30258 37660 30268 37716
rect 30324 37660 31052 37716
rect 31108 37660 31118 37716
rect 36306 37660 36316 37716
rect 36372 37660 37660 37716
rect 37716 37660 38220 37716
rect 38276 37660 38286 37716
rect 9650 37548 9660 37604
rect 9716 37548 10780 37604
rect 10836 37548 13804 37604
rect 13860 37548 13870 37604
rect 37090 37548 37100 37604
rect 37156 37548 38556 37604
rect 38612 37548 38622 37604
rect 41346 37548 41356 37604
rect 41412 37548 42700 37604
rect 42756 37548 42766 37604
rect 4466 37268 4476 37324
rect 4532 37268 4580 37324
rect 4636 37268 4684 37324
rect 4740 37268 4750 37324
rect 35186 37268 35196 37324
rect 35252 37268 35300 37324
rect 35356 37268 35404 37324
rect 35460 37268 35470 37324
rect 18162 37100 18172 37156
rect 18228 37100 20188 37156
rect 20244 37100 20254 37156
rect 49074 37100 49084 37156
rect 49140 37100 54348 37156
rect 54404 37100 54414 37156
rect 41234 36988 41244 37044
rect 41300 36988 41972 37044
rect 41916 36932 41972 36988
rect 1810 36876 1820 36932
rect 1876 36876 2716 36932
rect 2772 36876 4508 36932
rect 4564 36876 4574 36932
rect 9314 36876 9324 36932
rect 9380 36876 9884 36932
rect 9940 36876 9950 36932
rect 16706 36876 16716 36932
rect 16772 36876 20188 36932
rect 20244 36876 21644 36932
rect 21700 36876 23100 36932
rect 23156 36876 24220 36932
rect 24276 36876 24286 36932
rect 41916 36876 42588 36932
rect 42644 36876 42654 36932
rect 53106 36876 53116 36932
rect 53172 36876 53788 36932
rect 53844 36876 54348 36932
rect 54404 36876 54414 36932
rect 3602 36764 3612 36820
rect 3668 36764 5068 36820
rect 5124 36764 6076 36820
rect 6132 36764 6142 36820
rect 20738 36764 20748 36820
rect 20804 36764 21868 36820
rect 21924 36764 21934 36820
rect 3042 36652 3052 36708
rect 3108 36652 3836 36708
rect 3892 36652 5628 36708
rect 5684 36652 5694 36708
rect 19506 36652 19516 36708
rect 19572 36652 20860 36708
rect 20916 36652 24444 36708
rect 24500 36652 24510 36708
rect 24668 36652 26012 36708
rect 26068 36652 28420 36708
rect 37762 36652 37772 36708
rect 37828 36652 38556 36708
rect 38612 36652 38622 36708
rect 41234 36652 41244 36708
rect 41300 36652 45164 36708
rect 45220 36652 45230 36708
rect 50866 36652 50876 36708
rect 50932 36652 52780 36708
rect 52836 36652 52846 36708
rect 54114 36652 54124 36708
rect 54180 36652 55804 36708
rect 55860 36652 57148 36708
rect 57204 36652 57214 36708
rect 24668 36596 24724 36652
rect 28364 36596 28420 36652
rect 12786 36540 12796 36596
rect 12852 36540 13580 36596
rect 13636 36540 13646 36596
rect 18722 36540 18732 36596
rect 18788 36540 21196 36596
rect 21252 36540 21262 36596
rect 21858 36540 21868 36596
rect 21924 36540 23548 36596
rect 23604 36540 23996 36596
rect 24052 36540 24668 36596
rect 24724 36540 24734 36596
rect 25890 36540 25900 36596
rect 25956 36540 27356 36596
rect 27412 36540 27422 36596
rect 28354 36540 28364 36596
rect 28420 36540 29260 36596
rect 29316 36540 29326 36596
rect 46722 36540 46732 36596
rect 46788 36540 47852 36596
rect 47908 36540 50204 36596
rect 50260 36540 50316 36596
rect 50372 36540 51212 36596
rect 51268 36540 51278 36596
rect 10210 36428 10220 36484
rect 10276 36428 11340 36484
rect 11396 36428 13468 36484
rect 13524 36428 13534 36484
rect 26450 36428 26460 36484
rect 26516 36428 27916 36484
rect 27972 36428 27982 36484
rect 38882 36428 38892 36484
rect 38948 36428 41468 36484
rect 41524 36428 41534 36484
rect 0 36372 800 36400
rect 0 36316 4172 36372
rect 4228 36316 4238 36372
rect 0 36288 800 36316
rect 19826 36260 19836 36316
rect 19892 36260 19940 36316
rect 19996 36260 20044 36316
rect 20100 36260 20110 36316
rect 50546 36260 50556 36316
rect 50612 36260 50660 36316
rect 50716 36260 50764 36316
rect 50820 36260 50830 36316
rect 18386 36092 18396 36148
rect 18452 36092 19180 36148
rect 19236 36092 19246 36148
rect 19618 36092 19628 36148
rect 19684 36092 20636 36148
rect 20692 36092 20702 36148
rect 18834 35980 18844 36036
rect 18900 35980 19852 36036
rect 19908 35980 20748 36036
rect 20804 35980 20814 36036
rect 36194 35980 36204 36036
rect 36260 35980 37772 36036
rect 37828 35980 37838 36036
rect 55906 35980 55916 36036
rect 55972 35980 56700 36036
rect 56756 35980 56766 36036
rect 9874 35868 9884 35924
rect 9940 35868 11004 35924
rect 11060 35868 13020 35924
rect 13076 35868 14140 35924
rect 14196 35868 15260 35924
rect 15316 35868 16380 35924
rect 16436 35868 16446 35924
rect 37090 35868 37100 35924
rect 37156 35868 38332 35924
rect 38388 35868 38398 35924
rect 49410 35868 49420 35924
rect 49476 35868 50204 35924
rect 50260 35868 50270 35924
rect 24546 35756 24556 35812
rect 24612 35756 26348 35812
rect 26404 35756 27020 35812
rect 27076 35756 27086 35812
rect 29810 35756 29820 35812
rect 29876 35756 31836 35812
rect 31892 35756 40348 35812
rect 40404 35756 41244 35812
rect 41300 35756 42700 35812
rect 42756 35756 42766 35812
rect 53106 35756 53116 35812
rect 53172 35756 53900 35812
rect 53956 35756 53966 35812
rect 0 35700 800 35728
rect 27020 35700 27076 35756
rect 0 35644 16380 35700
rect 16436 35644 17724 35700
rect 17780 35644 18620 35700
rect 18676 35644 21420 35700
rect 21476 35644 21486 35700
rect 27020 35644 30604 35700
rect 30660 35644 30670 35700
rect 31378 35644 31388 35700
rect 31444 35644 33180 35700
rect 33236 35644 33516 35700
rect 33572 35644 34076 35700
rect 34132 35644 34142 35700
rect 41682 35644 41692 35700
rect 41748 35644 42364 35700
rect 42420 35644 44492 35700
rect 44548 35644 44558 35700
rect 48962 35644 48972 35700
rect 49028 35644 50092 35700
rect 50148 35644 51436 35700
rect 51492 35644 51502 35700
rect 0 35616 800 35644
rect 31388 35588 31444 35644
rect 29474 35532 29484 35588
rect 29540 35532 31444 35588
rect 38322 35532 38332 35588
rect 38388 35532 40124 35588
rect 40180 35532 40190 35588
rect 32722 35308 32732 35364
rect 32788 35308 34748 35364
rect 34804 35308 34814 35364
rect 43652 35308 43708 35364
rect 43764 35308 43774 35364
rect 44034 35308 44044 35364
rect 44100 35308 44940 35364
rect 44996 35308 45836 35364
rect 45892 35308 45902 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 43652 35252 43764 35308
rect 25666 35196 25676 35252
rect 25732 35196 26908 35252
rect 26964 35196 26974 35252
rect 27570 35196 27580 35252
rect 27636 35196 29708 35252
rect 29764 35196 29774 35252
rect 41794 35196 41804 35252
rect 41860 35196 44380 35252
rect 44436 35196 44446 35252
rect 51874 35196 51884 35252
rect 51940 35196 53004 35252
rect 53060 35196 53070 35252
rect 3378 35084 3388 35140
rect 3444 35084 5628 35140
rect 5684 35084 6300 35140
rect 6356 35084 6366 35140
rect 11890 35084 11900 35140
rect 11956 35084 13468 35140
rect 13524 35084 13534 35140
rect 14140 35084 16828 35140
rect 16884 35084 20188 35140
rect 20244 35084 20254 35140
rect 35298 35084 35308 35140
rect 35364 35084 35644 35140
rect 35700 35084 44268 35140
rect 44324 35084 44828 35140
rect 44884 35084 44894 35140
rect 0 35028 800 35056
rect 14140 35028 14196 35084
rect 0 34972 14196 35028
rect 51874 34972 51884 35028
rect 51940 34972 52556 35028
rect 52612 34972 53340 35028
rect 53396 34972 53406 35028
rect 0 34944 800 34972
rect 20412 34860 21644 34916
rect 21700 34860 21980 34916
rect 22036 34860 22046 34916
rect 42924 34860 44044 34916
rect 44100 34860 44110 34916
rect 44706 34860 44716 34916
rect 44772 34860 44940 34916
rect 44996 34860 46060 34916
rect 46116 34860 47180 34916
rect 47236 34860 48188 34916
rect 48244 34860 49420 34916
rect 49476 34860 49486 34916
rect 51202 34860 51212 34916
rect 51268 34860 52780 34916
rect 52836 34860 52846 34916
rect 52994 34860 53004 34916
rect 53060 34860 53788 34916
rect 53844 34860 54684 34916
rect 54740 34860 54750 34916
rect 55412 34860 56140 34916
rect 56196 34860 56206 34916
rect 20412 34804 20468 34860
rect 924 34748 20412 34804
rect 20468 34748 20478 34804
rect 21522 34748 21532 34804
rect 21588 34748 22876 34804
rect 22932 34748 23324 34804
rect 23380 34748 23390 34804
rect 26674 34748 26684 34804
rect 26740 34748 28028 34804
rect 28084 34748 29260 34804
rect 29316 34748 29326 34804
rect 33730 34748 33740 34804
rect 33796 34748 35196 34804
rect 35252 34748 36204 34804
rect 36260 34748 36270 34804
rect 37202 34748 37212 34804
rect 37268 34748 38108 34804
rect 38164 34748 38668 34804
rect 38724 34748 38734 34804
rect 0 34356 800 34384
rect 924 34356 980 34748
rect 4162 34636 4172 34692
rect 4228 34636 16604 34692
rect 16660 34636 19628 34692
rect 19684 34636 21308 34692
rect 21364 34636 22428 34692
rect 22484 34636 23772 34692
rect 23828 34636 23838 34692
rect 34850 34636 34860 34692
rect 34916 34636 35532 34692
rect 35588 34636 35598 34692
rect 42924 34580 42980 34860
rect 53004 34804 53060 34860
rect 55412 34804 55468 34860
rect 48850 34748 48860 34804
rect 48916 34748 49868 34804
rect 49924 34748 50652 34804
rect 50708 34748 51324 34804
rect 51380 34748 52108 34804
rect 52164 34748 53060 34804
rect 54898 34748 54908 34804
rect 54964 34748 55468 34804
rect 43652 34636 44492 34692
rect 44548 34636 49980 34692
rect 50036 34636 51548 34692
rect 51604 34636 52332 34692
rect 52388 34636 52398 34692
rect 55682 34636 55692 34692
rect 55748 34636 56588 34692
rect 56644 34636 56654 34692
rect 43652 34580 43708 34636
rect 3714 34524 3724 34580
rect 3780 34524 5740 34580
rect 5796 34524 5806 34580
rect 24658 34524 24668 34580
rect 24724 34524 26124 34580
rect 26180 34524 26190 34580
rect 28354 34524 28364 34580
rect 28420 34524 29372 34580
rect 29428 34524 29438 34580
rect 37650 34524 37660 34580
rect 37716 34524 41804 34580
rect 41860 34524 42924 34580
rect 42980 34524 42990 34580
rect 43138 34524 43148 34580
rect 43204 34524 43708 34580
rect 0 34300 980 34356
rect 22306 34300 22316 34356
rect 22372 34300 25340 34356
rect 25396 34300 25406 34356
rect 0 34272 800 34300
rect 19826 34244 19836 34300
rect 19892 34244 19940 34300
rect 19996 34244 20044 34300
rect 20100 34244 20110 34300
rect 50546 34244 50556 34300
rect 50612 34244 50660 34300
rect 50716 34244 50764 34300
rect 50820 34244 50830 34300
rect 23202 34076 23212 34132
rect 23268 34076 24108 34132
rect 24164 34076 24668 34132
rect 24724 34076 24734 34132
rect 55010 34076 55020 34132
rect 55076 34076 55692 34132
rect 55748 34076 55758 34132
rect 3266 33964 3276 34020
rect 3332 33964 4060 34020
rect 4116 33964 4126 34020
rect 20178 33964 20188 34020
rect 20244 33964 20860 34020
rect 20916 33964 21756 34020
rect 21812 33964 21822 34020
rect 24882 33964 24892 34020
rect 24948 33964 26236 34020
rect 26292 33964 26684 34020
rect 26740 33964 26750 34020
rect 38322 33964 38332 34020
rect 38388 33964 40348 34020
rect 40404 33964 40414 34020
rect 42252 33964 44716 34020
rect 44772 33964 44782 34020
rect 51538 33964 51548 34020
rect 51604 33964 54012 34020
rect 54068 33964 54078 34020
rect 42252 33908 42308 33964
rect 15092 33852 16380 33908
rect 16436 33852 18172 33908
rect 18228 33852 18844 33908
rect 18900 33852 20468 33908
rect 20962 33852 20972 33908
rect 21028 33852 22652 33908
rect 22708 33852 23660 33908
rect 23716 33852 23726 33908
rect 25778 33852 25788 33908
rect 25844 33852 27356 33908
rect 27412 33852 27916 33908
rect 27972 33852 27982 33908
rect 31826 33852 31836 33908
rect 31892 33852 37212 33908
rect 37268 33852 37278 33908
rect 41010 33852 41020 33908
rect 41076 33852 42252 33908
rect 42308 33852 42318 33908
rect 52770 33852 52780 33908
rect 52836 33852 54348 33908
rect 54404 33852 54414 33908
rect 5730 33740 5740 33796
rect 5796 33740 6412 33796
rect 6468 33740 6860 33796
rect 6916 33740 6926 33796
rect 0 33684 800 33712
rect 15092 33684 15148 33852
rect 20412 33796 20468 33852
rect 19170 33740 19180 33796
rect 19236 33740 20188 33796
rect 20244 33740 20254 33796
rect 20412 33740 30716 33796
rect 30772 33740 31276 33796
rect 31332 33740 31342 33796
rect 42354 33740 42364 33796
rect 42420 33740 43484 33796
rect 43540 33740 44268 33796
rect 44324 33740 44334 33796
rect 45714 33740 45724 33796
rect 45780 33740 46620 33796
rect 46676 33740 48860 33796
rect 48916 33740 48926 33796
rect 51874 33740 51884 33796
rect 51940 33740 52892 33796
rect 52948 33740 52958 33796
rect 0 33628 15148 33684
rect 16370 33628 16380 33684
rect 16436 33628 17948 33684
rect 18004 33628 18014 33684
rect 18946 33628 18956 33684
rect 19012 33628 19740 33684
rect 19796 33628 21420 33684
rect 21476 33628 21486 33684
rect 21644 33628 23548 33684
rect 23604 33628 24108 33684
rect 24164 33628 25116 33684
rect 25172 33628 25182 33684
rect 32386 33628 32396 33684
rect 32452 33628 34300 33684
rect 34356 33628 35308 33684
rect 35364 33628 35374 33684
rect 41346 33628 41356 33684
rect 41412 33628 43708 33684
rect 43764 33628 45164 33684
rect 45220 33628 46732 33684
rect 46788 33628 46798 33684
rect 53890 33628 53900 33684
rect 53956 33628 55804 33684
rect 55860 33628 55870 33684
rect 0 33600 800 33628
rect 21644 33572 21700 33628
rect 12226 33516 12236 33572
rect 12292 33516 14028 33572
rect 14084 33516 14094 33572
rect 21634 33516 21644 33572
rect 21700 33516 21710 33572
rect 49858 33404 49868 33460
rect 49924 33404 52220 33460
rect 52276 33404 52286 33460
rect 4466 33236 4476 33292
rect 4532 33236 4580 33292
rect 4636 33236 4684 33292
rect 4740 33236 4750 33292
rect 35186 33236 35196 33292
rect 35252 33236 35300 33292
rect 35356 33236 35404 33292
rect 35460 33236 35470 33292
rect 0 33012 800 33040
rect 0 32956 16940 33012
rect 16996 32956 19516 33012
rect 19572 32956 22092 33012
rect 22148 32956 28588 33012
rect 28644 32956 29484 33012
rect 29540 32956 29550 33012
rect 35746 32956 35756 33012
rect 35812 32956 47292 33012
rect 47348 32956 47358 33012
rect 0 32928 800 32956
rect 25890 32844 25900 32900
rect 25956 32844 29820 32900
rect 29876 32844 31164 32900
rect 31220 32844 31230 32900
rect 52658 32844 52668 32900
rect 52724 32844 53788 32900
rect 53844 32844 53854 32900
rect 20626 32732 20636 32788
rect 20692 32732 22204 32788
rect 22260 32732 22270 32788
rect 24322 32732 24332 32788
rect 24388 32732 25340 32788
rect 25396 32732 25406 32788
rect 25554 32732 25564 32788
rect 25620 32732 30268 32788
rect 30324 32732 30334 32788
rect 39778 32732 39788 32788
rect 39844 32732 43932 32788
rect 43988 32732 45276 32788
rect 45332 32732 45342 32788
rect 45714 32732 45724 32788
rect 45780 32732 47068 32788
rect 47124 32732 47134 32788
rect 22204 32676 22260 32732
rect 13570 32620 13580 32676
rect 13636 32620 20300 32676
rect 20356 32620 20366 32676
rect 22204 32620 25900 32676
rect 25956 32620 25966 32676
rect 30482 32620 30492 32676
rect 30548 32620 31276 32676
rect 31332 32620 31342 32676
rect 34066 32620 34076 32676
rect 34132 32620 35532 32676
rect 35588 32620 37100 32676
rect 37156 32620 37166 32676
rect 38882 32620 38892 32676
rect 38948 32620 40572 32676
rect 40628 32620 41020 32676
rect 41076 32620 41086 32676
rect 50978 32620 50988 32676
rect 51044 32620 55020 32676
rect 55076 32620 55086 32676
rect 3826 32508 3836 32564
rect 3892 32508 5628 32564
rect 5684 32508 5694 32564
rect 10882 32508 10892 32564
rect 10948 32508 13468 32564
rect 13524 32508 13534 32564
rect 22418 32508 22428 32564
rect 22484 32508 24668 32564
rect 24724 32508 24734 32564
rect 24882 32508 24892 32564
rect 24948 32508 26012 32564
rect 26068 32508 26078 32564
rect 37314 32508 37324 32564
rect 37380 32508 40460 32564
rect 40516 32508 40526 32564
rect 42018 32508 42028 32564
rect 42084 32508 42588 32564
rect 42644 32508 50204 32564
rect 50260 32508 51100 32564
rect 51156 32508 51166 32564
rect 53890 32508 53900 32564
rect 53956 32508 54124 32564
rect 54180 32508 54190 32564
rect 49298 32396 49308 32452
rect 49364 32396 50988 32452
rect 51044 32396 51054 32452
rect 0 32340 800 32368
rect 0 32284 7532 32340
rect 7588 32284 7598 32340
rect 0 32256 800 32284
rect 19826 32228 19836 32284
rect 19892 32228 19940 32284
rect 19996 32228 20044 32284
rect 20100 32228 20110 32284
rect 50546 32228 50556 32284
rect 50612 32228 50660 32284
rect 50716 32228 50764 32284
rect 50820 32228 50830 32284
rect 25218 32060 25228 32116
rect 25284 32060 26460 32116
rect 26516 32060 26526 32116
rect 8866 31948 8876 32004
rect 8932 31948 9772 32004
rect 9828 31948 9838 32004
rect 14130 31948 14140 32004
rect 14196 31948 17724 32004
rect 17780 31948 20188 32004
rect 20244 31948 20254 32004
rect 54114 31948 54124 32004
rect 54180 31948 57148 32004
rect 57204 31948 57214 32004
rect 12898 31836 12908 31892
rect 12964 31836 13804 31892
rect 13860 31836 13870 31892
rect 15362 31836 15372 31892
rect 15428 31836 19516 31892
rect 19572 31836 19582 31892
rect 22866 31836 22876 31892
rect 22932 31836 24220 31892
rect 24276 31836 25228 31892
rect 25284 31836 26348 31892
rect 26404 31836 29372 31892
rect 29428 31836 29438 31892
rect 34626 31836 34636 31892
rect 34692 31836 35644 31892
rect 35700 31836 35710 31892
rect 38994 31836 39004 31892
rect 39060 31836 41244 31892
rect 41300 31836 42140 31892
rect 42196 31836 43036 31892
rect 43092 31836 43102 31892
rect 51538 31836 51548 31892
rect 51604 31836 51884 31892
rect 51940 31836 56028 31892
rect 56084 31836 56094 31892
rect 56690 31836 56700 31892
rect 56756 31836 58156 31892
rect 58212 31836 58222 31892
rect 3378 31724 3388 31780
rect 3444 31724 4172 31780
rect 4228 31724 4238 31780
rect 6290 31724 6300 31780
rect 6356 31724 6972 31780
rect 7028 31724 7038 31780
rect 7410 31724 7420 31780
rect 7476 31724 8764 31780
rect 8820 31724 8830 31780
rect 15698 31724 15708 31780
rect 15764 31724 16380 31780
rect 16436 31724 17388 31780
rect 17444 31724 17454 31780
rect 24658 31724 24668 31780
rect 24724 31724 26012 31780
rect 26068 31724 26078 31780
rect 33506 31724 33516 31780
rect 33572 31724 36652 31780
rect 36708 31724 36718 31780
rect 38434 31724 38444 31780
rect 38500 31724 46060 31780
rect 46116 31724 46126 31780
rect 47954 31724 47964 31780
rect 48020 31724 50092 31780
rect 50148 31724 50158 31780
rect 51426 31724 51436 31780
rect 51492 31724 53900 31780
rect 53956 31724 53966 31780
rect 55458 31724 55468 31780
rect 55524 31724 56476 31780
rect 56532 31724 57036 31780
rect 57092 31724 57102 31780
rect 0 31668 800 31696
rect 0 31612 14364 31668
rect 14420 31612 14430 31668
rect 19058 31612 19068 31668
rect 19124 31612 20188 31668
rect 20244 31612 20254 31668
rect 37762 31612 37772 31668
rect 37828 31612 38220 31668
rect 38276 31612 38556 31668
rect 38612 31612 39900 31668
rect 39956 31612 40908 31668
rect 40964 31612 40974 31668
rect 47842 31612 47852 31668
rect 47908 31612 48748 31668
rect 48804 31612 48814 31668
rect 55682 31612 55692 31668
rect 55748 31612 56588 31668
rect 56644 31612 56654 31668
rect 0 31584 800 31612
rect 35634 31500 35644 31556
rect 35700 31500 36988 31556
rect 37044 31500 37054 31556
rect 50306 31500 50316 31556
rect 50372 31500 51324 31556
rect 51380 31500 52444 31556
rect 52500 31500 54124 31556
rect 54180 31500 54190 31556
rect 6178 31388 6188 31444
rect 6244 31388 6860 31444
rect 6916 31388 7308 31444
rect 7364 31388 7374 31444
rect 7522 31388 7532 31444
rect 7588 31388 21308 31444
rect 21364 31388 22204 31444
rect 22260 31388 22988 31444
rect 23044 31388 23054 31444
rect 4466 31220 4476 31276
rect 4532 31220 4580 31276
rect 4636 31220 4684 31276
rect 4740 31220 4750 31276
rect 35186 31220 35196 31276
rect 35252 31220 35300 31276
rect 35356 31220 35404 31276
rect 35460 31220 35470 31276
rect 32610 31164 32620 31220
rect 32676 31164 33852 31220
rect 33908 31164 33918 31220
rect 25106 31052 25116 31108
rect 25172 31052 27916 31108
rect 27972 31052 28476 31108
rect 28532 31052 28542 31108
rect 30482 31052 30492 31108
rect 30548 31052 35756 31108
rect 35812 31052 35822 31108
rect 0 30996 800 31024
rect 0 30940 9996 30996
rect 10052 30940 10062 30996
rect 26002 30940 26012 30996
rect 26068 30940 28140 30996
rect 28196 30940 28206 30996
rect 36642 30940 36652 30996
rect 36708 30940 37324 30996
rect 37380 30940 38556 30996
rect 38612 30940 38622 30996
rect 49074 30940 49084 30996
rect 49140 30940 51548 30996
rect 51604 30940 52220 30996
rect 52276 30940 52286 30996
rect 0 30912 800 30940
rect 12898 30828 12908 30884
rect 12964 30828 14924 30884
rect 14980 30828 14990 30884
rect 27010 30828 27020 30884
rect 27076 30828 31164 30884
rect 31220 30828 31230 30884
rect 32050 30828 32060 30884
rect 32116 30828 32732 30884
rect 32788 30828 32798 30884
rect 33730 30828 33740 30884
rect 33796 30828 34972 30884
rect 35028 30828 35038 30884
rect 36978 30828 36988 30884
rect 37044 30828 39004 30884
rect 39060 30828 39070 30884
rect 32060 30772 32116 30828
rect 3714 30716 3724 30772
rect 3780 30716 6076 30772
rect 6132 30716 6142 30772
rect 12450 30716 12460 30772
rect 12516 30716 18620 30772
rect 18676 30716 18686 30772
rect 30146 30716 30156 30772
rect 30212 30716 30492 30772
rect 30548 30716 30558 30772
rect 30930 30716 30940 30772
rect 30996 30716 32116 30772
rect 32498 30716 32508 30772
rect 32564 30716 36428 30772
rect 36484 30716 37996 30772
rect 38052 30716 38062 30772
rect 40562 30716 40572 30772
rect 40628 30716 41132 30772
rect 41188 30716 47964 30772
rect 48020 30716 48030 30772
rect 2370 30604 2380 30660
rect 2436 30604 5516 30660
rect 5572 30604 5582 30660
rect 29474 30604 29484 30660
rect 29540 30604 29932 30660
rect 29988 30604 30604 30660
rect 30660 30604 31276 30660
rect 31332 30604 33516 30660
rect 33572 30604 33582 30660
rect 33852 30604 38388 30660
rect 39442 30604 39452 30660
rect 39508 30604 48972 30660
rect 49028 30604 49038 30660
rect 54450 30604 54460 30660
rect 54516 30604 55468 30660
rect 55524 30604 55534 30660
rect 4050 30492 4060 30548
rect 4116 30492 4620 30548
rect 4676 30492 7308 30548
rect 7364 30492 8316 30548
rect 8372 30492 8382 30548
rect 10546 30492 10556 30548
rect 10612 30492 11116 30548
rect 11172 30492 12124 30548
rect 12180 30492 12190 30548
rect 13234 30492 13244 30548
rect 13300 30492 14028 30548
rect 14084 30492 14700 30548
rect 14756 30492 14766 30548
rect 20402 30492 20412 30548
rect 20468 30492 21420 30548
rect 21476 30492 21486 30548
rect 32834 30492 32844 30548
rect 32900 30492 33628 30548
rect 33684 30492 33694 30548
rect 33852 30436 33908 30604
rect 34178 30492 34188 30548
rect 34244 30492 35084 30548
rect 35140 30492 35150 30548
rect 35252 30492 37548 30548
rect 37604 30492 37614 30548
rect 35252 30436 35308 30492
rect 8372 30380 16268 30436
rect 16324 30380 16334 30436
rect 24210 30380 24220 30436
rect 24276 30380 26684 30436
rect 26740 30380 27468 30436
rect 27524 30380 27534 30436
rect 28130 30380 28140 30436
rect 28196 30380 29148 30436
rect 29204 30380 29214 30436
rect 30034 30380 30044 30436
rect 30100 30380 30110 30436
rect 31826 30380 31836 30436
rect 31892 30380 33908 30436
rect 34962 30380 34972 30436
rect 35028 30380 35308 30436
rect 36194 30380 36204 30436
rect 36260 30380 38108 30436
rect 38164 30380 38174 30436
rect 0 30324 800 30352
rect 8372 30324 8428 30380
rect 30044 30324 30100 30380
rect 38332 30324 38388 30604
rect 38546 30492 38556 30548
rect 38612 30492 39228 30548
rect 39284 30492 39294 30548
rect 45490 30492 45500 30548
rect 45556 30492 48188 30548
rect 48244 30492 51660 30548
rect 51716 30492 51726 30548
rect 46274 30380 46284 30436
rect 46340 30380 46620 30436
rect 46676 30380 50652 30436
rect 50708 30380 54236 30436
rect 54292 30380 54302 30436
rect 0 30268 8428 30324
rect 11676 30268 14140 30324
rect 14196 30268 14206 30324
rect 25778 30268 25788 30324
rect 25844 30268 30100 30324
rect 32386 30268 32396 30324
rect 32452 30268 34300 30324
rect 34356 30268 34366 30324
rect 34738 30268 34748 30324
rect 34804 30268 35084 30324
rect 35140 30268 36652 30324
rect 36708 30268 36718 30324
rect 37314 30268 37324 30324
rect 37380 30268 37772 30324
rect 37828 30268 37838 30324
rect 38332 30268 49420 30324
rect 49476 30268 49486 30324
rect 53788 30268 53900 30324
rect 53956 30268 57596 30324
rect 57652 30268 57662 30324
rect 0 30240 800 30268
rect 11676 30212 11732 30268
rect 19826 30212 19836 30268
rect 19892 30212 19940 30268
rect 19996 30212 20044 30268
rect 20100 30212 20110 30268
rect 50546 30212 50556 30268
rect 50612 30212 50660 30268
rect 50716 30212 50764 30268
rect 50820 30212 50830 30268
rect 53788 30212 53844 30268
rect 11666 30156 11676 30212
rect 11732 30156 11742 30212
rect 24546 30156 24556 30212
rect 24612 30156 26460 30212
rect 26516 30156 26526 30212
rect 33954 30156 33964 30212
rect 34020 30156 35420 30212
rect 35476 30156 35486 30212
rect 39778 30156 39788 30212
rect 39844 30156 40236 30212
rect 40292 30156 40302 30212
rect 46722 30156 46732 30212
rect 46788 30156 48748 30212
rect 48804 30156 50316 30212
rect 50372 30156 50382 30212
rect 53116 30156 53844 30212
rect 50316 30100 50372 30156
rect 53116 30100 53172 30156
rect 9986 30044 9996 30100
rect 10052 30044 12124 30100
rect 12180 30044 12190 30100
rect 15026 30044 15036 30100
rect 15092 30044 15932 30100
rect 15988 30044 15998 30100
rect 19618 30044 19628 30100
rect 19684 30044 21420 30100
rect 21476 30044 21486 30100
rect 21868 30044 27020 30100
rect 27076 30044 27086 30100
rect 50316 30044 51772 30100
rect 51828 30044 53116 30100
rect 53172 30044 53182 30100
rect 1810 29932 1820 29988
rect 1876 29932 2828 29988
rect 2884 29932 4060 29988
rect 4116 29932 4126 29988
rect 21868 29876 21924 30044
rect 24434 29932 24444 29988
rect 24500 29932 25900 29988
rect 25956 29932 30716 29988
rect 30772 29932 30782 29988
rect 36082 29932 36092 29988
rect 36148 29932 37100 29988
rect 37156 29932 37548 29988
rect 37604 29932 37614 29988
rect 37874 29932 37884 29988
rect 37940 29932 45724 29988
rect 45780 29932 45790 29988
rect 11554 29820 11564 29876
rect 11620 29820 12572 29876
rect 12628 29820 12638 29876
rect 14914 29820 14924 29876
rect 14980 29820 21868 29876
rect 21924 29820 21934 29876
rect 24658 29820 24668 29876
rect 24724 29820 25676 29876
rect 25732 29820 25742 29876
rect 27122 29820 27132 29876
rect 27188 29820 33852 29876
rect 33908 29820 33918 29876
rect 38322 29820 38332 29876
rect 38388 29820 40908 29876
rect 40964 29820 40974 29876
rect 44370 29820 44380 29876
rect 44436 29820 45388 29876
rect 45444 29820 45454 29876
rect 16370 29708 16380 29764
rect 16436 29708 21196 29764
rect 21252 29708 21262 29764
rect 23090 29708 23100 29764
rect 23156 29708 26124 29764
rect 26180 29708 26190 29764
rect 26338 29708 26348 29764
rect 26404 29708 28364 29764
rect 28420 29708 28812 29764
rect 28868 29708 28878 29764
rect 33618 29708 33628 29764
rect 33684 29708 34748 29764
rect 34804 29708 34814 29764
rect 35970 29708 35980 29764
rect 36036 29708 37884 29764
rect 37940 29708 47068 29764
rect 47124 29708 47404 29764
rect 47460 29708 47470 29764
rect 0 29652 800 29680
rect 0 29596 15484 29652
rect 15540 29596 15550 29652
rect 17378 29596 17388 29652
rect 17444 29596 18060 29652
rect 18116 29596 21084 29652
rect 21140 29596 21150 29652
rect 33842 29596 33852 29652
rect 33908 29596 36764 29652
rect 36820 29596 36830 29652
rect 39666 29596 39676 29652
rect 39732 29596 40348 29652
rect 40404 29596 43260 29652
rect 43316 29596 43326 29652
rect 51202 29596 51212 29652
rect 51268 29596 51996 29652
rect 52052 29596 52332 29652
rect 52388 29596 54012 29652
rect 54068 29596 54078 29652
rect 0 29568 800 29596
rect 4946 29484 4956 29540
rect 5012 29484 5740 29540
rect 5796 29484 5806 29540
rect 31602 29484 31612 29540
rect 31668 29484 33180 29540
rect 33236 29484 33246 29540
rect 41122 29484 41132 29540
rect 41188 29484 44268 29540
rect 44324 29484 44334 29540
rect 21746 29372 21756 29428
rect 21812 29372 25228 29428
rect 25284 29372 25294 29428
rect 28466 29372 28476 29428
rect 28532 29372 28812 29428
rect 28868 29372 35980 29428
rect 36036 29372 36046 29428
rect 42130 29372 42140 29428
rect 42196 29372 44380 29428
rect 44436 29372 46396 29428
rect 46452 29372 46732 29428
rect 46788 29372 46798 29428
rect 36194 29260 36204 29316
rect 36260 29260 36652 29316
rect 36708 29260 36718 29316
rect 4466 29204 4476 29260
rect 4532 29204 4580 29260
rect 4636 29204 4684 29260
rect 4740 29204 4750 29260
rect 35186 29204 35196 29260
rect 35252 29204 35300 29260
rect 35356 29204 35404 29260
rect 35460 29204 35470 29260
rect 13122 29148 13132 29204
rect 13188 29148 19180 29204
rect 19236 29148 19246 29204
rect 19618 29148 19628 29204
rect 19684 29148 27132 29204
rect 27188 29148 27198 29204
rect 12898 29036 12908 29092
rect 12964 29036 14924 29092
rect 14980 29036 17388 29092
rect 17444 29036 17454 29092
rect 21186 29036 21196 29092
rect 21252 29036 26348 29092
rect 26404 29036 26414 29092
rect 26786 29036 26796 29092
rect 26852 29036 29484 29092
rect 29540 29036 29550 29092
rect 30706 29036 30716 29092
rect 30772 29036 31164 29092
rect 31220 29036 39788 29092
rect 39844 29036 39854 29092
rect 0 28980 800 29008
rect 0 28924 16940 28980
rect 16996 28924 17006 28980
rect 17602 28924 17612 28980
rect 17668 28924 18508 28980
rect 18564 28924 18574 28980
rect 19842 28924 19852 28980
rect 19908 28924 20636 28980
rect 20692 28924 21532 28980
rect 21588 28924 22092 28980
rect 22148 28924 22158 28980
rect 29922 28924 29932 28980
rect 29988 28924 34748 28980
rect 34804 28924 36428 28980
rect 36484 28924 38668 28980
rect 0 28896 800 28924
rect 38612 28868 38668 28924
rect 16594 28812 16604 28868
rect 16660 28812 17724 28868
rect 17780 28812 17790 28868
rect 18172 28812 22316 28868
rect 22372 28812 22382 28868
rect 28018 28812 28028 28868
rect 28084 28812 37100 28868
rect 37156 28812 37166 28868
rect 38612 28812 41132 28868
rect 41188 28812 41198 28868
rect 46386 28812 46396 28868
rect 46452 28812 47068 28868
rect 47124 28812 47134 28868
rect 48066 28812 48076 28868
rect 48132 28812 50204 28868
rect 50260 28812 50540 28868
rect 50596 28812 51548 28868
rect 51604 28812 51614 28868
rect 51874 28812 51884 28868
rect 51940 28812 52780 28868
rect 52836 28812 53340 28868
rect 53396 28812 53406 28868
rect 54114 28812 54124 28868
rect 54180 28812 55468 28868
rect 18172 28756 18228 28812
rect 55412 28756 55468 28812
rect 2370 28700 2380 28756
rect 2436 28700 6188 28756
rect 6244 28700 6254 28756
rect 6738 28700 6748 28756
rect 6804 28700 14028 28756
rect 14084 28700 14094 28756
rect 15026 28700 15036 28756
rect 15092 28700 18228 28756
rect 18386 28700 18396 28756
rect 18452 28700 19516 28756
rect 19572 28700 20300 28756
rect 20356 28700 22988 28756
rect 23044 28700 23054 28756
rect 25442 28700 25452 28756
rect 25508 28700 28140 28756
rect 28196 28700 29148 28756
rect 29204 28700 29214 28756
rect 32946 28700 32956 28756
rect 33012 28700 34300 28756
rect 34356 28700 34366 28756
rect 48290 28700 48300 28756
rect 48356 28700 49756 28756
rect 49812 28700 49822 28756
rect 55412 28700 55692 28756
rect 55748 28700 55758 28756
rect 4946 28588 4956 28644
rect 5012 28588 6076 28644
rect 6132 28588 6142 28644
rect 12450 28588 12460 28644
rect 12516 28588 13468 28644
rect 13524 28588 13534 28644
rect 13682 28588 13692 28644
rect 13748 28588 14700 28644
rect 14756 28588 15932 28644
rect 15988 28588 15998 28644
rect 16482 28588 16492 28644
rect 16548 28588 24108 28644
rect 24164 28588 24174 28644
rect 27234 28588 27244 28644
rect 27300 28588 28252 28644
rect 28308 28588 28318 28644
rect 33506 28588 33516 28644
rect 33572 28588 34524 28644
rect 34580 28588 34590 28644
rect 35970 28588 35980 28644
rect 36036 28588 37436 28644
rect 37492 28588 37502 28644
rect 41682 28588 41692 28644
rect 41748 28588 42588 28644
rect 42644 28588 43708 28644
rect 47730 28588 47740 28644
rect 47796 28588 48972 28644
rect 49028 28588 49038 28644
rect 43652 28532 43708 28588
rect 1922 28476 1932 28532
rect 1988 28476 3164 28532
rect 3220 28476 5740 28532
rect 5796 28476 5806 28532
rect 19170 28476 19180 28532
rect 19236 28476 24332 28532
rect 24388 28476 24398 28532
rect 27122 28476 27132 28532
rect 27188 28476 29260 28532
rect 29316 28476 29326 28532
rect 32050 28476 32060 28532
rect 32116 28476 32508 28532
rect 32564 28476 33292 28532
rect 33348 28476 33358 28532
rect 37986 28476 37996 28532
rect 38052 28476 39452 28532
rect 39508 28476 42028 28532
rect 42084 28476 42094 28532
rect 43652 28476 44716 28532
rect 44772 28476 45500 28532
rect 45556 28476 45566 28532
rect 49298 28476 49308 28532
rect 49364 28476 51884 28532
rect 51940 28476 51950 28532
rect 53218 28476 53228 28532
rect 53284 28476 54348 28532
rect 54404 28476 54684 28532
rect 54740 28476 54750 28532
rect 18946 28364 18956 28420
rect 19012 28364 25340 28420
rect 25396 28364 25406 28420
rect 25564 28364 27580 28420
rect 27636 28364 27646 28420
rect 36530 28364 36540 28420
rect 36596 28364 38668 28420
rect 38724 28364 38734 28420
rect 43250 28364 43260 28420
rect 43316 28364 45052 28420
rect 45108 28364 45118 28420
rect 0 28308 800 28336
rect 25564 28308 25620 28364
rect 0 28252 13916 28308
rect 13972 28252 13982 28308
rect 22306 28252 22316 28308
rect 22372 28252 25620 28308
rect 26002 28252 26012 28308
rect 26068 28252 27916 28308
rect 27972 28252 27982 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 27122 28140 27132 28196
rect 27188 28140 35532 28196
rect 35588 28140 35598 28196
rect 17938 28028 17948 28084
rect 18004 28028 19404 28084
rect 19460 28028 19470 28084
rect 24882 28028 24892 28084
rect 24948 28028 25340 28084
rect 25396 28028 25406 28084
rect 35634 28028 35644 28084
rect 35700 28028 37884 28084
rect 37940 28028 37950 28084
rect 25554 27916 25564 27972
rect 25620 27916 26908 27972
rect 26964 27916 28476 27972
rect 28532 27916 28542 27972
rect 41020 27916 41692 27972
rect 41748 27916 41758 27972
rect 42130 27916 42140 27972
rect 42196 27916 42364 27972
rect 42420 27916 43260 27972
rect 43316 27916 43326 27972
rect 45154 27916 45164 27972
rect 45220 27916 46060 27972
rect 46116 27916 46508 27972
rect 46564 27916 46574 27972
rect 50642 27916 50652 27972
rect 50708 27916 51660 27972
rect 51716 27916 51726 27972
rect 52098 27916 52108 27972
rect 52164 27916 53116 27972
rect 53172 27916 54572 27972
rect 54628 27916 55356 27972
rect 55412 27916 55422 27972
rect 41020 27860 41076 27916
rect 16034 27804 16044 27860
rect 16100 27804 18956 27860
rect 19012 27804 19022 27860
rect 25890 27804 25900 27860
rect 25956 27804 25966 27860
rect 26226 27804 26236 27860
rect 26292 27804 27020 27860
rect 27076 27804 27086 27860
rect 28130 27804 28140 27860
rect 28196 27804 28812 27860
rect 28868 27804 28878 27860
rect 31490 27804 31500 27860
rect 31556 27804 32396 27860
rect 32452 27804 32462 27860
rect 33394 27804 33404 27860
rect 33460 27804 35644 27860
rect 35700 27804 36316 27860
rect 36372 27804 36382 27860
rect 38658 27804 38668 27860
rect 38724 27804 40012 27860
rect 40068 27804 41020 27860
rect 41076 27804 41086 27860
rect 41346 27804 41356 27860
rect 41412 27804 42812 27860
rect 42868 27804 43596 27860
rect 43652 27804 43662 27860
rect 45602 27804 45612 27860
rect 45668 27804 46956 27860
rect 47012 27804 47022 27860
rect 51090 27804 51100 27860
rect 51156 27804 52332 27860
rect 52388 27804 54908 27860
rect 54964 27804 54974 27860
rect 24546 27692 24556 27748
rect 24612 27692 25676 27748
rect 25732 27692 25742 27748
rect 0 27636 800 27664
rect 25900 27636 25956 27804
rect 38882 27692 38892 27748
rect 38948 27692 39788 27748
rect 39844 27692 42028 27748
rect 42084 27692 42094 27748
rect 0 27580 6748 27636
rect 6804 27580 6814 27636
rect 25900 27580 27020 27636
rect 27076 27580 27086 27636
rect 29698 27580 29708 27636
rect 29764 27580 31836 27636
rect 31892 27580 31902 27636
rect 33730 27580 33740 27636
rect 33796 27580 34412 27636
rect 34468 27580 35980 27636
rect 36036 27580 36988 27636
rect 37044 27580 38444 27636
rect 38500 27580 40348 27636
rect 40404 27580 41356 27636
rect 41412 27580 41422 27636
rect 0 27552 800 27580
rect 24658 27468 24668 27524
rect 24724 27468 28140 27524
rect 28196 27468 28206 27524
rect 29250 27468 29260 27524
rect 29316 27468 48524 27524
rect 48580 27468 48590 27524
rect 19506 27356 19516 27412
rect 19572 27356 26236 27412
rect 26292 27356 26302 27412
rect 26758 27356 26796 27412
rect 26852 27356 26862 27412
rect 30146 27356 30156 27412
rect 30212 27356 33404 27412
rect 33460 27356 33470 27412
rect 35634 27356 35644 27412
rect 35700 27356 36540 27412
rect 36596 27356 36606 27412
rect 37762 27356 37772 27412
rect 37828 27356 38556 27412
rect 38612 27356 38622 27412
rect 23426 27244 23436 27300
rect 23492 27244 32732 27300
rect 32788 27244 32798 27300
rect 4466 27188 4476 27244
rect 4532 27188 4580 27244
rect 4636 27188 4684 27244
rect 4740 27188 4750 27244
rect 35186 27188 35196 27244
rect 35252 27188 35300 27244
rect 35356 27188 35404 27244
rect 35460 27188 35470 27244
rect 25778 27132 25788 27188
rect 25844 27132 26124 27188
rect 26180 27132 26190 27188
rect 26450 27020 26460 27076
rect 26516 27020 28700 27076
rect 28756 27020 28766 27076
rect 32386 27020 32396 27076
rect 32452 27020 33292 27076
rect 33348 27020 33358 27076
rect 0 26964 800 26992
rect 0 26908 15036 26964
rect 15092 26908 15102 26964
rect 26114 26908 26124 26964
rect 26180 26908 26796 26964
rect 26852 26908 26862 26964
rect 31602 26908 31612 26964
rect 31668 26908 32508 26964
rect 32564 26908 32574 26964
rect 35252 26908 40404 26964
rect 0 26880 800 26908
rect 35252 26852 35308 26908
rect 40348 26852 40404 26908
rect 2706 26796 2716 26852
rect 2772 26796 4956 26852
rect 5012 26796 5022 26852
rect 8306 26796 8316 26852
rect 8372 26796 9324 26852
rect 9380 26796 10108 26852
rect 10164 26796 11228 26852
rect 11284 26796 11294 26852
rect 12786 26796 12796 26852
rect 12852 26796 13468 26852
rect 13524 26796 13534 26852
rect 25666 26796 25676 26852
rect 25732 26796 27356 26852
rect 27412 26796 27422 26852
rect 28476 26796 35308 26852
rect 37202 26796 37212 26852
rect 37268 26796 39116 26852
rect 39172 26796 40012 26852
rect 40068 26796 40078 26852
rect 40348 26796 44716 26852
rect 44772 26796 44782 26852
rect 48178 26796 48188 26852
rect 48244 26796 51548 26852
rect 51604 26796 51614 26852
rect 28476 26740 28532 26796
rect 12898 26684 12908 26740
rect 12964 26684 14028 26740
rect 14084 26684 14094 26740
rect 14242 26684 14252 26740
rect 14308 26684 16156 26740
rect 16212 26684 16222 26740
rect 28466 26684 28476 26740
rect 28532 26684 28542 26740
rect 30034 26684 30044 26740
rect 30100 26684 31948 26740
rect 33058 26684 33068 26740
rect 33124 26684 33740 26740
rect 33796 26684 33806 26740
rect 37090 26684 37100 26740
rect 37156 26684 38780 26740
rect 38836 26684 38846 26740
rect 39890 26684 39900 26740
rect 39956 26684 40572 26740
rect 40628 26684 40638 26740
rect 44258 26684 44268 26740
rect 44324 26684 45500 26740
rect 45556 26684 45566 26740
rect 49746 26684 49756 26740
rect 49812 26684 50428 26740
rect 50484 26684 50988 26740
rect 51044 26684 51054 26740
rect 51314 26684 51324 26740
rect 51380 26684 53676 26740
rect 53732 26684 53742 26740
rect 31892 26628 31948 26684
rect 39900 26628 39956 26684
rect 9762 26572 9772 26628
rect 9828 26572 11452 26628
rect 11508 26572 14476 26628
rect 14532 26572 14542 26628
rect 22194 26572 22204 26628
rect 22260 26572 24108 26628
rect 24164 26572 24174 26628
rect 27346 26572 27356 26628
rect 27412 26572 31388 26628
rect 31444 26572 31454 26628
rect 31892 26572 34188 26628
rect 34244 26572 34748 26628
rect 34804 26572 39956 26628
rect 40338 26572 40348 26628
rect 40404 26572 40684 26628
rect 40740 26572 42140 26628
rect 42196 26572 42924 26628
rect 42980 26572 42990 26628
rect 45602 26572 45612 26628
rect 45668 26572 50876 26628
rect 50932 26572 50942 26628
rect 51202 26572 51212 26628
rect 51268 26572 52108 26628
rect 52164 26572 53452 26628
rect 53508 26572 53518 26628
rect 13570 26460 13580 26516
rect 13636 26460 15484 26516
rect 15540 26460 16604 26516
rect 16660 26460 16670 26516
rect 26338 26460 26348 26516
rect 26404 26460 26796 26516
rect 26852 26460 27468 26516
rect 27524 26460 27534 26516
rect 28242 26460 28252 26516
rect 28308 26460 28812 26516
rect 28868 26460 28878 26516
rect 30034 26460 30044 26516
rect 30100 26460 31612 26516
rect 31668 26460 31678 26516
rect 32498 26460 32508 26516
rect 32564 26460 37548 26516
rect 37604 26460 37614 26516
rect 38434 26460 38444 26516
rect 38500 26460 39004 26516
rect 39060 26460 39564 26516
rect 39620 26460 47852 26516
rect 47908 26460 48636 26516
rect 48692 26460 48702 26516
rect 10994 26348 11004 26404
rect 11060 26348 12796 26404
rect 12852 26348 14364 26404
rect 14420 26348 14430 26404
rect 28914 26348 28924 26404
rect 28980 26348 29596 26404
rect 29652 26348 30940 26404
rect 30996 26348 31006 26404
rect 36530 26348 36540 26404
rect 36596 26348 38332 26404
rect 38388 26348 38398 26404
rect 38882 26348 38892 26404
rect 38948 26348 41244 26404
rect 41300 26348 41310 26404
rect 30482 26236 30492 26292
rect 30548 26236 31276 26292
rect 31332 26236 31612 26292
rect 31668 26236 31678 26292
rect 19826 26180 19836 26236
rect 19892 26180 19940 26236
rect 19996 26180 20044 26236
rect 20100 26180 20110 26236
rect 30492 26180 30548 26236
rect 50546 26180 50556 26236
rect 50612 26180 50660 26236
rect 50716 26180 50764 26236
rect 50820 26180 50830 26236
rect 21858 26124 21868 26180
rect 21924 26124 23324 26180
rect 23380 26124 25564 26180
rect 25620 26124 27020 26180
rect 27076 26124 30548 26180
rect 35970 26012 35980 26068
rect 36036 26012 36764 26068
rect 36820 26012 37772 26068
rect 37828 26012 37838 26068
rect 37986 26012 37996 26068
rect 38052 26012 39228 26068
rect 39284 26012 39294 26068
rect 1810 25900 1820 25956
rect 1876 25900 2716 25956
rect 2772 25900 2782 25956
rect 30706 25900 30716 25956
rect 30772 25900 38668 25956
rect 38724 25900 39116 25956
rect 39172 25900 39182 25956
rect 40002 25900 40012 25956
rect 40068 25900 42140 25956
rect 42196 25900 42206 25956
rect 53890 25900 53900 25956
rect 53956 25900 54908 25956
rect 54964 25900 55356 25956
rect 55412 25900 56700 25956
rect 56756 25900 56766 25956
rect 35522 25788 35532 25844
rect 35588 25788 35644 25844
rect 35700 25788 38332 25844
rect 38388 25788 38398 25844
rect 43810 25788 43820 25844
rect 43876 25788 45612 25844
rect 45668 25788 45678 25844
rect 47618 25788 47628 25844
rect 47684 25788 49644 25844
rect 49700 25788 49710 25844
rect 5730 25676 5740 25732
rect 5796 25676 7196 25732
rect 7252 25676 7262 25732
rect 8372 25676 8764 25732
rect 8820 25676 8830 25732
rect 19954 25676 19964 25732
rect 20020 25676 21420 25732
rect 21476 25676 21486 25732
rect 27794 25676 27804 25732
rect 27860 25676 28476 25732
rect 28532 25676 31164 25732
rect 31220 25676 32172 25732
rect 32228 25676 32238 25732
rect 42018 25676 42028 25732
rect 42084 25676 42476 25732
rect 42532 25676 42542 25732
rect 44370 25676 44380 25732
rect 44436 25676 46060 25732
rect 46116 25676 46126 25732
rect 48066 25676 48076 25732
rect 48132 25676 49084 25732
rect 49140 25676 49150 25732
rect 50194 25676 50204 25732
rect 50260 25676 52220 25732
rect 52276 25676 54460 25732
rect 54516 25676 54526 25732
rect 8372 25620 8428 25676
rect 2258 25564 2268 25620
rect 2324 25564 3948 25620
rect 4004 25564 4014 25620
rect 6178 25564 6188 25620
rect 6244 25564 8428 25620
rect 16818 25564 16828 25620
rect 16884 25564 17836 25620
rect 17892 25564 17902 25620
rect 22754 25564 22764 25620
rect 22820 25564 27468 25620
rect 27524 25564 30380 25620
rect 30436 25564 30446 25620
rect 26226 25452 26236 25508
rect 26292 25452 26908 25508
rect 26964 25452 26974 25508
rect 31826 25452 31836 25508
rect 31892 25452 33628 25508
rect 33684 25452 43820 25508
rect 43876 25452 43886 25508
rect 1810 25340 1820 25396
rect 1876 25340 3500 25396
rect 3556 25340 3566 25396
rect 9650 25340 9660 25396
rect 9716 25340 11340 25396
rect 11396 25340 12124 25396
rect 12180 25340 12190 25396
rect 21410 25340 21420 25396
rect 21476 25340 21868 25396
rect 21924 25340 21934 25396
rect 24770 25340 24780 25396
rect 24836 25340 25564 25396
rect 25620 25340 25630 25396
rect 28578 25340 28588 25396
rect 28644 25340 29372 25396
rect 29428 25340 29438 25396
rect 33842 25340 33852 25396
rect 33908 25340 34860 25396
rect 34916 25340 37548 25396
rect 37604 25340 37614 25396
rect 5842 25228 5852 25284
rect 5908 25228 8204 25284
rect 8260 25228 8270 25284
rect 20514 25228 20524 25284
rect 20580 25228 23324 25284
rect 23380 25228 23390 25284
rect 24556 25228 25452 25284
rect 25508 25228 25518 25284
rect 35532 25228 36988 25284
rect 37044 25228 37054 25284
rect 4466 25172 4476 25228
rect 4532 25172 4580 25228
rect 4636 25172 4684 25228
rect 4740 25172 4750 25228
rect 24556 25172 24612 25228
rect 35186 25172 35196 25228
rect 35252 25172 35300 25228
rect 35356 25172 35404 25228
rect 35460 25172 35470 25228
rect 24546 25116 24556 25172
rect 24612 25116 24622 25172
rect 28130 25116 28140 25172
rect 28196 25116 31052 25172
rect 31108 25116 31118 25172
rect 35532 25060 35588 25228
rect 39554 25116 39564 25172
rect 39620 25116 40572 25172
rect 40628 25116 40638 25172
rect 51650 25116 51660 25172
rect 51716 25116 52892 25172
rect 52948 25116 54908 25172
rect 54964 25116 55804 25172
rect 55860 25116 55870 25172
rect 31378 25004 31388 25060
rect 31444 25004 32508 25060
rect 32564 25004 32574 25060
rect 34514 25004 34524 25060
rect 34580 25004 35196 25060
rect 35252 25004 35588 25060
rect 21410 24892 21420 24948
rect 21476 24892 21980 24948
rect 22036 24892 22046 24948
rect 22978 24892 22988 24948
rect 23044 24892 30268 24948
rect 30324 24892 30334 24948
rect 36194 24892 36204 24948
rect 36260 24892 36764 24948
rect 36820 24892 36830 24948
rect 17602 24780 17612 24836
rect 17668 24780 19404 24836
rect 19460 24780 19964 24836
rect 20020 24780 20030 24836
rect 25554 24780 25564 24836
rect 25620 24780 27020 24836
rect 27076 24780 27086 24836
rect 28252 24780 30044 24836
rect 30100 24780 31948 24836
rect 32004 24780 32014 24836
rect 33954 24780 33964 24836
rect 34020 24780 35644 24836
rect 35700 24780 36540 24836
rect 36596 24780 36606 24836
rect 45266 24780 45276 24836
rect 45332 24780 45724 24836
rect 45780 24780 46396 24836
rect 46452 24780 46462 24836
rect 28252 24724 28308 24780
rect 4834 24668 4844 24724
rect 4900 24668 5628 24724
rect 5684 24668 5694 24724
rect 9314 24668 9324 24724
rect 9380 24668 10220 24724
rect 10276 24668 10892 24724
rect 10948 24668 10958 24724
rect 16258 24668 16268 24724
rect 16324 24668 17500 24724
rect 17556 24668 17566 24724
rect 17938 24668 17948 24724
rect 18004 24668 19068 24724
rect 19124 24668 19134 24724
rect 21970 24668 21980 24724
rect 22036 24668 28252 24724
rect 28308 24668 28318 24724
rect 29810 24668 29820 24724
rect 29876 24668 29886 24724
rect 32610 24668 32620 24724
rect 32676 24668 35644 24724
rect 35700 24668 35710 24724
rect 24882 24556 24892 24612
rect 24948 24556 27244 24612
rect 27300 24556 28140 24612
rect 28196 24556 28206 24612
rect 29820 24500 29876 24668
rect 36540 24500 36596 24780
rect 51874 24668 51884 24724
rect 51940 24668 53452 24724
rect 53508 24668 53518 24724
rect 56690 24668 56700 24724
rect 56756 24668 57932 24724
rect 57988 24668 57998 24724
rect 5058 24444 5068 24500
rect 5124 24444 6188 24500
rect 6244 24444 6524 24500
rect 6580 24444 6590 24500
rect 9538 24444 9548 24500
rect 9604 24444 12348 24500
rect 12404 24444 14028 24500
rect 14084 24444 14588 24500
rect 14644 24444 14654 24500
rect 22306 24444 22316 24500
rect 22372 24444 23548 24500
rect 23604 24444 23614 24500
rect 24098 24444 24108 24500
rect 24164 24444 25004 24500
rect 25060 24444 25070 24500
rect 25442 24444 25452 24500
rect 25508 24444 26124 24500
rect 26180 24444 26572 24500
rect 26628 24444 26638 24500
rect 28354 24444 28364 24500
rect 28420 24444 29260 24500
rect 29316 24444 29326 24500
rect 29820 24444 34524 24500
rect 34580 24444 35420 24500
rect 35476 24444 35486 24500
rect 36540 24444 40124 24500
rect 40180 24444 40796 24500
rect 40852 24444 41468 24500
rect 41524 24444 42140 24500
rect 42196 24444 43708 24500
rect 51874 24444 51884 24500
rect 51940 24444 52892 24500
rect 52948 24444 52958 24500
rect 37202 24332 37212 24388
rect 37268 24332 38108 24388
rect 38164 24332 38174 24388
rect 43652 24276 43708 24444
rect 55682 24332 55692 24388
rect 55748 24332 57484 24388
rect 57540 24332 57550 24388
rect 40226 24220 40236 24276
rect 40292 24220 41692 24276
rect 41748 24220 41758 24276
rect 43652 24220 44324 24276
rect 19826 24164 19836 24220
rect 19892 24164 19940 24220
rect 19996 24164 20044 24220
rect 20100 24164 20110 24220
rect 26338 24108 26348 24164
rect 26404 24108 35868 24164
rect 35924 24108 36764 24164
rect 36820 24108 36830 24164
rect 40450 24108 40460 24164
rect 40516 24108 41580 24164
rect 41636 24108 42364 24164
rect 42420 24108 43708 24164
rect 43652 23940 43708 24108
rect 44268 24052 44324 24220
rect 50546 24164 50556 24220
rect 50612 24164 50660 24220
rect 50716 24164 50764 24220
rect 50820 24164 50830 24220
rect 44258 23996 44268 24052
rect 44324 23996 46060 24052
rect 46116 23996 49980 24052
rect 50036 23996 50428 24052
rect 50484 23996 50494 24052
rect 1810 23884 1820 23940
rect 1876 23884 2604 23940
rect 2660 23884 2670 23940
rect 19058 23884 19068 23940
rect 19124 23884 22092 23940
rect 22148 23884 22158 23940
rect 23202 23884 23212 23940
rect 23268 23884 24556 23940
rect 24612 23884 24622 23940
rect 25890 23884 25900 23940
rect 25956 23884 26684 23940
rect 26740 23884 26750 23940
rect 39330 23884 39340 23940
rect 39396 23884 41244 23940
rect 41300 23884 41916 23940
rect 41972 23884 42476 23940
rect 42532 23884 42542 23940
rect 43652 23884 44380 23940
rect 44436 23884 44446 23940
rect 45602 23884 45612 23940
rect 45668 23884 53900 23940
rect 53956 23884 53966 23940
rect 54114 23884 54124 23940
rect 54180 23884 57148 23940
rect 57204 23884 57820 23940
rect 57876 23884 57886 23940
rect 44380 23828 44436 23884
rect 24770 23772 24780 23828
rect 24836 23772 26348 23828
rect 26404 23772 27580 23828
rect 27636 23772 27646 23828
rect 28690 23772 28700 23828
rect 28756 23772 30940 23828
rect 30996 23772 31612 23828
rect 31668 23772 32956 23828
rect 33012 23772 33022 23828
rect 44380 23772 45724 23828
rect 45780 23772 48860 23828
rect 48916 23772 49420 23828
rect 49476 23772 51772 23828
rect 51828 23772 51838 23828
rect 17490 23660 17500 23716
rect 17556 23660 18844 23716
rect 18900 23660 20300 23716
rect 20356 23660 20366 23716
rect 25106 23660 25116 23716
rect 25172 23660 25452 23716
rect 25508 23660 25518 23716
rect 28242 23660 28252 23716
rect 28308 23660 29036 23716
rect 29092 23660 29102 23716
rect 31892 23660 33292 23716
rect 33348 23660 33740 23716
rect 33796 23660 35196 23716
rect 35252 23660 35262 23716
rect 36194 23660 36204 23716
rect 36260 23660 37884 23716
rect 37940 23660 37950 23716
rect 49522 23660 49532 23716
rect 49588 23660 50204 23716
rect 50260 23660 50652 23716
rect 50708 23660 50718 23716
rect 31892 23604 31948 23660
rect 1922 23548 1932 23604
rect 1988 23548 3164 23604
rect 3220 23548 4844 23604
rect 4900 23548 4910 23604
rect 16818 23548 16828 23604
rect 16884 23548 18396 23604
rect 18452 23548 18462 23604
rect 22530 23548 22540 23604
rect 22596 23548 23436 23604
rect 23492 23548 24108 23604
rect 24164 23548 25788 23604
rect 25844 23548 26348 23604
rect 26404 23548 27804 23604
rect 27860 23548 28924 23604
rect 28980 23548 31948 23604
rect 32050 23548 32060 23604
rect 32116 23548 32620 23604
rect 32676 23548 34076 23604
rect 34132 23548 34142 23604
rect 56690 23548 56700 23604
rect 56756 23548 57596 23604
rect 57652 23548 57662 23604
rect 23874 23436 23884 23492
rect 23940 23436 24892 23492
rect 24948 23436 40348 23492
rect 40404 23436 40414 23492
rect 4466 23156 4476 23212
rect 4532 23156 4580 23212
rect 4636 23156 4684 23212
rect 4740 23156 4750 23212
rect 35186 23156 35196 23212
rect 35252 23156 35300 23212
rect 35356 23156 35404 23212
rect 35460 23156 35470 23212
rect 35746 22876 35756 22932
rect 35812 22876 36988 22932
rect 37044 22876 37054 22932
rect 4610 22764 4620 22820
rect 4676 22764 5740 22820
rect 5796 22764 5806 22820
rect 34402 22764 34412 22820
rect 34468 22764 37548 22820
rect 37604 22764 38220 22820
rect 38276 22764 38286 22820
rect 41010 22764 41020 22820
rect 41076 22764 41916 22820
rect 41972 22764 43036 22820
rect 43092 22764 43484 22820
rect 43540 22764 43550 22820
rect 21746 22652 21756 22708
rect 21812 22652 23884 22708
rect 23940 22652 23950 22708
rect 18386 22540 18396 22596
rect 18452 22540 20188 22596
rect 20244 22540 20636 22596
rect 20692 22540 20702 22596
rect 25218 22540 25228 22596
rect 25284 22540 25676 22596
rect 25732 22540 25742 22596
rect 35074 22540 35084 22596
rect 35140 22540 36092 22596
rect 36148 22540 36158 22596
rect 43484 22484 43540 22764
rect 31266 22428 31276 22484
rect 31332 22428 32508 22484
rect 32564 22428 33292 22484
rect 33348 22428 33358 22484
rect 43484 22428 44940 22484
rect 44996 22428 45006 22484
rect 55010 22428 55020 22484
rect 55076 22428 56476 22484
rect 56532 22428 56542 22484
rect 15250 22316 15260 22372
rect 15316 22316 26124 22372
rect 26180 22316 26190 22372
rect 19826 22148 19836 22204
rect 19892 22148 19940 22204
rect 19996 22148 20044 22204
rect 20100 22148 20110 22204
rect 50546 22148 50556 22204
rect 50612 22148 50660 22204
rect 50716 22148 50764 22204
rect 50820 22148 50830 22204
rect 16930 21868 16940 21924
rect 16996 21868 17948 21924
rect 18004 21868 18284 21924
rect 18340 21868 18350 21924
rect 33618 21868 33628 21924
rect 33684 21868 34748 21924
rect 34804 21868 35532 21924
rect 35588 21868 37940 21924
rect 37884 21812 37940 21868
rect 18610 21756 18620 21812
rect 18676 21756 19180 21812
rect 19236 21756 19246 21812
rect 37874 21756 37884 21812
rect 37940 21756 38220 21812
rect 38276 21756 39900 21812
rect 39956 21756 40460 21812
rect 40516 21756 41132 21812
rect 41188 21756 41198 21812
rect 49746 21756 49756 21812
rect 49812 21756 50764 21812
rect 50820 21756 51436 21812
rect 51492 21756 51502 21812
rect 51986 21756 51996 21812
rect 52052 21756 53564 21812
rect 53620 21756 53630 21812
rect 56690 21756 56700 21812
rect 56756 21756 57708 21812
rect 57764 21756 57774 21812
rect 20738 21644 20748 21700
rect 20804 21644 21196 21700
rect 21252 21644 22764 21700
rect 22820 21644 22830 21700
rect 24546 21644 24556 21700
rect 24612 21644 25564 21700
rect 25620 21644 25630 21700
rect 35634 21644 35644 21700
rect 35700 21644 36204 21700
rect 36260 21644 37100 21700
rect 37156 21644 37166 21700
rect 41234 21644 41244 21700
rect 41300 21644 43036 21700
rect 43092 21644 43102 21700
rect 46498 21644 46508 21700
rect 46564 21644 47740 21700
rect 47796 21644 48412 21700
rect 48468 21644 50204 21700
rect 50260 21644 50270 21700
rect 24210 21532 24220 21588
rect 24276 21532 26124 21588
rect 26180 21532 26190 21588
rect 28924 21532 30380 21588
rect 30436 21532 31388 21588
rect 31444 21532 31454 21588
rect 33170 21532 33180 21588
rect 33236 21532 34860 21588
rect 34916 21532 34926 21588
rect 41682 21532 41692 21588
rect 41748 21532 42252 21588
rect 42308 21532 42318 21588
rect 50642 21532 50652 21588
rect 50708 21532 51996 21588
rect 52052 21532 52062 21588
rect 28924 21476 28980 21532
rect 17938 21420 17948 21476
rect 18004 21420 26236 21476
rect 26292 21420 26796 21476
rect 26852 21420 28924 21476
rect 28980 21420 28990 21476
rect 29362 21420 29372 21476
rect 29428 21420 41468 21476
rect 41524 21420 41534 21476
rect 41570 21308 41580 21364
rect 41636 21308 42700 21364
rect 42756 21308 47404 21364
rect 47460 21308 48188 21364
rect 48244 21308 48254 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 41794 20972 41804 21028
rect 41860 20972 43036 21028
rect 43092 20972 43102 21028
rect 54786 20972 54796 21028
rect 54852 20972 56476 21028
rect 56532 20972 56542 21028
rect 38770 20860 38780 20916
rect 38836 20860 40124 20916
rect 40180 20860 40684 20916
rect 40740 20860 43372 20916
rect 43428 20860 43438 20916
rect 16258 20748 16268 20804
rect 16324 20748 16940 20804
rect 16996 20748 17006 20804
rect 19842 20748 19852 20804
rect 19908 20748 20188 20804
rect 46722 20748 46732 20804
rect 46788 20748 47628 20804
rect 47684 20748 48412 20804
rect 48468 20748 48478 20804
rect 20132 20692 20188 20748
rect 20132 20636 21420 20692
rect 21476 20636 22540 20692
rect 22596 20636 23212 20692
rect 23268 20636 23278 20692
rect 23650 20636 23660 20692
rect 23716 20636 24780 20692
rect 24836 20636 24846 20692
rect 31892 20636 36428 20692
rect 36484 20636 38556 20692
rect 38612 20636 38622 20692
rect 45042 20636 45052 20692
rect 45108 20636 46172 20692
rect 46228 20636 48076 20692
rect 48132 20636 49308 20692
rect 49364 20636 50092 20692
rect 50148 20636 50764 20692
rect 50820 20636 50830 20692
rect 55906 20636 55916 20692
rect 55972 20636 56812 20692
rect 56868 20636 56878 20692
rect 20290 20524 20300 20580
rect 20356 20524 21644 20580
rect 21700 20524 24220 20580
rect 24276 20524 24286 20580
rect 19170 20412 19180 20468
rect 19236 20412 20188 20468
rect 20244 20412 20748 20468
rect 20804 20412 20814 20468
rect 27458 20300 27468 20356
rect 27524 20300 28476 20356
rect 28532 20300 30156 20356
rect 30212 20300 30222 20356
rect 31892 20244 31948 20636
rect 55916 20580 55972 20636
rect 37090 20524 37100 20580
rect 37156 20524 37660 20580
rect 37716 20524 40012 20580
rect 40068 20524 41580 20580
rect 41636 20524 41646 20580
rect 51986 20524 51996 20580
rect 52052 20524 53564 20580
rect 53620 20524 54908 20580
rect 54964 20524 55468 20580
rect 55524 20524 55972 20580
rect 42802 20412 42812 20468
rect 42868 20412 43708 20468
rect 43764 20412 43774 20468
rect 54114 20412 54124 20468
rect 54180 20412 55692 20468
rect 55748 20412 56700 20468
rect 56756 20412 56766 20468
rect 14690 20188 14700 20244
rect 14756 20188 15260 20244
rect 15316 20188 16828 20244
rect 16884 20188 16894 20244
rect 25554 20188 25564 20244
rect 25620 20188 29708 20244
rect 29764 20188 31948 20244
rect 19826 20132 19836 20188
rect 19892 20132 19940 20188
rect 19996 20132 20044 20188
rect 20100 20132 20110 20188
rect 36306 20132 36316 20188
rect 36372 20132 36382 20188
rect 50546 20132 50556 20188
rect 50612 20132 50660 20188
rect 50716 20132 50764 20188
rect 50820 20132 50830 20188
rect 25330 20076 25340 20132
rect 25396 20076 25900 20132
rect 25956 20076 26460 20132
rect 26516 20076 27468 20132
rect 27524 20076 27534 20132
rect 30258 20076 30268 20132
rect 30324 20076 31724 20132
rect 31780 20076 32060 20132
rect 32116 20076 32126 20132
rect 36316 20076 37660 20132
rect 37716 20076 37726 20132
rect 36316 20020 36372 20076
rect 22530 19964 22540 20020
rect 22596 19964 26236 20020
rect 26292 19964 26302 20020
rect 33170 19964 33180 20020
rect 33236 19964 34188 20020
rect 34244 19964 35868 20020
rect 35924 19964 36372 20020
rect 36642 19964 36652 20020
rect 36708 19964 37772 20020
rect 37828 19964 38668 20020
rect 38724 19964 38734 20020
rect 52770 19964 52780 20020
rect 52836 19964 54796 20020
rect 54852 19964 54862 20020
rect 16706 19852 16716 19908
rect 16772 19852 18172 19908
rect 18228 19852 18238 19908
rect 33394 19852 33404 19908
rect 33460 19852 34524 19908
rect 34580 19852 34590 19908
rect 48514 19852 48524 19908
rect 48580 19852 49756 19908
rect 49812 19852 49822 19908
rect 19618 19740 19628 19796
rect 19684 19740 20300 19796
rect 20356 19740 20366 19796
rect 34178 19740 34188 19796
rect 34244 19740 39452 19796
rect 39508 19740 39518 19796
rect 48290 19740 48300 19796
rect 48356 19740 50204 19796
rect 50260 19740 50270 19796
rect 51650 19740 51660 19796
rect 51716 19740 53340 19796
rect 53396 19740 54572 19796
rect 54628 19740 55132 19796
rect 55188 19740 55198 19796
rect 19282 19628 19292 19684
rect 19348 19628 20188 19684
rect 20244 19628 20254 19684
rect 24322 19628 24332 19684
rect 24388 19628 26236 19684
rect 26292 19628 26302 19684
rect 31714 19628 31724 19684
rect 31780 19628 31948 19684
rect 36082 19628 36092 19684
rect 36148 19628 37100 19684
rect 37156 19628 37166 19684
rect 39218 19628 39228 19684
rect 39284 19628 41020 19684
rect 41076 19628 41086 19684
rect 41346 19628 41356 19684
rect 41412 19628 41804 19684
rect 41860 19628 41870 19684
rect 47954 19628 47964 19684
rect 48020 19628 48748 19684
rect 48804 19628 48814 19684
rect 31892 19572 31948 19628
rect 22082 19516 22092 19572
rect 22148 19516 22764 19572
rect 22820 19516 25564 19572
rect 25620 19516 25630 19572
rect 31892 19516 32172 19572
rect 32228 19516 32238 19572
rect 18610 19292 18620 19348
rect 18676 19292 24892 19348
rect 24948 19292 24958 19348
rect 4466 19124 4476 19180
rect 4532 19124 4580 19180
rect 4636 19124 4684 19180
rect 4740 19124 4750 19180
rect 35186 19124 35196 19180
rect 35252 19124 35300 19180
rect 35356 19124 35404 19180
rect 35460 19124 35470 19180
rect 27122 18732 27132 18788
rect 27188 18732 30156 18788
rect 30212 18732 30222 18788
rect 33618 18732 33628 18788
rect 33684 18732 34524 18788
rect 34580 18732 36204 18788
rect 36260 18732 36652 18788
rect 36708 18732 36718 18788
rect 37762 18732 37772 18788
rect 37828 18732 39116 18788
rect 39172 18732 39182 18788
rect 31042 18620 31052 18676
rect 31108 18620 32508 18676
rect 32564 18620 34972 18676
rect 35028 18620 35038 18676
rect 36316 18620 38780 18676
rect 38836 18620 38846 18676
rect 51874 18620 51884 18676
rect 51940 18620 52668 18676
rect 52724 18620 54348 18676
rect 54404 18620 54684 18676
rect 54740 18620 54750 18676
rect 36316 18564 36372 18620
rect 26002 18508 26012 18564
rect 26068 18508 28588 18564
rect 28644 18508 30044 18564
rect 30100 18508 31500 18564
rect 31556 18508 34076 18564
rect 34132 18508 34748 18564
rect 34804 18508 36316 18564
rect 36372 18508 36382 18564
rect 38658 18508 38668 18564
rect 38724 18508 40124 18564
rect 40180 18508 41020 18564
rect 41076 18508 41244 18564
rect 41300 18508 41310 18564
rect 43474 18508 43484 18564
rect 43540 18508 46172 18564
rect 46228 18508 46238 18564
rect 50530 18508 50540 18564
rect 50596 18508 51996 18564
rect 52052 18508 52892 18564
rect 52948 18508 52958 18564
rect 53218 18508 53228 18564
rect 53284 18508 54124 18564
rect 54180 18508 54190 18564
rect 56914 18508 56924 18564
rect 56980 18508 57708 18564
rect 57764 18508 57774 18564
rect 39778 18396 39788 18452
rect 39844 18396 41132 18452
rect 41188 18396 41198 18452
rect 19826 18116 19836 18172
rect 19892 18116 19940 18172
rect 19996 18116 20044 18172
rect 20100 18116 20110 18172
rect 50546 18116 50556 18172
rect 50612 18116 50660 18172
rect 50716 18116 50764 18172
rect 50820 18116 50830 18172
rect 42242 17948 42252 18004
rect 42308 17948 43708 18004
rect 43652 17892 43708 17948
rect 26786 17836 26796 17892
rect 26852 17836 27804 17892
rect 27860 17836 27870 17892
rect 28354 17836 28364 17892
rect 28420 17836 34636 17892
rect 34692 17836 34702 17892
rect 38770 17836 38780 17892
rect 38836 17836 39452 17892
rect 39508 17836 39900 17892
rect 39956 17836 39966 17892
rect 41458 17836 41468 17892
rect 41524 17836 42140 17892
rect 42196 17836 43260 17892
rect 43316 17836 43326 17892
rect 43652 17836 44492 17892
rect 44548 17836 44558 17892
rect 51538 17836 51548 17892
rect 51604 17836 53676 17892
rect 53732 17836 53742 17892
rect 39900 17780 39956 17836
rect 28466 17724 28476 17780
rect 28532 17724 29596 17780
rect 29652 17724 29662 17780
rect 39900 17724 41244 17780
rect 41300 17724 42252 17780
rect 42308 17724 42318 17780
rect 32162 17612 32172 17668
rect 32228 17612 34188 17668
rect 34244 17612 34254 17668
rect 41682 17612 41692 17668
rect 41748 17612 42700 17668
rect 42756 17612 42766 17668
rect 43652 17556 43708 17780
rect 43764 17724 43774 17780
rect 50866 17612 50876 17668
rect 50932 17612 53452 17668
rect 53508 17612 53518 17668
rect 32498 17500 32508 17556
rect 32564 17500 33516 17556
rect 33572 17500 35644 17556
rect 35700 17500 36764 17556
rect 36820 17500 39788 17556
rect 39844 17500 39854 17556
rect 40338 17500 40348 17556
rect 40404 17500 40908 17556
rect 40964 17500 41916 17556
rect 41972 17500 43708 17556
rect 45602 17500 45612 17556
rect 45668 17500 47180 17556
rect 47236 17500 48972 17556
rect 49028 17500 49532 17556
rect 49588 17500 49598 17556
rect 34738 17276 34748 17332
rect 34804 17276 36764 17332
rect 36820 17276 36830 17332
rect 4466 17108 4476 17164
rect 4532 17108 4580 17164
rect 4636 17108 4684 17164
rect 4740 17108 4750 17164
rect 35186 17108 35196 17164
rect 35252 17108 35300 17164
rect 35356 17108 35404 17164
rect 35460 17108 35470 17164
rect 18722 16828 18732 16884
rect 18788 16828 19516 16884
rect 19572 16828 23268 16884
rect 23212 16772 23268 16828
rect 21858 16716 21868 16772
rect 21924 16716 22988 16772
rect 23044 16716 23054 16772
rect 23202 16716 23212 16772
rect 23268 16716 23660 16772
rect 23716 16716 24220 16772
rect 24276 16716 26012 16772
rect 26068 16716 26078 16772
rect 31490 16716 31500 16772
rect 31556 16716 31948 16772
rect 32004 16716 32014 16772
rect 22082 16604 22092 16660
rect 22148 16604 24108 16660
rect 24164 16604 24444 16660
rect 24500 16604 24510 16660
rect 24770 16604 24780 16660
rect 24836 16604 26796 16660
rect 26852 16604 26862 16660
rect 39218 16604 39228 16660
rect 39284 16604 39900 16660
rect 39956 16604 45052 16660
rect 45108 16604 45118 16660
rect 45714 16604 45724 16660
rect 45780 16604 47404 16660
rect 47460 16604 47470 16660
rect 54562 16604 54572 16660
rect 54628 16604 55020 16660
rect 55076 16604 55580 16660
rect 55636 16604 56140 16660
rect 56196 16604 56206 16660
rect 24780 16548 24836 16604
rect 22530 16492 22540 16548
rect 22596 16492 23436 16548
rect 23492 16492 23502 16548
rect 23986 16492 23996 16548
rect 24052 16492 24836 16548
rect 27794 16492 27804 16548
rect 27860 16492 29260 16548
rect 29316 16492 30828 16548
rect 30884 16492 32284 16548
rect 32340 16492 32350 16548
rect 41122 16492 41132 16548
rect 41188 16492 44604 16548
rect 44660 16492 46956 16548
rect 47012 16492 47022 16548
rect 47282 16492 47292 16548
rect 47348 16492 48524 16548
rect 48580 16492 48590 16548
rect 54114 16492 54124 16548
rect 54180 16492 54460 16548
rect 54516 16492 55356 16548
rect 55412 16492 56588 16548
rect 56644 16492 56654 16548
rect 23436 16436 23492 16492
rect 27804 16436 27860 16492
rect 23436 16380 27860 16436
rect 38546 16380 38556 16436
rect 38612 16380 40684 16436
rect 40740 16380 40750 16436
rect 47618 16380 47628 16436
rect 47684 16380 48412 16436
rect 48468 16380 48860 16436
rect 48916 16380 48926 16436
rect 49186 16380 49196 16436
rect 49252 16380 50092 16436
rect 50148 16380 51212 16436
rect 51268 16380 51278 16436
rect 52098 16380 52108 16436
rect 52164 16380 53228 16436
rect 53284 16380 53900 16436
rect 53956 16380 54908 16436
rect 54964 16380 54974 16436
rect 48860 16324 48916 16380
rect 28914 16268 28924 16324
rect 28980 16268 30380 16324
rect 30436 16268 30446 16324
rect 48860 16268 49420 16324
rect 49476 16268 49644 16324
rect 49700 16268 50540 16324
rect 50596 16268 52332 16324
rect 52388 16268 53676 16324
rect 53732 16268 55132 16324
rect 55188 16268 57484 16324
rect 57540 16268 57550 16324
rect 19826 16100 19836 16156
rect 19892 16100 19940 16156
rect 19996 16100 20044 16156
rect 20100 16100 20110 16156
rect 50546 16100 50556 16156
rect 50612 16100 50660 16156
rect 50716 16100 50764 16156
rect 50820 16100 50830 16156
rect 20178 16044 20188 16100
rect 20244 16044 20254 16100
rect 20188 15876 20244 16044
rect 27010 15932 27020 15988
rect 27076 15932 31276 15988
rect 31332 15932 31342 15988
rect 49074 15932 49084 15988
rect 49140 15932 51100 15988
rect 51156 15932 51166 15988
rect 20188 15820 23660 15876
rect 23716 15820 29148 15876
rect 29204 15820 29708 15876
rect 29764 15820 29774 15876
rect 35970 15820 35980 15876
rect 36036 15820 37100 15876
rect 37156 15820 37166 15876
rect 40226 15820 40236 15876
rect 40292 15820 41244 15876
rect 41300 15820 41310 15876
rect 48290 15820 48300 15876
rect 48356 15820 49196 15876
rect 49252 15820 49262 15876
rect 50082 15820 50092 15876
rect 50148 15820 50988 15876
rect 51044 15820 52108 15876
rect 52164 15820 52174 15876
rect 20188 15764 20244 15820
rect 19730 15708 19740 15764
rect 19796 15708 20244 15764
rect 28242 15708 28252 15764
rect 28308 15708 37548 15764
rect 37604 15708 37614 15764
rect 47506 15708 47516 15764
rect 47572 15708 48636 15764
rect 48692 15708 53004 15764
rect 53060 15708 53070 15764
rect 17714 15596 17724 15652
rect 17780 15596 19852 15652
rect 19908 15596 22092 15652
rect 22148 15596 22158 15652
rect 32050 15596 32060 15652
rect 32116 15596 32956 15652
rect 33012 15596 34412 15652
rect 34468 15596 34478 15652
rect 36306 15596 36316 15652
rect 36372 15596 37996 15652
rect 38052 15596 38062 15652
rect 48402 15596 48412 15652
rect 48468 15596 49868 15652
rect 49924 15596 54236 15652
rect 54292 15596 54302 15652
rect 24098 15484 24108 15540
rect 24164 15484 25228 15540
rect 25284 15484 25294 15540
rect 30930 15484 30940 15540
rect 30996 15484 33180 15540
rect 33236 15484 33246 15540
rect 47730 15484 47740 15540
rect 47796 15484 48972 15540
rect 49028 15484 49038 15540
rect 51202 15484 51212 15540
rect 51268 15484 51884 15540
rect 51940 15484 54460 15540
rect 54516 15484 54526 15540
rect 30594 15372 30604 15428
rect 30660 15372 31276 15428
rect 31332 15372 33628 15428
rect 33684 15372 34188 15428
rect 34244 15372 34254 15428
rect 31938 15260 31948 15316
rect 32004 15260 32396 15316
rect 32452 15260 32462 15316
rect 47068 15148 47628 15204
rect 47684 15148 47694 15204
rect 4466 15092 4476 15148
rect 4532 15092 4580 15148
rect 4636 15092 4684 15148
rect 4740 15092 4750 15148
rect 35186 15092 35196 15148
rect 35252 15092 35300 15148
rect 35356 15092 35404 15148
rect 35460 15092 35470 15148
rect 47068 15092 47124 15148
rect 19180 15036 20748 15092
rect 20804 15036 21420 15092
rect 21476 15036 21486 15092
rect 28354 15036 28364 15092
rect 28420 15036 31500 15092
rect 31556 15036 32508 15092
rect 32564 15036 33740 15092
rect 33796 15036 33806 15092
rect 45154 15036 45164 15092
rect 45220 15036 47124 15092
rect 19180 14756 19236 15036
rect 33170 14924 33180 14980
rect 33236 14924 36428 14980
rect 36484 14924 37884 14980
rect 37940 14924 37950 14980
rect 20178 14812 20188 14868
rect 20244 14812 25004 14868
rect 25060 14812 25070 14868
rect 17826 14700 17836 14756
rect 17892 14700 19180 14756
rect 19236 14700 19246 14756
rect 25330 14700 25340 14756
rect 25396 14700 26684 14756
rect 26740 14700 27132 14756
rect 27188 14700 27580 14756
rect 27636 14700 27646 14756
rect 32386 14700 32396 14756
rect 32452 14700 33292 14756
rect 33348 14700 37324 14756
rect 37380 14700 38668 14756
rect 38724 14700 38734 14756
rect 52658 14700 52668 14756
rect 52724 14700 56252 14756
rect 56308 14700 56318 14756
rect 17490 14588 17500 14644
rect 17556 14588 19628 14644
rect 19684 14588 20188 14644
rect 33730 14588 33740 14644
rect 33796 14588 35084 14644
rect 35140 14588 38220 14644
rect 38276 14588 38286 14644
rect 43474 14588 43484 14644
rect 43540 14588 43820 14644
rect 43876 14588 44940 14644
rect 44996 14588 45006 14644
rect 50530 14588 50540 14644
rect 50596 14588 52892 14644
rect 52948 14588 52958 14644
rect 20132 14420 20188 14588
rect 21410 14476 21420 14532
rect 21476 14476 23324 14532
rect 23380 14476 23390 14532
rect 25890 14476 25900 14532
rect 25956 14476 26684 14532
rect 26740 14476 28252 14532
rect 28308 14476 28318 14532
rect 41682 14476 41692 14532
rect 41748 14476 44268 14532
rect 44324 14476 45500 14532
rect 45556 14476 47068 14532
rect 47124 14476 47134 14532
rect 18386 14364 18396 14420
rect 18452 14364 19964 14420
rect 20020 14364 20030 14420
rect 20132 14364 21756 14420
rect 21812 14364 21822 14420
rect 22530 14364 22540 14420
rect 22596 14364 23548 14420
rect 23604 14364 23614 14420
rect 29698 14364 29708 14420
rect 29764 14364 30492 14420
rect 30548 14364 30940 14420
rect 30996 14364 31006 14420
rect 35522 14364 35532 14420
rect 35588 14364 36652 14420
rect 36708 14364 37772 14420
rect 37828 14364 37838 14420
rect 51538 14252 51548 14308
rect 51604 14252 51996 14308
rect 52052 14252 52668 14308
rect 52724 14252 52734 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 24434 13804 24444 13860
rect 24500 13804 25676 13860
rect 25732 13804 25742 13860
rect 52546 13804 52556 13860
rect 52612 13804 54572 13860
rect 54628 13804 56028 13860
rect 56084 13804 56094 13860
rect 16818 13692 16828 13748
rect 16884 13692 18284 13748
rect 18340 13692 18350 13748
rect 25330 13692 25340 13748
rect 25396 13692 28588 13748
rect 28644 13692 29708 13748
rect 29764 13692 29774 13748
rect 40002 13692 40012 13748
rect 40068 13692 45388 13748
rect 45444 13692 45454 13748
rect 20962 13580 20972 13636
rect 21028 13580 21756 13636
rect 21812 13580 21822 13636
rect 38994 13580 39004 13636
rect 39060 13580 39452 13636
rect 39508 13580 41132 13636
rect 41188 13580 43484 13636
rect 43540 13580 43550 13636
rect 24882 13468 24892 13524
rect 24948 13468 26236 13524
rect 26292 13468 27020 13524
rect 27076 13468 27086 13524
rect 23650 13356 23660 13412
rect 23716 13356 27244 13412
rect 27300 13356 30380 13412
rect 30436 13356 30446 13412
rect 4466 13076 4476 13132
rect 4532 13076 4580 13132
rect 4636 13076 4684 13132
rect 4740 13076 4750 13132
rect 35186 13076 35196 13132
rect 35252 13076 35300 13132
rect 35356 13076 35404 13132
rect 35460 13076 35470 13132
rect 27010 12684 27020 12740
rect 27076 12684 31612 12740
rect 31668 12684 33404 12740
rect 33460 12684 33740 12740
rect 33796 12684 33806 12740
rect 52770 12684 52780 12740
rect 52836 12684 55356 12740
rect 55412 12684 55422 12740
rect 35522 12348 35532 12404
rect 35588 12348 35980 12404
rect 36036 12348 37324 12404
rect 37380 12348 37660 12404
rect 37716 12348 38220 12404
rect 38276 12348 38892 12404
rect 38948 12348 38958 12404
rect 45378 12348 45388 12404
rect 45444 12348 46396 12404
rect 46452 12348 48860 12404
rect 48916 12348 48926 12404
rect 19826 12068 19836 12124
rect 19892 12068 19940 12124
rect 19996 12068 20044 12124
rect 20100 12068 20110 12124
rect 50546 12068 50556 12124
rect 50612 12068 50660 12124
rect 50716 12068 50764 12124
rect 50820 12068 50830 12124
rect 25218 11676 25228 11732
rect 25284 11676 25900 11732
rect 25956 11676 27132 11732
rect 27188 11676 30828 11732
rect 30884 11676 30894 11732
rect 37762 11676 37772 11732
rect 37828 11676 38556 11732
rect 38612 11676 38622 11732
rect 51874 11676 51884 11732
rect 51940 11676 53340 11732
rect 53396 11676 53406 11732
rect 18610 11564 18620 11620
rect 18676 11564 19740 11620
rect 19796 11564 21812 11620
rect 24434 11564 24444 11620
rect 24500 11564 25452 11620
rect 25508 11564 28812 11620
rect 28868 11564 29820 11620
rect 29876 11564 30380 11620
rect 30436 11564 30446 11620
rect 48850 11564 48860 11620
rect 48916 11564 52332 11620
rect 52388 11564 53116 11620
rect 53172 11564 53676 11620
rect 53732 11564 53742 11620
rect 21756 11508 21812 11564
rect 19394 11452 19404 11508
rect 19460 11452 20524 11508
rect 20580 11452 20590 11508
rect 21746 11452 21756 11508
rect 21812 11452 22988 11508
rect 23044 11452 23054 11508
rect 31154 11452 31164 11508
rect 31220 11452 33068 11508
rect 33124 11452 33134 11508
rect 29474 11340 29484 11396
rect 29540 11340 31948 11396
rect 32004 11340 35868 11396
rect 35924 11340 35934 11396
rect 4466 11060 4476 11116
rect 4532 11060 4580 11116
rect 4636 11060 4684 11116
rect 4740 11060 4750 11116
rect 35186 11060 35196 11116
rect 35252 11060 35300 11116
rect 35356 11060 35404 11116
rect 35460 11060 35470 11116
rect 22866 10892 22876 10948
rect 22932 10892 23996 10948
rect 24052 10892 24062 10948
rect 37314 10780 37324 10836
rect 37380 10780 38668 10836
rect 38724 10780 39228 10836
rect 39284 10780 41020 10836
rect 41076 10780 41580 10836
rect 41636 10780 42364 10836
rect 42420 10780 43596 10836
rect 43652 10780 45388 10836
rect 45444 10780 45454 10836
rect 18946 10668 18956 10724
rect 19012 10668 21420 10724
rect 21476 10668 21486 10724
rect 30370 10668 30380 10724
rect 30436 10668 31724 10724
rect 31780 10668 31948 10724
rect 35970 10668 35980 10724
rect 36036 10668 37772 10724
rect 37828 10668 37838 10724
rect 42018 10668 42028 10724
rect 42084 10668 43484 10724
rect 43540 10668 44492 10724
rect 44548 10668 44558 10724
rect 31892 10612 31948 10668
rect 31892 10556 32508 10612
rect 32564 10556 34188 10612
rect 34244 10556 34254 10612
rect 36530 10556 36540 10612
rect 36596 10556 38444 10612
rect 38500 10556 39116 10612
rect 39172 10556 41132 10612
rect 41188 10556 44044 10612
rect 44100 10556 44380 10612
rect 44436 10556 45164 10612
rect 45220 10556 45230 10612
rect 20738 10444 20748 10500
rect 20804 10444 22316 10500
rect 22372 10444 22382 10500
rect 32386 10444 32396 10500
rect 32452 10444 33628 10500
rect 33684 10444 33694 10500
rect 30156 10108 31164 10164
rect 31220 10108 31230 10164
rect 36428 10108 37324 10164
rect 37380 10108 37390 10164
rect 19826 10052 19836 10108
rect 19892 10052 19940 10108
rect 19996 10052 20044 10108
rect 20100 10052 20110 10108
rect 30156 10052 30212 10108
rect 36428 10052 36484 10108
rect 50546 10052 50556 10108
rect 50612 10052 50660 10108
rect 50716 10052 50764 10108
rect 50820 10052 50830 10108
rect 20290 9996 20300 10052
rect 20356 9996 21644 10052
rect 21700 9996 21710 10052
rect 26002 9996 26012 10052
rect 26068 9996 26796 10052
rect 26852 9996 29708 10052
rect 29764 9996 30212 10052
rect 33954 9996 33964 10052
rect 34020 9996 35196 10052
rect 35252 9996 36428 10052
rect 36484 9996 36494 10052
rect 18162 9772 18172 9828
rect 18228 9772 19068 9828
rect 19124 9772 19134 9828
rect 23426 9772 23436 9828
rect 23492 9772 23772 9828
rect 23828 9772 25676 9828
rect 25732 9772 25742 9828
rect 23986 9660 23996 9716
rect 24052 9660 24668 9716
rect 24724 9660 25228 9716
rect 25284 9660 26572 9716
rect 26628 9660 28140 9716
rect 28196 9660 28206 9716
rect 4466 9044 4476 9100
rect 4532 9044 4580 9100
rect 4636 9044 4684 9100
rect 4740 9044 4750 9100
rect 35186 9044 35196 9100
rect 35252 9044 35300 9100
rect 35356 9044 35404 9100
rect 35460 9044 35470 9100
rect 22082 8652 22092 8708
rect 22148 8652 22540 8708
rect 22596 8652 23772 8708
rect 23828 8652 23838 8708
rect 28130 8652 28140 8708
rect 28196 8652 29148 8708
rect 29204 8652 29596 8708
rect 29652 8652 29662 8708
rect 22978 8540 22988 8596
rect 23044 8540 23660 8596
rect 23716 8540 23726 8596
rect 28578 8540 28588 8596
rect 28644 8540 29260 8596
rect 29316 8540 29326 8596
rect 22866 8428 22876 8484
rect 22932 8428 23996 8484
rect 24052 8428 24062 8484
rect 27682 8428 27692 8484
rect 27748 8428 28700 8484
rect 28756 8428 28766 8484
rect 19826 8036 19836 8092
rect 19892 8036 19940 8092
rect 19996 8036 20044 8092
rect 20100 8036 20110 8092
rect 50546 8036 50556 8092
rect 50612 8036 50660 8092
rect 50716 8036 50764 8092
rect 50820 8036 50830 8092
rect 28252 7868 31612 7924
rect 31668 7868 31836 7924
rect 31892 7868 31902 7924
rect 28252 7812 28308 7868
rect 21298 7756 21308 7812
rect 21364 7756 22316 7812
rect 22372 7756 24892 7812
rect 24948 7756 28252 7812
rect 28308 7756 28318 7812
rect 29586 7756 29596 7812
rect 29652 7756 30380 7812
rect 30436 7756 30446 7812
rect 29138 7644 29148 7700
rect 29204 7644 30604 7700
rect 30660 7644 30670 7700
rect 30258 7532 30268 7588
rect 30324 7532 31724 7588
rect 31780 7532 31790 7588
rect 0 7476 800 7504
rect 0 7420 4284 7476
rect 4340 7420 4350 7476
rect 0 7392 800 7420
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 0 6804 800 6832
rect 0 6748 3836 6804
rect 3892 6748 3902 6804
rect 0 6720 800 6748
rect 19826 6020 19836 6076
rect 19892 6020 19940 6076
rect 19996 6020 20044 6076
rect 20100 6020 20110 6076
rect 50546 6020 50556 6076
rect 50612 6020 50660 6076
rect 50716 6020 50764 6076
rect 50820 6020 50830 6076
rect 4466 5012 4476 5068
rect 4532 5012 4580 5068
rect 4636 5012 4684 5068
rect 4740 5012 4750 5068
rect 35186 5012 35196 5068
rect 35252 5012 35300 5068
rect 35356 5012 35404 5068
rect 35460 5012 35470 5068
rect 19826 4004 19836 4060
rect 19892 4004 19940 4060
rect 19996 4004 20044 4060
rect 20100 4004 20110 4060
rect 50546 4004 50556 4060
rect 50612 4004 50660 4060
rect 50716 4004 50764 4060
rect 50820 4004 50830 4060
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55412 4532 55468
rect 4580 55412 4636 55468
rect 4684 55412 4740 55468
rect 35196 55412 35252 55468
rect 35300 55412 35356 55468
rect 35404 55412 35460 55468
rect 19836 54404 19892 54460
rect 19940 54404 19996 54460
rect 20044 54404 20100 54460
rect 50556 54404 50612 54460
rect 50660 54404 50716 54460
rect 50764 54404 50820 54460
rect 4476 53396 4532 53452
rect 4580 53396 4636 53452
rect 4684 53396 4740 53452
rect 35196 53396 35252 53452
rect 35300 53396 35356 53452
rect 35404 53396 35460 53452
rect 19836 52388 19892 52444
rect 19940 52388 19996 52444
rect 20044 52388 20100 52444
rect 50556 52388 50612 52444
rect 50660 52388 50716 52444
rect 50764 52388 50820 52444
rect 4476 51380 4532 51436
rect 4580 51380 4636 51436
rect 4684 51380 4740 51436
rect 35196 51380 35252 51436
rect 35300 51380 35356 51436
rect 35404 51380 35460 51436
rect 19836 50372 19892 50428
rect 19940 50372 19996 50428
rect 20044 50372 20100 50428
rect 50556 50372 50612 50428
rect 50660 50372 50716 50428
rect 50764 50372 50820 50428
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48356 19892 48412
rect 19940 48356 19996 48412
rect 20044 48356 20100 48412
rect 50556 48356 50612 48412
rect 50660 48356 50716 48412
rect 50764 48356 50820 48412
rect 4476 47348 4532 47404
rect 4580 47348 4636 47404
rect 4684 47348 4740 47404
rect 35196 47348 35252 47404
rect 35300 47348 35356 47404
rect 35404 47348 35460 47404
rect 19836 46340 19892 46396
rect 19940 46340 19996 46396
rect 20044 46340 20100 46396
rect 50556 46340 50612 46396
rect 50660 46340 50716 46396
rect 50764 46340 50820 46396
rect 4476 45332 4532 45388
rect 4580 45332 4636 45388
rect 4684 45332 4740 45388
rect 35196 45332 35252 45388
rect 35300 45332 35356 45388
rect 35404 45332 35460 45388
rect 19836 44324 19892 44380
rect 19940 44324 19996 44380
rect 20044 44324 20100 44380
rect 50556 44324 50612 44380
rect 50660 44324 50716 44380
rect 50764 44324 50820 44380
rect 4476 43316 4532 43372
rect 4580 43316 4636 43372
rect 4684 43316 4740 43372
rect 35196 43316 35252 43372
rect 35300 43316 35356 43372
rect 35404 43316 35460 43372
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41300 4532 41356
rect 4580 41300 4636 41356
rect 4684 41300 4740 41356
rect 35196 41300 35252 41356
rect 35300 41300 35356 41356
rect 35404 41300 35460 41356
rect 19836 40292 19892 40348
rect 19940 40292 19996 40348
rect 20044 40292 20100 40348
rect 50556 40292 50612 40348
rect 50660 40292 50716 40348
rect 50764 40292 50820 40348
rect 4476 39284 4532 39340
rect 4580 39284 4636 39340
rect 4684 39284 4740 39340
rect 35196 39284 35252 39340
rect 35300 39284 35356 39340
rect 35404 39284 35460 39340
rect 50204 38780 50260 38836
rect 19836 38276 19892 38332
rect 19940 38276 19996 38332
rect 20044 38276 20100 38332
rect 50556 38276 50612 38332
rect 50660 38276 50716 38332
rect 50764 38276 50820 38332
rect 4476 37268 4532 37324
rect 4580 37268 4636 37324
rect 4684 37268 4740 37324
rect 35196 37268 35252 37324
rect 35300 37268 35356 37324
rect 35404 37268 35460 37324
rect 50316 36540 50372 36596
rect 19836 36260 19892 36316
rect 19940 36260 19996 36316
rect 20044 36260 20100 36316
rect 50556 36260 50612 36316
rect 50660 36260 50716 36316
rect 50764 36260 50820 36316
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34244 19892 34300
rect 19940 34244 19996 34300
rect 20044 34244 20100 34300
rect 50556 34244 50612 34300
rect 50660 34244 50716 34300
rect 50764 34244 50820 34300
rect 4476 33236 4532 33292
rect 4580 33236 4636 33292
rect 4684 33236 4740 33292
rect 35196 33236 35252 33292
rect 35300 33236 35356 33292
rect 35404 33236 35460 33292
rect 19836 32228 19892 32284
rect 19940 32228 19996 32284
rect 20044 32228 20100 32284
rect 50556 32228 50612 32284
rect 50660 32228 50716 32284
rect 50764 32228 50820 32284
rect 4476 31220 4532 31276
rect 4580 31220 4636 31276
rect 4684 31220 4740 31276
rect 35196 31220 35252 31276
rect 35300 31220 35356 31276
rect 35404 31220 35460 31276
rect 19836 30212 19892 30268
rect 19940 30212 19996 30268
rect 20044 30212 20100 30268
rect 50556 30212 50612 30268
rect 50660 30212 50716 30268
rect 50764 30212 50820 30268
rect 4476 29204 4532 29260
rect 4580 29204 4636 29260
rect 4684 29204 4740 29260
rect 35196 29204 35252 29260
rect 35300 29204 35356 29260
rect 35404 29204 35460 29260
rect 26796 29036 26852 29092
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 35644 27804 35700 27860
rect 26796 27356 26852 27412
rect 4476 27188 4532 27244
rect 4580 27188 4636 27244
rect 4684 27188 4740 27244
rect 35196 27188 35252 27244
rect 35300 27188 35356 27244
rect 35404 27188 35460 27244
rect 19836 26180 19892 26236
rect 19940 26180 19996 26236
rect 20044 26180 20100 26236
rect 50556 26180 50612 26236
rect 50660 26180 50716 26236
rect 50764 26180 50820 26236
rect 35644 25788 35700 25844
rect 4476 25172 4532 25228
rect 4580 25172 4636 25228
rect 4684 25172 4740 25228
rect 35196 25172 35252 25228
rect 35300 25172 35356 25228
rect 35404 25172 35460 25228
rect 35644 24668 35700 24724
rect 19836 24164 19892 24220
rect 19940 24164 19996 24220
rect 20044 24164 20100 24220
rect 50556 24164 50612 24220
rect 50660 24164 50716 24220
rect 50764 24164 50820 24220
rect 4476 23156 4532 23212
rect 4580 23156 4636 23212
rect 4684 23156 4740 23212
rect 35196 23156 35252 23212
rect 35300 23156 35356 23212
rect 35404 23156 35460 23212
rect 19836 22148 19892 22204
rect 19940 22148 19996 22204
rect 20044 22148 20100 22204
rect 50556 22148 50612 22204
rect 50660 22148 50716 22204
rect 50764 22148 50820 22204
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20132 19892 20188
rect 19940 20132 19996 20188
rect 20044 20132 20100 20188
rect 50556 20132 50612 20188
rect 50660 20132 50716 20188
rect 50764 20132 50820 20188
rect 20188 19628 20244 19684
rect 4476 19124 4532 19180
rect 4580 19124 4636 19180
rect 4684 19124 4740 19180
rect 35196 19124 35252 19180
rect 35300 19124 35356 19180
rect 35404 19124 35460 19180
rect 19836 18116 19892 18172
rect 19940 18116 19996 18172
rect 20044 18116 20100 18172
rect 50556 18116 50612 18172
rect 50660 18116 50716 18172
rect 50764 18116 50820 18172
rect 4476 17108 4532 17164
rect 4580 17108 4636 17164
rect 4684 17108 4740 17164
rect 35196 17108 35252 17164
rect 35300 17108 35356 17164
rect 35404 17108 35460 17164
rect 19836 16100 19892 16156
rect 19940 16100 19996 16156
rect 20044 16100 20100 16156
rect 50556 16100 50612 16156
rect 50660 16100 50716 16156
rect 50764 16100 50820 16156
rect 20188 16044 20244 16100
rect 4476 15092 4532 15148
rect 4580 15092 4636 15148
rect 4684 15092 4740 15148
rect 35196 15092 35252 15148
rect 35300 15092 35356 15148
rect 35404 15092 35460 15148
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13076 4532 13132
rect 4580 13076 4636 13132
rect 4684 13076 4740 13132
rect 35196 13076 35252 13132
rect 35300 13076 35356 13132
rect 35404 13076 35460 13132
rect 19836 12068 19892 12124
rect 19940 12068 19996 12124
rect 20044 12068 20100 12124
rect 50556 12068 50612 12124
rect 50660 12068 50716 12124
rect 50764 12068 50820 12124
rect 4476 11060 4532 11116
rect 4580 11060 4636 11116
rect 4684 11060 4740 11116
rect 35196 11060 35252 11116
rect 35300 11060 35356 11116
rect 35404 11060 35460 11116
rect 19836 10052 19892 10108
rect 19940 10052 19996 10108
rect 20044 10052 20100 10108
rect 50556 10052 50612 10108
rect 50660 10052 50716 10108
rect 50764 10052 50820 10108
rect 4476 9044 4532 9100
rect 4580 9044 4636 9100
rect 4684 9044 4740 9100
rect 35196 9044 35252 9100
rect 35300 9044 35356 9100
rect 35404 9044 35460 9100
rect 19836 8036 19892 8092
rect 19940 8036 19996 8092
rect 20044 8036 20100 8092
rect 50556 8036 50612 8092
rect 50660 8036 50716 8092
rect 50764 8036 50820 8092
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6020 19892 6076
rect 19940 6020 19996 6076
rect 20044 6020 20100 6076
rect 50556 6020 50612 6076
rect 50660 6020 50716 6076
rect 50764 6020 50820 6076
rect 4476 5012 4532 5068
rect 4580 5012 4636 5068
rect 4684 5012 4740 5068
rect 35196 5012 35252 5068
rect 35300 5012 35356 5068
rect 35404 5012 35460 5068
rect 19836 4004 19892 4060
rect 19940 4004 19996 4060
rect 20044 4004 20100 4060
rect 50556 4004 50612 4060
rect 50660 4004 50716 4060
rect 50764 4004 50820 4060
<< metal4 >>
rect 4448 55468 4768 56508
rect 4448 55412 4476 55468
rect 4532 55412 4580 55468
rect 4636 55412 4684 55468
rect 4740 55412 4768 55468
rect 4448 53452 4768 55412
rect 4448 53396 4476 53452
rect 4532 53396 4580 53452
rect 4636 53396 4684 53452
rect 4740 53396 4768 53452
rect 4448 51436 4768 53396
rect 4448 51380 4476 51436
rect 4532 51380 4580 51436
rect 4636 51380 4684 51436
rect 4740 51380 4768 51436
rect 4448 49420 4768 51380
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47404 4768 49364
rect 4448 47348 4476 47404
rect 4532 47348 4580 47404
rect 4636 47348 4684 47404
rect 4740 47348 4768 47404
rect 4448 45388 4768 47348
rect 4448 45332 4476 45388
rect 4532 45332 4580 45388
rect 4636 45332 4684 45388
rect 4740 45332 4768 45388
rect 4448 43372 4768 45332
rect 4448 43316 4476 43372
rect 4532 43316 4580 43372
rect 4636 43316 4684 43372
rect 4740 43316 4768 43372
rect 4448 41356 4768 43316
rect 4448 41300 4476 41356
rect 4532 41300 4580 41356
rect 4636 41300 4684 41356
rect 4740 41300 4768 41356
rect 4448 39340 4768 41300
rect 4448 39284 4476 39340
rect 4532 39284 4580 39340
rect 4636 39284 4684 39340
rect 4740 39284 4768 39340
rect 4448 37324 4768 39284
rect 4448 37268 4476 37324
rect 4532 37268 4580 37324
rect 4636 37268 4684 37324
rect 4740 37268 4768 37324
rect 4448 35308 4768 37268
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33292 4768 35252
rect 4448 33236 4476 33292
rect 4532 33236 4580 33292
rect 4636 33236 4684 33292
rect 4740 33236 4768 33292
rect 4448 31276 4768 33236
rect 4448 31220 4476 31276
rect 4532 31220 4580 31276
rect 4636 31220 4684 31276
rect 4740 31220 4768 31276
rect 4448 29260 4768 31220
rect 4448 29204 4476 29260
rect 4532 29204 4580 29260
rect 4636 29204 4684 29260
rect 4740 29204 4768 29260
rect 4448 27244 4768 29204
rect 4448 27188 4476 27244
rect 4532 27188 4580 27244
rect 4636 27188 4684 27244
rect 4740 27188 4768 27244
rect 4448 25228 4768 27188
rect 4448 25172 4476 25228
rect 4532 25172 4580 25228
rect 4636 25172 4684 25228
rect 4740 25172 4768 25228
rect 4448 23212 4768 25172
rect 4448 23156 4476 23212
rect 4532 23156 4580 23212
rect 4636 23156 4684 23212
rect 4740 23156 4768 23212
rect 4448 21196 4768 23156
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19180 4768 21140
rect 4448 19124 4476 19180
rect 4532 19124 4580 19180
rect 4636 19124 4684 19180
rect 4740 19124 4768 19180
rect 4448 17164 4768 19124
rect 4448 17108 4476 17164
rect 4532 17108 4580 17164
rect 4636 17108 4684 17164
rect 4740 17108 4768 17164
rect 4448 15148 4768 17108
rect 4448 15092 4476 15148
rect 4532 15092 4580 15148
rect 4636 15092 4684 15148
rect 4740 15092 4768 15148
rect 4448 13132 4768 15092
rect 4448 13076 4476 13132
rect 4532 13076 4580 13132
rect 4636 13076 4684 13132
rect 4740 13076 4768 13132
rect 4448 11116 4768 13076
rect 4448 11060 4476 11116
rect 4532 11060 4580 11116
rect 4636 11060 4684 11116
rect 4740 11060 4768 11116
rect 4448 9100 4768 11060
rect 4448 9044 4476 9100
rect 4532 9044 4580 9100
rect 4636 9044 4684 9100
rect 4740 9044 4768 9100
rect 4448 7084 4768 9044
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5068 4768 7028
rect 4448 5012 4476 5068
rect 4532 5012 4580 5068
rect 4636 5012 4684 5068
rect 4740 5012 4768 5068
rect 4448 3972 4768 5012
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54460 20128 56420
rect 19808 54404 19836 54460
rect 19892 54404 19940 54460
rect 19996 54404 20044 54460
rect 20100 54404 20128 54460
rect 19808 52444 20128 54404
rect 19808 52388 19836 52444
rect 19892 52388 19940 52444
rect 19996 52388 20044 52444
rect 20100 52388 20128 52444
rect 19808 50428 20128 52388
rect 19808 50372 19836 50428
rect 19892 50372 19940 50428
rect 19996 50372 20044 50428
rect 20100 50372 20128 50428
rect 19808 48412 20128 50372
rect 19808 48356 19836 48412
rect 19892 48356 19940 48412
rect 19996 48356 20044 48412
rect 20100 48356 20128 48412
rect 19808 46396 20128 48356
rect 19808 46340 19836 46396
rect 19892 46340 19940 46396
rect 19996 46340 20044 46396
rect 20100 46340 20128 46396
rect 19808 44380 20128 46340
rect 19808 44324 19836 44380
rect 19892 44324 19940 44380
rect 19996 44324 20044 44380
rect 20100 44324 20128 44380
rect 19808 42364 20128 44324
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40348 20128 42308
rect 19808 40292 19836 40348
rect 19892 40292 19940 40348
rect 19996 40292 20044 40348
rect 20100 40292 20128 40348
rect 19808 38332 20128 40292
rect 19808 38276 19836 38332
rect 19892 38276 19940 38332
rect 19996 38276 20044 38332
rect 20100 38276 20128 38332
rect 19808 36316 20128 38276
rect 19808 36260 19836 36316
rect 19892 36260 19940 36316
rect 19996 36260 20044 36316
rect 20100 36260 20128 36316
rect 19808 34300 20128 36260
rect 19808 34244 19836 34300
rect 19892 34244 19940 34300
rect 19996 34244 20044 34300
rect 20100 34244 20128 34300
rect 19808 32284 20128 34244
rect 19808 32228 19836 32284
rect 19892 32228 19940 32284
rect 19996 32228 20044 32284
rect 20100 32228 20128 32284
rect 19808 30268 20128 32228
rect 19808 30212 19836 30268
rect 19892 30212 19940 30268
rect 19996 30212 20044 30268
rect 20100 30212 20128 30268
rect 19808 28252 20128 30212
rect 35168 55468 35488 56508
rect 35168 55412 35196 55468
rect 35252 55412 35300 55468
rect 35356 55412 35404 55468
rect 35460 55412 35488 55468
rect 35168 53452 35488 55412
rect 35168 53396 35196 53452
rect 35252 53396 35300 53452
rect 35356 53396 35404 53452
rect 35460 53396 35488 53452
rect 35168 51436 35488 53396
rect 35168 51380 35196 51436
rect 35252 51380 35300 51436
rect 35356 51380 35404 51436
rect 35460 51380 35488 51436
rect 35168 49420 35488 51380
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47404 35488 49364
rect 35168 47348 35196 47404
rect 35252 47348 35300 47404
rect 35356 47348 35404 47404
rect 35460 47348 35488 47404
rect 35168 45388 35488 47348
rect 35168 45332 35196 45388
rect 35252 45332 35300 45388
rect 35356 45332 35404 45388
rect 35460 45332 35488 45388
rect 35168 43372 35488 45332
rect 35168 43316 35196 43372
rect 35252 43316 35300 43372
rect 35356 43316 35404 43372
rect 35460 43316 35488 43372
rect 35168 41356 35488 43316
rect 35168 41300 35196 41356
rect 35252 41300 35300 41356
rect 35356 41300 35404 41356
rect 35460 41300 35488 41356
rect 35168 39340 35488 41300
rect 35168 39284 35196 39340
rect 35252 39284 35300 39340
rect 35356 39284 35404 39340
rect 35460 39284 35488 39340
rect 35168 37324 35488 39284
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54460 50848 56420
rect 50528 54404 50556 54460
rect 50612 54404 50660 54460
rect 50716 54404 50764 54460
rect 50820 54404 50848 54460
rect 50528 52444 50848 54404
rect 50528 52388 50556 52444
rect 50612 52388 50660 52444
rect 50716 52388 50764 52444
rect 50820 52388 50848 52444
rect 50528 50428 50848 52388
rect 50528 50372 50556 50428
rect 50612 50372 50660 50428
rect 50716 50372 50764 50428
rect 50820 50372 50848 50428
rect 50528 48412 50848 50372
rect 50528 48356 50556 48412
rect 50612 48356 50660 48412
rect 50716 48356 50764 48412
rect 50820 48356 50848 48412
rect 50528 46396 50848 48356
rect 50528 46340 50556 46396
rect 50612 46340 50660 46396
rect 50716 46340 50764 46396
rect 50820 46340 50848 46396
rect 50528 44380 50848 46340
rect 50528 44324 50556 44380
rect 50612 44324 50660 44380
rect 50716 44324 50764 44380
rect 50820 44324 50848 44380
rect 50528 42364 50848 44324
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40348 50848 42308
rect 50528 40292 50556 40348
rect 50612 40292 50660 40348
rect 50716 40292 50764 40348
rect 50820 40292 50848 40348
rect 50204 38836 50260 38846
rect 50204 38668 50260 38780
rect 50204 38612 50372 38668
rect 35168 37268 35196 37324
rect 35252 37268 35300 37324
rect 35356 37268 35404 37324
rect 35460 37268 35488 37324
rect 35168 35308 35488 37268
rect 50316 36596 50372 38612
rect 50316 36530 50372 36540
rect 50528 38332 50848 40292
rect 50528 38276 50556 38332
rect 50612 38276 50660 38332
rect 50716 38276 50764 38332
rect 50820 38276 50848 38332
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33292 35488 35252
rect 35168 33236 35196 33292
rect 35252 33236 35300 33292
rect 35356 33236 35404 33292
rect 35460 33236 35488 33292
rect 35168 31276 35488 33236
rect 35168 31220 35196 31276
rect 35252 31220 35300 31276
rect 35356 31220 35404 31276
rect 35460 31220 35488 31276
rect 35168 29260 35488 31220
rect 35168 29204 35196 29260
rect 35252 29204 35300 29260
rect 35356 29204 35404 29260
rect 35460 29204 35488 29260
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26236 20128 28196
rect 26796 29092 26852 29102
rect 26796 27412 26852 29036
rect 26796 27346 26852 27356
rect 19808 26180 19836 26236
rect 19892 26180 19940 26236
rect 19996 26180 20044 26236
rect 20100 26180 20128 26236
rect 19808 24220 20128 26180
rect 19808 24164 19836 24220
rect 19892 24164 19940 24220
rect 19996 24164 20044 24220
rect 20100 24164 20128 24220
rect 19808 22204 20128 24164
rect 19808 22148 19836 22204
rect 19892 22148 19940 22204
rect 19996 22148 20044 22204
rect 20100 22148 20128 22204
rect 19808 20188 20128 22148
rect 19808 20132 19836 20188
rect 19892 20132 19940 20188
rect 19996 20132 20044 20188
rect 20100 20132 20128 20188
rect 19808 18172 20128 20132
rect 35168 27244 35488 29204
rect 50528 36316 50848 38276
rect 50528 36260 50556 36316
rect 50612 36260 50660 36316
rect 50716 36260 50764 36316
rect 50820 36260 50848 36316
rect 50528 34300 50848 36260
rect 50528 34244 50556 34300
rect 50612 34244 50660 34300
rect 50716 34244 50764 34300
rect 50820 34244 50848 34300
rect 50528 32284 50848 34244
rect 50528 32228 50556 32284
rect 50612 32228 50660 32284
rect 50716 32228 50764 32284
rect 50820 32228 50848 32284
rect 50528 30268 50848 32228
rect 50528 30212 50556 30268
rect 50612 30212 50660 30268
rect 50716 30212 50764 30268
rect 50820 30212 50848 30268
rect 50528 28252 50848 30212
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 35168 27188 35196 27244
rect 35252 27188 35300 27244
rect 35356 27188 35404 27244
rect 35460 27188 35488 27244
rect 35168 25228 35488 27188
rect 35168 25172 35196 25228
rect 35252 25172 35300 25228
rect 35356 25172 35404 25228
rect 35460 25172 35488 25228
rect 35168 23212 35488 25172
rect 35644 27860 35700 27870
rect 35644 25844 35700 27804
rect 35644 24724 35700 25788
rect 35644 24658 35700 24668
rect 50528 26236 50848 28196
rect 50528 26180 50556 26236
rect 50612 26180 50660 26236
rect 50716 26180 50764 26236
rect 50820 26180 50848 26236
rect 35168 23156 35196 23212
rect 35252 23156 35300 23212
rect 35356 23156 35404 23212
rect 35460 23156 35488 23212
rect 35168 21196 35488 23156
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 18116 19836 18172
rect 19892 18116 19940 18172
rect 19996 18116 20044 18172
rect 20100 18116 20128 18172
rect 19808 16156 20128 18116
rect 19808 16100 19836 16156
rect 19892 16100 19940 16156
rect 19996 16100 20044 16156
rect 20100 16100 20128 16156
rect 19808 14140 20128 16100
rect 20188 19684 20244 19694
rect 20188 16100 20244 19628
rect 20188 16034 20244 16044
rect 35168 19180 35488 21140
rect 35168 19124 35196 19180
rect 35252 19124 35300 19180
rect 35356 19124 35404 19180
rect 35460 19124 35488 19180
rect 35168 17164 35488 19124
rect 35168 17108 35196 17164
rect 35252 17108 35300 17164
rect 35356 17108 35404 17164
rect 35460 17108 35488 17164
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12124 20128 14084
rect 19808 12068 19836 12124
rect 19892 12068 19940 12124
rect 19996 12068 20044 12124
rect 20100 12068 20128 12124
rect 19808 10108 20128 12068
rect 19808 10052 19836 10108
rect 19892 10052 19940 10108
rect 19996 10052 20044 10108
rect 20100 10052 20128 10108
rect 19808 8092 20128 10052
rect 19808 8036 19836 8092
rect 19892 8036 19940 8092
rect 19996 8036 20044 8092
rect 20100 8036 20128 8092
rect 19808 6076 20128 8036
rect 19808 6020 19836 6076
rect 19892 6020 19940 6076
rect 19996 6020 20044 6076
rect 20100 6020 20128 6076
rect 19808 4060 20128 6020
rect 19808 4004 19836 4060
rect 19892 4004 19940 4060
rect 19996 4004 20044 4060
rect 20100 4004 20128 4060
rect 19808 3972 20128 4004
rect 35168 15148 35488 17108
rect 35168 15092 35196 15148
rect 35252 15092 35300 15148
rect 35356 15092 35404 15148
rect 35460 15092 35488 15148
rect 35168 13132 35488 15092
rect 35168 13076 35196 13132
rect 35252 13076 35300 13132
rect 35356 13076 35404 13132
rect 35460 13076 35488 13132
rect 35168 11116 35488 13076
rect 35168 11060 35196 11116
rect 35252 11060 35300 11116
rect 35356 11060 35404 11116
rect 35460 11060 35488 11116
rect 35168 9100 35488 11060
rect 35168 9044 35196 9100
rect 35252 9044 35300 9100
rect 35356 9044 35404 9100
rect 35460 9044 35488 9100
rect 35168 7084 35488 9044
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5068 35488 7028
rect 35168 5012 35196 5068
rect 35252 5012 35300 5068
rect 35356 5012 35404 5068
rect 35460 5012 35488 5068
rect 35168 3972 35488 5012
rect 50528 24220 50848 26180
rect 50528 24164 50556 24220
rect 50612 24164 50660 24220
rect 50716 24164 50764 24220
rect 50820 24164 50848 24220
rect 50528 22204 50848 24164
rect 50528 22148 50556 22204
rect 50612 22148 50660 22204
rect 50716 22148 50764 22204
rect 50820 22148 50848 22204
rect 50528 20188 50848 22148
rect 50528 20132 50556 20188
rect 50612 20132 50660 20188
rect 50716 20132 50764 20188
rect 50820 20132 50848 20188
rect 50528 18172 50848 20132
rect 50528 18116 50556 18172
rect 50612 18116 50660 18172
rect 50716 18116 50764 18172
rect 50820 18116 50848 18172
rect 50528 16156 50848 18116
rect 50528 16100 50556 16156
rect 50612 16100 50660 16156
rect 50716 16100 50764 16156
rect 50820 16100 50848 16156
rect 50528 14140 50848 16100
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12124 50848 14084
rect 50528 12068 50556 12124
rect 50612 12068 50660 12124
rect 50716 12068 50764 12124
rect 50820 12068 50848 12124
rect 50528 10108 50848 12068
rect 50528 10052 50556 10108
rect 50612 10052 50660 10108
rect 50716 10052 50764 10108
rect 50820 10052 50848 10108
rect 50528 8092 50848 10052
rect 50528 8036 50556 8092
rect 50612 8036 50660 8092
rect 50716 8036 50764 8092
rect 50820 8036 50848 8092
rect 50528 6076 50848 8036
rect 50528 6020 50556 6076
rect 50612 6020 50660 6076
rect 50716 6020 50764 6076
rect 50820 6020 50848 6076
rect 50528 4060 50848 6020
rect 50528 4004 50556 4060
rect 50612 4004 50660 4060
rect 50716 4004 50764 4060
rect 50820 4004 50848 4060
rect 50528 3972 50848 4004
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _244_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _245_
timestamp 1698431365
transform 1 0 28000 0 -1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _246_
timestamp 1698431365
transform -1 0 28336 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _247_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 40544 0 -1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _248_
timestamp 1698431365
transform -1 0 40544 0 -1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _249_
timestamp 1698431365
transform 1 0 45248 0 1 16128
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _250_
timestamp 1698431365
transform -1 0 37520 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _251_
timestamp 1698431365
transform 1 0 39312 0 1 18144
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _252_
timestamp 1698431365
transform 1 0 46816 0 1 16128
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _253_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 -1 18144
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _254_
timestamp 1698431365
transform 1 0 52528 0 -1 16128
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _255_
timestamp 1698431365
transform 1 0 46816 0 1 18144
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _256_
timestamp 1698431365
transform 1 0 48160 0 1 14112
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _257_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 35056 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _258_
timestamp 1698431365
transform 1 0 45024 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _259_
timestamp 1698431365
transform -1 0 48384 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _260_
timestamp 1698431365
transform 1 0 38080 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _261_
timestamp 1698431365
transform 1 0 40656 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _262_
timestamp 1698431365
transform -1 0 48160 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _263_
timestamp 1698431365
transform 1 0 48608 0 -1 20160
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _264_
timestamp 1698431365
transform -1 0 35280 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _265_
timestamp 1698431365
transform -1 0 35056 0 1 24192
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _266_
timestamp 1698431365
transform -1 0 40432 0 1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _267_
timestamp 1698431365
transform -1 0 30240 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _268_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29344 0 -1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _269_
timestamp 1698431365
transform -1 0 31920 0 -1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _270_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 30128 0 -1 22176
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _271_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 30016 0 1 24192
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _272_
timestamp 1698431365
transform -1 0 34832 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _273_
timestamp 1698431365
transform -1 0 36624 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _274_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 26208
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _275_
timestamp 1698431365
transform -1 0 29008 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _276_
timestamp 1698431365
transform 1 0 40208 0 1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _277_
timestamp 1698431365
transform 1 0 42896 0 -1 22176
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _278_
timestamp 1698431365
transform 1 0 44912 0 -1 14112
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _279_
timestamp 1698431365
transform 1 0 33152 0 -1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _280_
timestamp 1698431365
transform 1 0 43008 0 1 20160
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _281_
timestamp 1698431365
transform -1 0 42000 0 -1 22176
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _282_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 -1 26208
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _283_
timestamp 1698431365
transform -1 0 24864 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _284_
timestamp 1698431365
transform -1 0 27328 0 1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _285_
timestamp 1698431365
transform 1 0 14560 0 1 30240
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _286_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 16576 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _287_
timestamp 1698431365
transform -1 0 28336 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _288_
timestamp 1698431365
transform 1 0 29008 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _289_
timestamp 1698431365
transform -1 0 41440 0 -1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _290_
timestamp 1698431365
transform 1 0 39312 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _291_
timestamp 1698431365
transform 1 0 39088 0 1 44352
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _292_
timestamp 1698431365
transform 1 0 48832 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _293_
timestamp 1698431365
transform -1 0 50848 0 1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _294_
timestamp 1698431365
transform 1 0 42896 0 -1 42336
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _295_
timestamp 1698431365
transform -1 0 44464 0 1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _296_
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _297_
timestamp 1698431365
transform 1 0 38976 0 1 46368
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _298_
timestamp 1698431365
transform 1 0 42672 0 1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _299_
timestamp 1698431365
transform -1 0 50064 0 1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _300_
timestamp 1698431365
transform 1 0 48608 0 -1 46368
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _301_
timestamp 1698431365
transform 1 0 41664 0 -1 44352
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _302_
timestamp 1698431365
transform 1 0 41440 0 -1 42336
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _303_
timestamp 1698431365
transform -1 0 31024 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _304_
timestamp 1698431365
transform 1 0 40768 0 -1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _305_
timestamp 1698431365
transform -1 0 26880 0 1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _306_
timestamp 1698431365
transform 1 0 39536 0 1 16128
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _307_
timestamp 1698431365
transform 1 0 34048 0 -1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _308_
timestamp 1698431365
transform 1 0 35168 0 -1 14112
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _309_
timestamp 1698431365
transform 1 0 37520 0 -1 16128
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _310_
timestamp 1698431365
transform -1 0 33600 0 1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _311_
timestamp 1698431365
transform -1 0 38976 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _312_
timestamp 1698431365
transform -1 0 39088 0 -1 24192
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__nand3_1  _313_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32256 0 1 24192
box -86 -90 870 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _314_
timestamp 1698431365
transform -1 0 40208 0 1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _315_
timestamp 1698431365
transform 1 0 32928 0 -1 40320
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _316_
timestamp 1698431365
transform -1 0 32256 0 -1 28224
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_1  _317_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 31808 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _318_
timestamp 1698431365
transform -1 0 28784 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _319_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 28000 0 1 26208
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__nor3_1  _320_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _321_
timestamp 1698431365
transform 1 0 15456 0 1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _322_
timestamp 1698431365
transform 1 0 33040 0 -1 18144
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _323_
timestamp 1698431365
transform -1 0 32032 0 -1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _324_
timestamp 1698431365
transform -1 0 30688 0 1 18144
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _325_
timestamp 1698431365
transform -1 0 34048 0 -1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _326_
timestamp 1698431365
transform 1 0 29904 0 1 12096
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _327_
timestamp 1698431365
transform 1 0 31248 0 -1 16128
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _328_
timestamp 1698431365
transform -1 0 30912 0 1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _329_
timestamp 1698431365
transform -1 0 27888 0 1 24192
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _330_
timestamp 1698431365
transform 1 0 15232 0 1 22176
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _331_
timestamp 1698431365
transform 1 0 26096 0 -1 24192
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _332_
timestamp 1698431365
transform -1 0 38640 0 1 24192
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _333_
timestamp 1698431365
transform 1 0 33152 0 1 22176
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _334_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 38416 0 -1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _335_
timestamp 1698431365
transform 1 0 37408 0 -1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _336_
timestamp 1698431365
transform 1 0 36848 0 1 24192
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _337_
timestamp 1698431365
transform 1 0 30240 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _338_
timestamp 1698431365
transform -1 0 41440 0 1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _339_
timestamp 1698431365
transform 1 0 39088 0 -1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _340_
timestamp 1698431365
transform 1 0 38976 0 1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _341_
timestamp 1698431365
transform 1 0 36064 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _342_
timestamp 1698431365
transform 1 0 36736 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _343_
timestamp 1698431365
transform -1 0 39312 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _344_
timestamp 1698431365
transform 1 0 36848 0 1 38304
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _345_
timestamp 1698431365
transform 1 0 36848 0 1 34272
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _346_
timestamp 1698431365
transform -1 0 38192 0 -1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _347_
timestamp 1698431365
transform -1 0 34272 0 1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _348_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _349_
timestamp 1698431365
transform 1 0 31920 0 -1 40320
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _350_
timestamp 1698431365
transform 1 0 33152 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _351_
timestamp 1698431365
transform 1 0 32256 0 1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _352_
timestamp 1698431365
transform -1 0 33264 0 1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _353_
timestamp 1698431365
transform -1 0 44464 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _354_
timestamp 1698431365
transform -1 0 51184 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _355_
timestamp 1698431365
transform 1 0 44576 0 -1 30240
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _356_
timestamp 1698431365
transform -1 0 38080 0 1 30240
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _357_
timestamp 1698431365
transform 1 0 34160 0 1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_1  _358_
timestamp 1698431365
transform 1 0 35280 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _359_
timestamp 1698431365
transform -1 0 29344 0 -1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _360_
timestamp 1698431365
transform 1 0 26544 0 -1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _361_
timestamp 1698431365
transform 1 0 16912 0 1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _362_
timestamp 1698431365
transform 1 0 26656 0 -1 18144
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _363_
timestamp 1698431365
transform 1 0 23184 0 1 12096
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _364_
timestamp 1698431365
transform -1 0 31696 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _365_
timestamp 1698431365
transform 1 0 25760 0 -1 20160
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _366_
timestamp 1698431365
transform -1 0 18704 0 -1 20160
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _367_
timestamp 1698431365
transform 1 0 24640 0 1 22176
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _368_
timestamp 1698431365
transform 1 0 48496 0 1 38304
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _369_
timestamp 1698431365
transform 1 0 52640 0 1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _370_
timestamp 1698431365
transform 1 0 52528 0 1 40320
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _371_
timestamp 1698431365
transform 1 0 48608 0 -1 40320
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _372_
timestamp 1698431365
transform 1 0 52528 0 1 44352
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _373_
timestamp 1698431365
transform 1 0 51408 0 1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _374_
timestamp 1698431365
transform 1 0 52752 0 -1 40320
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _375_
timestamp 1698431365
transform 1 0 49504 0 1 40320
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _376_
timestamp 1698431365
transform 1 0 47264 0 1 40320
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _377_
timestamp 1698431365
transform -1 0 30352 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _378_
timestamp 1698431365
transform 1 0 25088 0 1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _379_
timestamp 1698431365
transform 1 0 13888 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _380_
timestamp 1698431365
transform 1 0 15008 0 -1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _381_
timestamp 1698431365
transform 1 0 22736 0 1 14112
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _382_
timestamp 1698431365
transform -1 0 30912 0 -1 40320
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _383_
timestamp 1698431365
transform 1 0 31808 0 -1 46368
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _384_
timestamp 1698431365
transform 1 0 23520 0 1 48384
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _385_
timestamp 1698431365
transform -1 0 26096 0 1 24192
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _386_
timestamp 1698431365
transform 1 0 25088 0 -1 22176
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _387_
timestamp 1698431365
transform 1 0 26096 0 1 24192
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _388_
timestamp 1698431365
transform 1 0 25088 0 -1 24192
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _389_
timestamp 1698431365
transform -1 0 38640 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _390_
timestamp 1698431365
transform 1 0 36400 0 -1 24192
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _391_
timestamp 1698431365
transform 1 0 41216 0 1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _392_
timestamp 1698431365
transform -1 0 39088 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _393_
timestamp 1698431365
transform 1 0 40320 0 1 38304
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _394_
timestamp 1698431365
transform -1 0 39088 0 1 34272
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _395_
timestamp 1698431365
transform 1 0 36960 0 1 26208
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _396_
timestamp 1698431365
transform 1 0 34608 0 1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _397_
timestamp 1698431365
transform 1 0 35952 0 -1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _398_
timestamp 1698431365
transform 1 0 34608 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _399_
timestamp 1698431365
transform -1 0 34496 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _400_
timestamp 1698431365
transform 1 0 44912 0 -1 32256
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _401_
timestamp 1698431365
transform -1 0 38640 0 1 30240
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _402_
timestamp 1698431365
transform 1 0 35280 0 -1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_1  _403_
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _404_
timestamp 1698431365
transform 1 0 27328 0 1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _405_
timestamp 1698431365
transform 1 0 14000 0 1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _406_
timestamp 1698431365
transform -1 0 29680 0 1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _407_
timestamp 1698431365
transform 1 0 30352 0 1 44352
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _408_
timestamp 1698431365
transform 1 0 32928 0 -1 46368
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _409_
timestamp 1698431365
transform 1 0 29792 0 -1 42336
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _410_
timestamp 1698431365
transform 1 0 27328 0 1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _411_
timestamp 1698431365
transform 1 0 26656 0 -1 34272
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _412_
timestamp 1698431365
transform 1 0 52080 0 -1 38304
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _413_
timestamp 1698431365
transform -1 0 55216 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _414_
timestamp 1698431365
transform 1 0 52752 0 -1 32256
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _415_
timestamp 1698431365
transform 1 0 50848 0 1 32256
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _416_
timestamp 1698431365
transform 1 0 52752 0 -1 36288
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _417_
timestamp 1698431365
transform 1 0 52528 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _418_
timestamp 1698431365
transform 1 0 52752 0 -1 30240
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _419_
timestamp 1698431365
transform 1 0 52192 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _420_
timestamp 1698431365
transform 1 0 49392 0 -1 32256
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _421_
timestamp 1698431365
transform -1 0 31696 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _422_
timestamp 1698431365
transform -1 0 27664 0 1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _423_
timestamp 1698431365
transform 1 0 13888 0 -1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _424_
timestamp 1698431365
transform 1 0 23632 0 1 38304
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _425_
timestamp 1698431365
transform 1 0 22960 0 1 42336
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _426_
timestamp 1698431365
transform 1 0 26992 0 -1 42336
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _427_
timestamp 1698431365
transform 1 0 25424 0 -1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _428_
timestamp 1698431365
transform 1 0 24752 0 1 34272
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _429_
timestamp 1698431365
transform -1 0 37744 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _430_
timestamp 1698431365
transform -1 0 36400 0 -1 24192
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _431_
timestamp 1698431365
transform 1 0 39760 0 1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _432_
timestamp 1698431365
transform -1 0 39536 0 1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _433_
timestamp 1698431365
transform 1 0 38976 0 1 36288
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _434_
timestamp 1698431365
transform -1 0 38528 0 1 34272
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _435_
timestamp 1698431365
transform 1 0 36512 0 -1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _436_
timestamp 1698431365
transform 1 0 34384 0 -1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _437_
timestamp 1698431365
transform 1 0 35168 0 -1 26208
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _438_
timestamp 1698431365
transform -1 0 32704 0 -1 38304
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _439_
timestamp 1698431365
transform 1 0 33264 0 1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _440_
timestamp 1698431365
transform 1 0 39312 0 1 32256
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _441_
timestamp 1698431365
transform -1 0 37520 0 -1 32256
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _442_
timestamp 1698431365
transform 1 0 34832 0 1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_1  _443_
timestamp 1698431365
transform -1 0 34272 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _444_
timestamp 1698431365
transform 1 0 26544 0 -1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _445_
timestamp 1698431365
transform 1 0 14336 0 -1 32256
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _446_
timestamp 1698431365
transform 1 0 52528 0 1 22176
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _447_
timestamp 1698431365
transform 1 0 52528 0 1 26208
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _448_
timestamp 1698431365
transform 1 0 50848 0 1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _449_
timestamp 1698431365
transform 1 0 52752 0 -1 24192
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _450_
timestamp 1698431365
transform 1 0 44912 0 -1 26208
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _451_
timestamp 1698431365
transform -1 0 44912 0 -1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _452_
timestamp 1698431365
transform 1 0 44688 0 1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _453_
timestamp 1698431365
transform -1 0 28672 0 1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _454_
timestamp 1698431365
transform 1 0 21168 0 1 22176
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _455_
timestamp 1698431365
transform 1 0 21056 0 -1 26208
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _456_
timestamp 1698431365
transform -1 0 24640 0 1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _457_
timestamp 1698431365
transform -1 0 26656 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi221_1  _458_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 26544 0 -1 28224
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__nor3_1  _459_
timestamp 1698431365
transform -1 0 25088 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _460_
timestamp 1698431365
transform 1 0 12096 0 -1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _461_
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _462_
timestamp 1698431365
transform 1 0 22848 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__or4_1  _463_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 26544 0 -1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _464_
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _465_
timestamp 1698431365
transform 1 0 21392 0 -1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _466_
timestamp 1698431365
transform 1 0 18480 0 -1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _467_
timestamp 1698431365
transform 1 0 18704 0 1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _468_
timestamp 1698431365
transform 1 0 17472 0 1 30240
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _469_
timestamp 1698431365
transform -1 0 12656 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _470_
timestamp 1698431365
transform -1 0 22624 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _471_
timestamp 1698431365
transform -1 0 23072 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _472_
timestamp 1698431365
transform 1 0 20720 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__oai31_1  _473_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21840 0 -1 34272
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _474_
timestamp 1698431365
transform -1 0 26096 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _475_
timestamp 1698431365
transform -1 0 27216 0 1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _476_
timestamp 1698431365
transform -1 0 30576 0 1 32256
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _477_
timestamp 1698431365
transform -1 0 32368 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _478_
timestamp 1698431365
transform 1 0 20272 0 1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _479_
timestamp 1698431365
transform 1 0 21168 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _480_
timestamp 1698431365
transform -1 0 26096 0 -1 34272
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _481_
timestamp 1698431365
transform -1 0 25424 0 1 32256
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _482_
timestamp 1698431365
transform -1 0 24416 0 1 32256
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _483_
timestamp 1698431365
transform 1 0 23408 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _484_
timestamp 1698431365
transform -1 0 21280 0 -1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _485_
timestamp 1698431365
transform 1 0 21168 0 1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _486_
timestamp 1698431365
transform 1 0 17248 0 1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _487_
timestamp 1698431365
transform 1 0 18704 0 1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _488_
timestamp 1698431365
transform 1 0 17696 0 -1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _489_
timestamp 1698431365
transform 1 0 19152 0 -1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _490_
timestamp 1698431365
transform 1 0 20048 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  _491_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 13776 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__nand4_1  _492_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 22176 0 1 34272
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _493_
timestamp 1698431365
transform 1 0 20384 0 -1 32256
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _494_
timestamp 1698431365
transform 1 0 18592 0 1 32256
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _495_
timestamp 1698431365
transform 1 0 17808 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _496_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 26880 0 -1 36288
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _497_
timestamp 1698431365
transform 1 0 30576 0 1 32256
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _498_
timestamp 1698431365
transform 1 0 30800 0 1 34272
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _499_
timestamp 1698431365
transform 1 0 29568 0 -1 32256
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _500_
timestamp 1698431365
transform 1 0 25088 0 -1 32256
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _501_
timestamp 1698431365
transform 1 0 23072 0 1 30240
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _502_
timestamp 1698431365
transform -1 0 24864 0 -1 36288
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _503_
timestamp 1698431365
transform -1 0 19712 0 1 36288
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _504_
timestamp 1698431365
transform 1 0 16352 0 1 40320
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _505_
timestamp 1698431365
transform -1 0 20160 0 1 38304
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _506_
timestamp 1698431365
transform 1 0 17248 0 -1 40320
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _507_
timestamp 1698431365
transform 1 0 17472 0 -1 38304
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _508_
timestamp 1698431365
transform 1 0 9968 0 1 32256
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _509_
timestamp 1698431365
transform -1 0 21392 0 -1 30240
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _510_
timestamp 1698431365
transform 1 0 17248 0 -1 32256
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _511_
timestamp 1698431365
transform 1 0 15456 0 1 32256
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  _512_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 9632 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  _513_
timestamp 1698431365
transform -1 0 4144 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  _514_
timestamp 1698431365
transform 1 0 55776 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  _515_
timestamp 1698431365
transform -1 0 4144 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  _516_
timestamp 1698431365
transform -1 0 4592 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__249__I test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 45024 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__250__I
timestamp 1698431365
transform 1 0 36624 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__262__I
timestamp 1698431365
transform 1 0 48384 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__263__S0
timestamp 1698431365
transform 1 0 48832 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__263__S1
timestamp 1698431365
transform -1 0 48384 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__264__I
timestamp 1698431365
transform -1 0 34832 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__269__I
timestamp 1698431365
transform 1 0 32144 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__270__S
timestamp 1698431365
transform 1 0 30352 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__280__S
timestamp 1698431365
transform 1 0 42784 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__281__A1
timestamp 1698431365
transform 1 0 42672 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__284__A2
timestamp 1698431365
transform 1 0 29232 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__290__I
timestamp 1698431365
transform -1 0 39312 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__291__S0
timestamp 1698431365
transform 1 0 44016 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__291__S1
timestamp 1698431365
transform -1 0 43904 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__292__I
timestamp 1698431365
transform 1 0 49728 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__294__S0
timestamp 1698431365
transform 1 0 42672 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__294__S1
timestamp 1698431365
transform 1 0 46592 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__297__S0
timestamp 1698431365
transform -1 0 43232 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__297__S1
timestamp 1698431365
transform 1 0 44128 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__300__S1
timestamp 1698431365
transform 1 0 54096 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__302__S
timestamp 1698431365
transform -1 0 41440 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__303__A2
timestamp 1698431365
transform -1 0 32144 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__305__I
timestamp 1698431365
transform -1 0 26208 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__308__S0
timestamp 1698431365
transform 1 0 39200 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__309__S
timestamp 1698431365
transform 1 0 37296 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__319__A2
timestamp 1698431365
transform 1 0 28000 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__322__S0
timestamp 1698431365
transform 1 0 36736 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__324__I
timestamp 1698431365
transform 1 0 30912 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__326__S1
timestamp 1698431365
transform -1 0 33824 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__327__S
timestamp 1698431365
transform -1 0 33376 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__328__I
timestamp 1698431365
transform 1 0 31136 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__330__S
timestamp 1698431365
transform 1 0 16912 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__333__I
timestamp 1698431365
transform 1 0 32480 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__338__I
timestamp 1698431365
transform 1 0 43008 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__339__S
timestamp 1698431365
transform 1 0 41216 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__340__B
timestamp 1698431365
transform 1 0 40320 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__349__I
timestamp 1698431365
transform 1 0 31696 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__357__B
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__363__S1
timestamp 1698431365
transform -1 0 27104 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__365__S
timestamp 1698431365
transform -1 0 27440 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__366__S
timestamp 1698431365
transform 1 0 18256 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__368__S1
timestamp 1698431365
transform 1 0 51968 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__372__S1
timestamp 1698431365
transform -1 0 52752 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__376__S
timestamp 1698431365
transform 1 0 47040 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__377__A2
timestamp 1698431365
transform -1 0 30576 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__381__S1
timestamp 1698431365
transform 1 0 26208 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__382__I
timestamp 1698431365
transform 1 0 31136 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__383__I
timestamp 1698431365
transform -1 0 32704 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__385__I1
timestamp 1698431365
transform 1 0 26992 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__385__S
timestamp 1698431365
transform 1 0 28112 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__386__S
timestamp 1698431365
transform 1 0 26768 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__391__S
timestamp 1698431365
transform 1 0 42896 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__392__B
timestamp 1698431365
transform 1 0 39088 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__402__B
timestamp 1698431365
transform 1 0 37856 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__406__I
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__409__S
timestamp 1698431365
transform 1 0 31472 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__420__S
timestamp 1698431365
transform 1 0 50176 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__421__A2
timestamp 1698431365
transform -1 0 31920 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__424__S1
timestamp 1698431365
transform 1 0 27328 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__426__S
timestamp 1698431365
transform -1 0 28896 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__432__B
timestamp 1698431365
transform 1 0 39760 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__442__B
timestamp 1698431365
transform 1 0 35952 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__451__S
timestamp 1698431365
transform -1 0 44016 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__452__S
timestamp 1698431365
transform 1 0 44240 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__454__S0
timestamp 1698431365
transform -1 0 23968 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__455__S0
timestamp 1698431365
transform 1 0 24864 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__470__I
timestamp 1698431365
transform 1 0 23744 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__471__I
timestamp 1698431365
transform 1 0 23296 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__472__I
timestamp 1698431365
transform 1 0 22064 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__473__B
timestamp 1698431365
transform -1 0 21840 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__475__I0
timestamp 1698431365
transform -1 0 24752 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__476__I0
timestamp 1698431365
transform 1 0 28560 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__477__I0
timestamp 1698431365
transform 1 0 30688 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__478__I
timestamp 1698431365
transform -1 0 21504 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__483__I0
timestamp 1698431365
transform 1 0 23184 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__483__I1
timestamp 1698431365
transform 1 0 23184 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__485__I0
timestamp 1698431365
transform -1 0 21952 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__485__I1
timestamp 1698431365
transform 1 0 20160 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__486__I0
timestamp 1698431365
transform -1 0 16352 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__486__I1
timestamp 1698431365
transform 1 0 17024 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__487__I0
timestamp 1698431365
transform 1 0 16576 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__487__I1
timestamp 1698431365
transform 1 0 20160 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__488__I0
timestamp 1698431365
transform 1 0 16352 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__488__I1
timestamp 1698431365
transform -1 0 17696 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__489__I0
timestamp 1698431365
transform 1 0 16800 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__489__I1
timestamp 1698431365
transform 1 0 20608 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__492__A1
timestamp 1698431365
transform -1 0 19936 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__492__A2
timestamp 1698431365
transform -1 0 17808 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__492__A3
timestamp 1698431365
transform 1 0 16800 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__492__A4
timestamp 1698431365
transform 1 0 21504 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__493__I0
timestamp 1698431365
transform -1 0 22288 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__494__I0
timestamp 1698431365
transform -1 0 17024 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__495__I0
timestamp 1698431365
transform 1 0 16352 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__496__CLK
timestamp 1698431365
transform 1 0 26432 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__497__CLK
timestamp 1698431365
transform 1 0 30240 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__498__CLK
timestamp 1698431365
transform 1 0 30576 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__499__CLK
timestamp 1698431365
transform 1 0 29344 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__500__CLK
timestamp 1698431365
transform 1 0 24192 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__501__CLK
timestamp 1698431365
transform 1 0 22848 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__502__CLK
timestamp 1698431365
transform 1 0 20832 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__503__CLK
timestamp 1698431365
transform 1 0 16352 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__504__CLK
timestamp 1698431365
transform 1 0 16128 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__505__CLK
timestamp 1698431365
transform 1 0 16800 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__506__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__507__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__508__CLK
timestamp 1698431365
transform 1 0 9744 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__509__CLK
timestamp 1698431365
transform 1 0 18032 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__510__CLK
timestamp 1698431365
transform 1 0 16352 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__511__CLK
timestamp 1698431365
transform 1 0 15232 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_1_inst_A
timestamp 1698431365
transform 1 0 37968 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_1_inst_B
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_1_inst_CI
timestamp 1698431365
transform 1 0 37520 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_2_inst_A
timestamp 1698431365
transform 1 0 44912 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_2_inst_B
timestamp 1698431365
transform 1 0 44464 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_2_inst_CI
timestamp 1698431365
transform 1 0 44016 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_4_inst_A
timestamp 1698431365
transform 1 0 45360 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_4_inst_B
timestamp 1698431365
transform 1 0 44240 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_4_inst_CI
timestamp 1698431365
transform 1 0 44912 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_1_inst_A
timestamp 1698431365
transform 1 0 57232 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_1_inst_B
timestamp 1698431365
transform 1 0 56784 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_2_inst_A
timestamp 1698431365
transform 1 0 33936 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_2_inst_B
timestamp 1698431365
transform 1 0 34384 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_4_inst_A
timestamp 1698431365
transform 1 0 43568 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_4_inst_B
timestamp 1698431365
transform 1 0 43120 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_1_inst_A1
timestamp 1698431365
transform 1 0 31584 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_1_inst_A2
timestamp 1698431365
transform 1 0 32032 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_2_inst_A1
timestamp 1698431365
transform 1 0 50848 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_2_inst_A2
timestamp 1698431365
transform 1 0 51296 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_4_inst_A1
timestamp 1698431365
transform 1 0 33152 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_4_inst_A2
timestamp 1698431365
transform 1 0 32480 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_1_inst_A1
timestamp 1698431365
transform 1 0 50960 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_1_inst_A2
timestamp 1698431365
transform 1 0 51632 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_1_inst_A3
timestamp 1698431365
transform 1 0 49840 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_2_inst_A1
timestamp 1698431365
transform 1 0 34160 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_2_inst_A2
timestamp 1698431365
transform 1 0 33712 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_2_inst_A3
timestamp 1698431365
transform 1 0 33264 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_4_inst_A1
timestamp 1698431365
transform 1 0 44912 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_4_inst_A2
timestamp 1698431365
transform 1 0 44240 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_4_inst_A3
timestamp 1698431365
transform 1 0 44352 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_1_inst_A1
timestamp 1698431365
transform 1 0 48832 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_1_inst_A2
timestamp 1698431365
transform 1 0 47264 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_1_inst_A3
timestamp 1698431365
transform 1 0 48160 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_1_inst_A4
timestamp 1698431365
transform 1 0 47712 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_2_inst_A1
timestamp 1698431365
transform 1 0 47712 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_2_inst_A2
timestamp 1698431365
transform 1 0 47264 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_2_inst_A3
timestamp 1698431365
transform 1 0 46816 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_2_inst_A4
timestamp 1698431365
transform 1 0 46368 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_4_inst_A1
timestamp 1698431365
transform 1 0 30464 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_4_inst_A2
timestamp 1698431365
transform 1 0 30016 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_4_inst_A3
timestamp 1698431365
transform 1 0 29568 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_4_inst_A4
timestamp 1698431365
transform 1 0 30240 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_1_inst_A1
timestamp 1698431365
transform 1 0 43456 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_1_inst_A2
timestamp 1698431365
transform 1 0 42224 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_1_inst_B
timestamp 1698431365
transform 1 0 41104 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_2_inst_A1
timestamp 1698431365
transform 1 0 57568 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_2_inst_A2
timestamp 1698431365
transform 1 0 57120 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_2_inst_B
timestamp 1698431365
transform 1 0 56672 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_4_inst_A1
timestamp 1698431365
transform 1 0 43008 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_4_inst_A2
timestamp 1698431365
transform 1 0 43904 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_4_inst_B
timestamp 1698431365
transform 1 0 42560 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_1_inst_A1
timestamp 1698431365
transform 1 0 58128 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_1_inst_A2
timestamp 1698431365
transform 1 0 57008 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_1_inst_B1
timestamp 1698431365
transform 1 0 55776 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_1_inst_B2
timestamp 1698431365
transform 1 0 57680 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_2_inst_A1
timestamp 1698431365
transform 1 0 43680 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_2_inst_A2
timestamp 1698431365
transform 1 0 42560 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_2_inst_B1
timestamp 1698431365
transform 1 0 43232 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_2_inst_B2
timestamp 1698431365
transform 1 0 42112 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_4_inst_A1
timestamp 1698431365
transform 1 0 56672 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_4_inst_A2
timestamp 1698431365
transform 1 0 55776 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_4_inst_B1
timestamp 1698431365
transform 1 0 55328 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_4_inst_B2
timestamp 1698431365
transform 1 0 54880 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_1_inst_A1
timestamp 1698431365
transform 1 0 56000 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_1_inst_A2
timestamp 1698431365
transform 1 0 53760 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_1_inst_B
timestamp 1698431365
transform 1 0 55552 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_1_inst_C
timestamp 1698431365
transform 1 0 53312 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_2_inst_A1
timestamp 1698431365
transform 1 0 43568 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_2_inst_A2
timestamp 1698431365
transform 1 0 42336 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_2_inst_B
timestamp 1698431365
transform 1 0 41888 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_2_inst_C
timestamp 1698431365
transform 1 0 42672 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_4_inst_A1
timestamp 1698431365
transform 1 0 40992 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_4_inst_A2
timestamp 1698431365
transform 1 0 39984 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_4_inst_B
timestamp 1698431365
transform 1 0 39872 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_4_inst_C
timestamp 1698431365
transform 1 0 39424 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_1_inst_A1
timestamp 1698431365
transform 1 0 57120 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_1_inst_A2
timestamp 1698431365
transform 1 0 54880 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_1_inst_B1
timestamp 1698431365
transform 1 0 57792 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_1_inst_B2
timestamp 1698431365
transform 1 0 57344 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_1_inst_C
timestamp 1698431365
transform 1 0 56896 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_2_inst_A1
timestamp 1698431365
transform 1 0 43344 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_2_inst_A2
timestamp 1698431365
transform 1 0 40768 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_2_inst_B1
timestamp 1698431365
transform 1 0 40320 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_2_inst_B2
timestamp 1698431365
transform 1 0 39872 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_2_inst_C
timestamp 1698431365
transform 1 0 40208 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_A1
timestamp 1698431365
transform 1 0 51632 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_A2
timestamp 1698431365
transform 1 0 53088 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_B1
timestamp 1698431365
transform 1 0 52080 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_B2
timestamp 1698431365
transform 1 0 53200 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_C
timestamp 1698431365
transform 1 0 52752 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_A1
timestamp 1698431365
transform 1 0 42784 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_A2
timestamp 1698431365
transform 1 0 41664 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_B1
timestamp 1698431365
transform 1 0 39312 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_B2
timestamp 1698431365
transform 1 0 38864 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_C1
timestamp 1698431365
transform 1 0 38416 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_C2
timestamp 1698431365
transform 1 0 37968 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_A1
timestamp 1698431365
transform 1 0 56672 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_A2
timestamp 1698431365
transform 1 0 53648 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_B1
timestamp 1698431365
transform 1 0 53200 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_B2
timestamp 1698431365
transform 1 0 52752 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_C1
timestamp 1698431365
transform 1 0 49280 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_C2
timestamp 1698431365
transform 1 0 50624 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_A1
timestamp 1698431365
transform 1 0 52304 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_A2
timestamp 1698431365
transform 1 0 50064 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_B1
timestamp 1698431365
transform 1 0 52752 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_B2
timestamp 1698431365
transform 1 0 51856 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_C1
timestamp 1698431365
transform -1 0 51632 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_C2
timestamp 1698431365
transform 1 0 50512 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_1_inst_I
timestamp 1698431365
transform 1 0 34720 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_2_inst_I
timestamp 1698431365
transform 1 0 56224 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_3_inst_I
timestamp 1698431365
transform 1 0 34048 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_4_inst_I
timestamp 1698431365
transform 1 0 54992 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_8_inst_I
timestamp 1698431365
transform 1 0 31472 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_12_inst_I
timestamp 1698431365
transform 1 0 45248 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_16_inst_I
timestamp 1698431365
transform 1 0 48832 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_20_inst_I
timestamp 1698431365
transform 1 0 45136 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_1_inst_EN
timestamp 1698431365
transform 1 0 27104 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_1_inst_I
timestamp 1698431365
transform 1 0 26656 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_2_inst_EN
timestamp 1698431365
transform 1 0 29232 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_2_inst_I
timestamp 1698431365
transform 1 0 28560 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_3_inst_EN
timestamp 1698431365
transform 1 0 28560 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_3_inst_I
timestamp 1698431365
transform -1 0 29232 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_4_inst_EN
timestamp 1698431365
transform 1 0 19600 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_4_inst_I
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_8_inst_EN
timestamp 1698431365
transform 1 0 21392 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_8_inst_I
timestamp 1698431365
transform 1 0 21392 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_12_inst_EN
timestamp 1698431365
transform 1 0 24080 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_12_inst_I
timestamp 1698431365
transform 1 0 23632 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_16_inst_EN
timestamp 1698431365
transform 1 0 32032 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_16_inst_I
timestamp 1698431365
transform 1 0 32480 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_1_inst_I
timestamp 1698431365
transform 1 0 21840 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_2_inst_I
timestamp 1698431365
transform 1 0 32144 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_3_inst_I
timestamp 1698431365
transform 1 0 24640 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_4_inst_I
timestamp 1698431365
transform 1 0 23184 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_8_inst_I
timestamp 1698431365
transform 1 0 27440 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_12_inst_I
timestamp 1698431365
transform 1 0 30128 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_16_inst_I
timestamp 1698431365
transform 1 0 19152 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_20_inst_I
timestamp 1698431365
transform 1 0 20272 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_1_inst_I
timestamp 1698431365
transform 1 0 24976 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_2_inst_I
timestamp 1698431365
transform 1 0 28784 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_3_inst_I
timestamp 1698431365
transform 1 0 29232 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_4_inst_I
timestamp 1698431365
transform 1 0 25536 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_8_inst_I
timestamp 1698431365
transform 1 0 28560 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_12_inst_I
timestamp 1698431365
transform 1 0 31248 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_16_inst_I
timestamp 1698431365
transform 1 0 16800 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_20_inst_I
timestamp 1698431365
transform 1 0 16800 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_1_inst_CLKN
timestamp 1698431365
transform 1 0 24528 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_1_inst_D
timestamp 1698431365
transform 1 0 20720 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_2_inst_CLKN
timestamp 1698431365
transform 1 0 43792 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_2_inst_D
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_4_inst_CLKN
timestamp 1698431365
transform 1 0 33488 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_4_inst_D
timestamp 1698431365
transform 1 0 33936 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_CLKN
timestamp 1698431365
transform 1 0 28560 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_D
timestamp 1698431365
transform 1 0 28112 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_RN
timestamp 1698431365
transform 1 0 27664 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_CLKN
timestamp 1698431365
transform 1 0 25760 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_D
timestamp 1698431365
transform 1 0 20720 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_RN
timestamp 1698431365
transform 1 0 20272 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_CLKN
timestamp 1698431365
transform 1 0 21616 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_D
timestamp 1698431365
transform 1 0 21840 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_RN
timestamp 1698431365
transform 1 0 22288 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_CLKN
timestamp 1698431365
transform 1 0 28560 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_D
timestamp 1698431365
transform 1 0 28112 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_RN
timestamp 1698431365
transform 1 0 27664 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 27328 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_CLKN
timestamp 1698431365
transform 1 0 25648 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_D
timestamp 1698431365
transform 1 0 21616 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_RN
timestamp 1698431365
transform 1 0 20272 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 19824 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_CLKN
timestamp 1698431365
transform 1 0 20272 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_D
timestamp 1698431365
transform 1 0 20720 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_RN
timestamp 1698431365
transform 1 0 22512 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 22064 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_CLKN
timestamp 1698431365
transform 1 0 41440 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_D
timestamp 1698431365
transform 1 0 40992 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 40208 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_CLKN
timestamp 1698431365
transform 1 0 31248 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_D
timestamp 1698431365
transform 1 0 30800 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 30352 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_CLKN
timestamp 1698431365
transform 1 0 25648 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_D
timestamp 1698431365
transform 1 0 24640 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 24192 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_1_inst_CLK
timestamp 1698431365
transform 1 0 23408 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_1_inst_D
timestamp 1698431365
transform 1 0 19376 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_2_inst_CLK
timestamp 1698431365
transform 1 0 21392 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_2_inst_D
timestamp 1698431365
transform 1 0 17360 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_4_inst_CLK
timestamp 1698431365
transform 1 0 26432 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_4_inst_D
timestamp 1698431365
transform 1 0 25984 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_1_inst_CLK
timestamp 1698431365
transform 1 0 20720 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_1_inst_D
timestamp 1698431365
transform 1 0 17136 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_1_inst_RN
timestamp 1698431365
transform 1 0 21168 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_2_inst_CLK
timestamp 1698431365
transform 1 0 21840 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_2_inst_D
timestamp 1698431365
transform 1 0 16800 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_2_inst_RN
timestamp 1698431365
transform 1 0 21392 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_4_inst_CLK
timestamp 1698431365
transform 1 0 42000 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_4_inst_D
timestamp 1698431365
transform 1 0 41552 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_4_inst_RN
timestamp 1698431365
transform 1 0 41104 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_CLK
timestamp 1698431365
transform 1 0 31136 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_D
timestamp 1698431365
transform 1 0 31584 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_RN
timestamp 1698431365
transform 1 0 32480 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 32032 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_CLK
timestamp 1698431365
transform 1 0 26320 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_D
timestamp 1698431365
transform 1 0 25872 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_RN
timestamp 1698431365
transform 1 0 25424 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 24640 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_CLK
timestamp 1698431365
transform 1 0 22512 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_D
timestamp 1698431365
transform 1 0 18144 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_RN
timestamp 1698431365
transform 1 0 22960 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 23632 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_1_inst_CLK
timestamp 1698431365
transform 1 0 23968 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_1_inst_D
timestamp 1698431365
transform 1 0 19040 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 23520 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_2_inst_CLK
timestamp 1698431365
transform 1 0 27216 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_2_inst_D
timestamp 1698431365
transform 1 0 27216 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 26880 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_4_inst_CLK
timestamp 1698431365
transform 1 0 22064 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_4_inst_D
timestamp 1698431365
transform 1 0 17472 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 22624 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlya_1_inst_I
timestamp 1698431365
transform 1 0 38640 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlya_2_inst_I
timestamp 1698431365
transform 1 0 38192 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlya_4_inst_I
timestamp 1698431365
transform 1 0 31696 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyb_1_inst_I
timestamp 1698431365
transform 1 0 24192 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyb_2_inst_I
timestamp 1698431365
transform 1 0 22960 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyb_4_inst_I
timestamp 1698431365
transform 1 0 28672 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyc_1_inst_I
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyc_2_inst_I
timestamp 1698431365
transform 1 0 20720 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyc_4_inst_I
timestamp 1698431365
transform 1 0 41440 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyd_1_inst_I
timestamp 1698431365
transform 1 0 35504 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyd_2_inst_I
timestamp 1698431365
transform 1 0 30912 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyd_4_inst_I
timestamp 1698431365
transform 1 0 24640 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_1_inst_CLKN
timestamp 1698431365
transform 1 0 25872 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_1_inst_E
timestamp 1698431365
transform 1 0 20272 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_1_inst_TE
timestamp 1698431365
transform 1 0 19824 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_2_inst_CLKN
timestamp 1698431365
transform 1 0 24640 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_2_inst_E
timestamp 1698431365
transform 1 0 24192 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_2_inst_TE
timestamp 1698431365
transform 1 0 23744 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_4_inst_CLKN
timestamp 1698431365
transform 1 0 23520 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_4_inst_E
timestamp 1698431365
transform 1 0 23072 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_4_inst_TE
timestamp 1698431365
transform 1 0 23072 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_2_inst_CLK
timestamp 1698431365
transform 1 0 24640 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_2_inst_E
timestamp 1698431365
transform 1 0 24192 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_2_inst_TE
timestamp 1698431365
transform 1 0 24080 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_4_inst_CLK
timestamp 1698431365
transform 1 0 28672 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_4_inst_E
timestamp 1698431365
transform 1 0 28224 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_4_inst_TE
timestamp 1698431365
transform 1 0 27776 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_1_inst_I
timestamp 1698431365
transform 1 0 33152 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_2_inst_I
timestamp 1698431365
transform 1 0 56896 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_3_inst_I
timestamp 1698431365
transform 1 0 35504 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_4_inst_I
timestamp 1698431365
transform 1 0 56672 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_8_inst_I
timestamp 1698431365
transform 1 0 31024 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_12_inst_I
timestamp 1698431365
transform 1 0 45696 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_16_inst_I
timestamp 1698431365
transform 1 0 46368 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_20_inst_I
timestamp 1698431365
transform 1 0 47040 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_1_inst_EN
timestamp 1698431365
transform 1 0 34160 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_1_inst_I
timestamp 1698431365
transform 1 0 34048 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_2_inst_EN
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_2_inst_I
timestamp 1698431365
transform 1 0 24640 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_3_inst_EN
timestamp 1698431365
transform 1 0 21280 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_3_inst_I
timestamp 1698431365
transform 1 0 20832 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_4_inst_EN
timestamp 1698431365
transform 1 0 22064 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_4_inst_I
timestamp 1698431365
transform -1 0 19376 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_8_inst_EN
timestamp 1698431365
transform 1 0 24640 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_8_inst_I
timestamp 1698431365
transform 1 0 20720 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_12_inst_EN
timestamp 1698431365
transform 1 0 23408 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_12_inst_I
timestamp 1698431365
transform 1 0 23632 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_1_inst_D
timestamp 1698431365
transform 1 0 45360 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_1_inst_E
timestamp 1698431365
transform 1 0 45360 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_2_inst_D
timestamp 1698431365
transform 1 0 36624 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_2_inst_E
timestamp 1698431365
transform 1 0 37632 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_4_inst_D
timestamp 1698431365
transform 1 0 47712 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_4_inst_E
timestamp 1698431365
transform 1 0 48160 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_1_inst_D
timestamp 1698431365
transform 1 0 36176 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_1_inst_E
timestamp 1698431365
transform 1 0 37072 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_1_inst_RN
timestamp 1698431365
transform 1 0 36624 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_2_inst_D
timestamp 1698431365
transform 1 0 49280 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_2_inst_E
timestamp 1698431365
transform 1 0 50176 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_2_inst_RN
timestamp 1698431365
transform 1 0 49728 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_4_inst_D
timestamp 1698431365
transform 1 0 44464 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_4_inst_E
timestamp 1698431365
transform 1 0 43568 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_4_inst_RN
timestamp 1698431365
transform 1 0 44016 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_D
timestamp 1698431365
transform 1 0 37072 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_E
timestamp 1698431365
transform 1 0 36400 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_RN
timestamp 1698431365
transform 1 0 36400 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 35952 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_D
timestamp 1698431365
transform 1 0 29568 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_E
timestamp 1698431365
transform 1 0 29120 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_RN
timestamp 1698431365
transform 1 0 28672 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 28224 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_D
timestamp 1698431365
transform 1 0 22064 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_E
timestamp 1698431365
transform 1 0 22736 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_RN
timestamp 1698431365
transform 1 0 21616 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 22288 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_1_inst_D
timestamp 1698431365
transform 1 0 24192 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_1_inst_E
timestamp 1698431365
transform 1 0 23744 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 23296 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_2_inst_D
timestamp 1698431365
transform 1 0 33488 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_2_inst_E
timestamp 1698431365
transform 1 0 33040 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 32032 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_4_inst_D
timestamp 1698431365
transform 1 0 26096 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_4_inst_E
timestamp 1698431365
transform 1 0 24640 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 24192 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_1_inst_I0
timestamp 1698431365
transform 1 0 50624 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_1_inst_I1
timestamp 1698431365
transform 1 0 50736 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_1_inst_S
timestamp 1698431365
transform 1 0 50288 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_2_inst_I0
timestamp 1698431365
transform 1 0 37072 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_2_inst_I1
timestamp 1698431365
transform 1 0 36400 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_2_inst_S
timestamp 1698431365
transform 1 0 37072 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_4_inst_I0
timestamp 1698431365
transform 1 0 52304 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_4_inst_I1
timestamp 1698431365
transform 1 0 51408 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_4_inst_S
timestamp 1698431365
transform 1 0 51856 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_I0
timestamp 1698431365
transform 1 0 56672 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_I1
timestamp 1698431365
transform 1 0 52080 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_I2
timestamp 1698431365
transform 1 0 51184 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_I3
timestamp 1698431365
transform 1 0 51632 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_S0
timestamp 1698431365
transform 1 0 50512 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_S1
timestamp 1698431365
transform 1 0 50960 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_I0
timestamp 1698431365
transform 1 0 39424 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_I1
timestamp 1698431365
transform 1 0 38976 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_I2
timestamp 1698431365
transform 1 0 38528 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_I3
timestamp 1698431365
transform 1 0 38080 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_S0
timestamp 1698431365
transform -1 0 37856 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_S1
timestamp 1698431365
transform -1 0 37408 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_I0
timestamp 1698431365
transform 1 0 35504 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_I1
timestamp 1698431365
transform 1 0 35280 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_I2
timestamp 1698431365
transform 1 0 35056 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_I3
timestamp 1698431365
transform 1 0 34832 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_S0
timestamp 1698431365
transform 1 0 34608 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_S1
timestamp 1698431365
transform 1 0 33376 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_1_inst_A1
timestamp 1698431365
transform 1 0 56448 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_1_inst_A2
timestamp 1698431365
transform 1 0 56000 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_2_inst_A1
timestamp 1698431365
transform 1 0 38416 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_2_inst_A2
timestamp 1698431365
transform 1 0 38304 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_4_inst_A1
timestamp 1698431365
transform 1 0 50064 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_4_inst_A2
timestamp 1698431365
transform 1 0 50512 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_1_inst_A1
timestamp 1698431365
transform 1 0 32928 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_1_inst_A2
timestamp 1698431365
transform 1 0 34048 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_1_inst_A3
timestamp 1698431365
transform 1 0 33152 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_2_inst_A1
timestamp 1698431365
transform 1 0 46368 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_2_inst_A2
timestamp 1698431365
transform 1 0 44688 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_2_inst_A3
timestamp 1698431365
transform 1 0 45136 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_4_inst_A1
timestamp 1698431365
transform 1 0 48160 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_4_inst_A2
timestamp 1698431365
transform 1 0 47712 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_4_inst_A3
timestamp 1698431365
transform 1 0 47600 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_1_inst_A1
timestamp 1698431365
transform 1 0 41440 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_1_inst_A2
timestamp 1698431365
transform 1 0 40992 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_1_inst_A3
timestamp 1698431365
transform 1 0 40320 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_1_inst_A4
timestamp 1698431365
transform 1 0 40096 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_2_inst_A1
timestamp 1698431365
transform 1 0 48944 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_2_inst_A2
timestamp 1698431365
transform 1 0 45584 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_2_inst_A3
timestamp 1698431365
transform 1 0 46032 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_2_inst_A4
timestamp 1698431365
transform 1 0 46368 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_4_inst_A1
timestamp 1698431365
transform 1 0 56672 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_4_inst_A2
timestamp 1698431365
transform 1 0 53200 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_4_inst_A3
timestamp 1698431365
transform 1 0 52080 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_4_inst_A4
timestamp 1698431365
transform 1 0 52752 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_1_inst_A1
timestamp 1698431365
transform 1 0 48832 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_1_inst_A2
timestamp 1698431365
transform 1 0 48160 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_2_inst_A1
timestamp 1698431365
transform 1 0 56560 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_2_inst_A2
timestamp 1698431365
transform 1 0 56112 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_4_inst_A1
timestamp 1698431365
transform 1 0 40320 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_4_inst_A2
timestamp 1698431365
transform 1 0 40992 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_1_inst_A1
timestamp 1698431365
transform 1 0 57120 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_1_inst_A2
timestamp 1698431365
transform 1 0 57120 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_1_inst_A3
timestamp 1698431365
transform 1 0 56672 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_2_inst_A1
timestamp 1698431365
transform 1 0 48384 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_2_inst_A2
timestamp 1698431365
transform 1 0 47264 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_2_inst_A3
timestamp 1698431365
transform 1 0 47712 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_4_inst_A1
timestamp 1698431365
transform 1 0 38304 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_4_inst_A2
timestamp 1698431365
transform 1 0 39200 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_4_inst_A3
timestamp 1698431365
transform 1 0 38752 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_1_inst_A1
timestamp 1698431365
transform 1 0 46256 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_1_inst_A2
timestamp 1698431365
transform 1 0 47152 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_1_inst_A3
timestamp 1698431365
transform 1 0 45808 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_1_inst_A4
timestamp 1698431365
transform 1 0 46704 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_2_inst_A1
timestamp 1698431365
transform 1 0 53424 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_2_inst_A2
timestamp 1698431365
transform 1 0 55328 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_2_inst_A3
timestamp 1698431365
transform 1 0 52976 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_2_inst_A4
timestamp 1698431365
transform 1 0 53648 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_4_inst_A1
timestamp 1698431365
transform 1 0 45920 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_4_inst_A2
timestamp 1698431365
transform 1 0 45472 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_4_inst_A3
timestamp 1698431365
transform 1 0 45024 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_4_inst_A4
timestamp 1698431365
transform 1 0 44352 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_1_inst_A1
timestamp 1698431365
transform 1 0 46592 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_1_inst_A2
timestamp 1698431365
transform 1 0 46144 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_1_inst_B
timestamp 1698431365
transform 1 0 44912 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_2_inst_A1
timestamp 1698431365
transform 1 0 31584 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_2_inst_A2
timestamp 1698431365
transform 1 0 32032 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_2_inst_B
timestamp 1698431365
transform 1 0 34496 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_4_inst_A1
timestamp 1698431365
transform 1 0 51520 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_4_inst_A2
timestamp 1698431365
transform 1 0 51072 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_4_inst_B
timestamp 1698431365
transform 1 0 50400 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_1_inst_A1
timestamp 1698431365
transform 1 0 39312 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_1_inst_A2
timestamp 1698431365
transform 1 0 40096 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_1_inst_B1
timestamp 1698431365
transform 1 0 30688 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_1_inst_B2
timestamp 1698431365
transform 1 0 35056 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_2_inst_A1
timestamp 1698431365
transform 1 0 52304 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_2_inst_A2
timestamp 1698431365
transform 1 0 50176 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_2_inst_B1
timestamp 1698431365
transform 1 0 53872 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_2_inst_B2
timestamp 1698431365
transform 1 0 51520 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_4_inst_A1
timestamp 1698431365
transform 1 0 32032 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_4_inst_A2
timestamp 1698431365
transform 1 0 32480 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_4_inst_B1
timestamp 1698431365
transform 1 0 33600 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_4_inst_B2
timestamp 1698431365
transform 1 0 33152 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_1_inst_A1
timestamp 1698431365
transform 1 0 49728 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_1_inst_A2
timestamp 1698431365
transform 1 0 50176 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_1_inst_A3
timestamp 1698431365
transform 1 0 51072 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_1_inst_B
timestamp 1698431365
transform 1 0 50624 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_2_inst_A1
timestamp 1698431365
transform 1 0 49616 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_2_inst_A2
timestamp 1698431365
transform 1 0 50960 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_2_inst_A3
timestamp 1698431365
transform 1 0 50064 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_2_inst_B
timestamp 1698431365
transform 1 0 51408 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_4_inst_A1
timestamp 1698431365
transform 1 0 42560 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_4_inst_A2
timestamp 1698431365
transform 1 0 43232 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_4_inst_A3
timestamp 1698431365
transform 1 0 42784 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_4_inst_B
timestamp 1698431365
transform 1 0 40320 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_1_inst_A1
timestamp 1698431365
transform 1 0 35952 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_1_inst_A2
timestamp 1698431365
transform 1 0 35504 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_1_inst_A3
timestamp 1698431365
transform 1 0 35056 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_1_inst_B1
timestamp 1698431365
transform 1 0 34608 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_1_inst_B2
timestamp 1698431365
transform 1 0 34160 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_2_inst_A1
timestamp 1698431365
transform 1 0 48944 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_2_inst_A2
timestamp 1698431365
transform 1 0 56448 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_2_inst_A3
timestamp 1698431365
transform 1 0 52304 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_2_inst_B1
timestamp 1698431365
transform 1 0 50176 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_2_inst_B2
timestamp 1698431365
transform 1 0 51968 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_4_inst_A1
timestamp 1698431365
transform 1 0 35392 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_4_inst_A2
timestamp 1698431365
transform 1 0 34944 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_4_inst_A3
timestamp 1698431365
transform 1 0 34496 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_4_inst_B1
timestamp 1698431365
transform 1 0 34048 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_4_inst_B2
timestamp 1698431365
transform 1 0 33152 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_A1
timestamp 1698431365
transform 1 0 51184 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_A2
timestamp 1698431365
transform 1 0 51072 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_A3
timestamp 1698431365
transform 1 0 50736 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_B1
timestamp 1698431365
transform 1 0 50288 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_B2
timestamp 1698431365
transform 1 0 50624 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_B3
timestamp 1698431365
transform 1 0 50176 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_A1
timestamp 1698431365
transform 1 0 38304 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_A2
timestamp 1698431365
transform 1 0 37072 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_A3
timestamp 1698431365
transform 1 0 37856 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_B1
timestamp 1698431365
transform 1 0 36288 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_B2
timestamp 1698431365
transform 1 0 35840 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_B3
timestamp 1698431365
transform 1 0 36400 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_A1
timestamp 1698431365
transform 1 0 50176 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_A2
timestamp 1698431365
transform 1 0 48832 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_A3
timestamp 1698431365
transform 1 0 48832 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_B1
timestamp 1698431365
transform 1 0 49728 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_B2
timestamp 1698431365
transform 1 0 48048 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_B3
timestamp 1698431365
transform 1 0 47600 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_1_inst_A1
timestamp 1698431365
transform 1 0 57456 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_1_inst_A2
timestamp 1698431365
transform 1 0 57008 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_1_inst_B
timestamp 1698431365
transform 1 0 56560 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_1_inst_C
timestamp 1698431365
transform 1 0 56112 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_2_inst_A1
timestamp 1698431365
transform 1 0 43120 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_2_inst_A2
timestamp 1698431365
transform 1 0 41888 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_2_inst_B
timestamp 1698431365
transform 1 0 40992 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_2_inst_C
timestamp 1698431365
transform 1 0 41440 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_4_inst_A1
timestamp 1698431365
transform 1 0 37072 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_4_inst_A2
timestamp 1698431365
transform 1 0 36400 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_4_inst_B
timestamp 1698431365
transform 1 0 36400 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_4_inst_C
timestamp 1698431365
transform 1 0 35952 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_1_inst_A1
timestamp 1698431365
transform 1 0 51184 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_1_inst_A2
timestamp 1698431365
transform 1 0 49840 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_1_inst_B1
timestamp 1698431365
transform 1 0 49392 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_1_inst_B2
timestamp 1698431365
transform 1 0 49168 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_1_inst_C
timestamp 1698431365
transform 1 0 48160 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_2_inst_A1
timestamp 1698431365
transform 1 0 42672 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_2_inst_A2
timestamp 1698431365
transform 1 0 42224 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_2_inst_B1
timestamp 1698431365
transform 1 0 41776 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_2_inst_B2
timestamp 1698431365
transform 1 0 41328 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_2_inst_C
timestamp 1698431365
transform 1 0 41664 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_4_inst_A1
timestamp 1698431365
transform 1 0 55776 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_4_inst_A2
timestamp 1698431365
transform 1 0 54656 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_4_inst_B1
timestamp 1698431365
transform 1 0 54208 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_4_inst_B2
timestamp 1698431365
transform 1 0 53200 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_4_inst_C
timestamp 1698431365
transform 1 0 52752 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_A1
timestamp 1698431365
transform 1 0 41888 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_A2
timestamp 1698431365
transform 1 0 40656 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_B1
timestamp 1698431365
transform 1 0 41440 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_B2
timestamp 1698431365
transform 1 0 40992 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_C1
timestamp 1698431365
transform 1 0 40208 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_C2
timestamp 1698431365
transform 1 0 39760 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_A1
timestamp 1698431365
transform 1 0 51184 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_A2
timestamp 1698431365
transform 1 0 52304 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_B1
timestamp 1698431365
transform 1 0 51408 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_B2
timestamp 1698431365
transform 1 0 51632 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_C1
timestamp 1698431365
transform 1 0 52080 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_C2
timestamp 1698431365
transform 1 0 51856 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_A1
timestamp 1698431365
transform 1 0 50512 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_A2
timestamp 1698431365
transform 1 0 52304 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_B1
timestamp 1698431365
transform 1 0 51856 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_B2
timestamp 1698431365
transform 1 0 50960 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_C1
timestamp 1698431365
transform 1 0 51408 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_C2
timestamp 1698431365
transform 1 0 50736 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_1_inst_A1
timestamp 1698431365
transform 1 0 55664 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_1_inst_A2
timestamp 1698431365
transform 1 0 54320 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_2_inst_A1
timestamp 1698431365
transform 1 0 41664 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_2_inst_A2
timestamp 1698431365
transform 1 0 40432 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_4_inst_A1
timestamp 1698431365
transform 1 0 57120 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_4_inst_A2
timestamp 1698431365
transform 1 0 56672 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_1_inst_A1
timestamp 1698431365
transform 1 0 45024 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_1_inst_A2
timestamp 1698431365
transform 1 0 45920 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_1_inst_A3
timestamp 1698431365
transform 1 0 45472 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_2_inst_A1
timestamp 1698431365
transform 1 0 36960 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_2_inst_A2
timestamp 1698431365
transform 1 0 37520 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_2_inst_A3
timestamp 1698431365
transform 1 0 37072 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_4_inst_A1
timestamp 1698431365
transform 1 0 43456 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_4_inst_A2
timestamp 1698431365
transform 1 0 42112 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_4_inst_A3
timestamp 1698431365
transform 1 0 43008 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_1_inst_A1
timestamp 1698431365
transform 1 0 50624 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_1_inst_A2
timestamp 1698431365
transform 1 0 50176 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_1_inst_A3
timestamp 1698431365
transform 1 0 48160 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_1_inst_A4
timestamp 1698431365
transform 1 0 49728 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_2_inst_A1
timestamp 1698431365
transform 1 0 45360 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_2_inst_A2
timestamp 1698431365
transform 1 0 44912 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_2_inst_A3
timestamp 1698431365
transform 1 0 44016 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_2_inst_A4
timestamp 1698431365
transform 1 0 43792 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_4_inst_A1
timestamp 1698431365
transform 1 0 49840 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_4_inst_A2
timestamp 1698431365
transform 1 0 49392 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_4_inst_A3
timestamp 1698431365
transform 1 0 49392 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_4_inst_A4
timestamp 1698431365
transform 1 0 48944 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_1_inst_CLK
timestamp 1698431365
transform 1 0 22736 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_1_inst_D
timestamp 1698431365
transform 1 0 16800 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_1_inst_SE
timestamp 1698431365
transform 1 0 23408 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_1_inst_SI
timestamp 1698431365
transform 1 0 22960 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_2_inst_CLK
timestamp 1698431365
transform 1 0 42112 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_2_inst_D
timestamp 1698431365
transform 1 0 41664 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_2_inst_SE
timestamp 1698431365
transform 1 0 41216 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_2_inst_SI
timestamp 1698431365
transform 1 0 39424 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_4_inst_CLK
timestamp 1698431365
transform 1 0 35952 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_4_inst_D
timestamp 1698431365
transform 1 0 37296 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_4_inst_SE
timestamp 1698431365
transform 1 0 36400 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_4_inst_SI
timestamp 1698431365
transform 1 0 37744 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_CLK
timestamp 1698431365
transform 1 0 33600 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_D
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_RN
timestamp 1698431365
transform 1 0 32256 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_SE
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_SI
timestamp 1698431365
transform 1 0 30912 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_CLK
timestamp 1698431365
transform 1 0 23856 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_D
timestamp 1698431365
transform 1 0 22960 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_RN
timestamp 1698431365
transform 1 0 22512 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SE
timestamp 1698431365
transform 1 0 23184 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SI
timestamp 1698431365
transform 1 0 22064 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_CLK
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_D
timestamp 1698431365
transform 1 0 20048 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_RN
timestamp 1698431365
transform 1 0 19152 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_SE
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_SI
timestamp 1698431365
transform 1 0 25312 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_CLK
timestamp 1698431365
transform 1 0 28560 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_D
timestamp 1698431365
transform 1 0 28112 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_RN
timestamp 1698431365
transform 1 0 27664 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SETN
timestamp 1698431365
transform -1 0 28112 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SE
timestamp 1698431365
transform 1 0 27216 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SI
timestamp 1698431365
transform 1 0 26768 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_CLK
timestamp 1698431365
transform 1 0 27104 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_D
timestamp 1698431365
transform 1 0 20720 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_RN
timestamp 1698431365
transform 1 0 20272 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SE
timestamp 1698431365
transform 1 0 19824 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 20608 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SI
timestamp 1698431365
transform 1 0 20384 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_CLK
timestamp 1698431365
transform 1 0 26432 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_D
timestamp 1698431365
transform 1 0 17808 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_RN
timestamp 1698431365
transform 1 0 26320 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 25536 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SE
timestamp 1698431365
transform 1 0 25984 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SI
timestamp 1698431365
transform 1 0 25536 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_CLK
timestamp 1698431365
transform 1 0 40992 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_D
timestamp 1698431365
transform 1 0 41552 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SE
timestamp 1698431365
transform 1 0 40320 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 39872 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SI
timestamp 1698431365
transform 1 0 39088 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_CLK
timestamp 1698431365
transform 1 0 37296 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_D
timestamp 1698431365
transform 1 0 35056 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 35952 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SE
timestamp 1698431365
transform 1 0 35504 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SI
timestamp 1698431365
transform 1 0 36400 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_CLK
timestamp 1698431365
transform 1 0 30576 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_D
timestamp 1698431365
transform 1 0 31024 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 31472 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SE
timestamp 1698431365
transform 1 0 30128 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SI
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_1_inst_A1
timestamp 1698431365
transform 1 0 37072 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_1_inst_A2
timestamp 1698431365
transform 1 0 37520 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_2_inst_A1
timestamp 1698431365
transform 1 0 49504 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_2_inst_A2
timestamp 1698431365
transform 1 0 49952 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_4_inst_A1
timestamp 1698431365
transform 1 0 46032 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_4_inst_A2
timestamp 1698431365
transform 1 0 45584 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_1_inst_A1
timestamp 1698431365
transform 1 0 37968 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_1_inst_A2
timestamp 1698431365
transform 1 0 37520 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_1_inst_A3
timestamp 1698431365
transform 1 0 37072 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_2_inst_A1
timestamp 1698431365
transform 1 0 42560 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_2_inst_A2
timestamp 1698431365
transform 1 0 39872 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_2_inst_A3
timestamp 1698431365
transform 1 0 40320 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_4_inst_A1
timestamp 1698431365
transform 1 0 49056 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_4_inst_A2
timestamp 1698431365
transform 1 0 48608 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_4_inst_A3
timestamp 1698431365
transform 1 0 48160 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_1_inst_A1
timestamp 1698431365
transform 1 0 44240 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_1_inst_A2
timestamp 1698431365
transform 1 0 44688 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_2_inst_A1
timestamp 1698431365
transform 1 0 51968 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_2_inst_A2
timestamp 1698431365
transform 1 0 51184 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_4_inst_A1
timestamp 1698431365
transform 1 0 37968 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_4_inst_A2
timestamp 1698431365
transform 1 0 37744 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_1_inst_A1
timestamp 1698431365
transform 1 0 50400 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_1_inst_A2
timestamp 1698431365
transform 1 0 49952 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_1_inst_A3
timestamp 1698431365
transform 1 0 49504 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_2_inst_A1
timestamp 1698431365
transform 1 0 53088 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_2_inst_A2
timestamp 1698431365
transform 1 0 50960 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_2_inst_A3
timestamp 1698431365
transform 1 0 52752 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_4_inst_A1
timestamp 1698431365
transform 1 0 43568 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_4_inst_A2
timestamp 1698431365
transform 1 0 43120 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_4_inst_A3
timestamp 1698431365
transform 1 0 39872 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[1\].div_flop_RN
timestamp 1698431365
transform 1 0 11200 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[2\].div_flop_RN
timestamp 1698431365
transform 1 0 10528 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[3\].div_flop_RN
timestamp 1698431365
transform 1 0 14000 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[4\].div_flop_RN
timestamp 1698431365
transform 1 0 9296 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[5\].div_flop_RN
timestamp 1698431365
transform 1 0 9632 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[6\].div_flop_RN
timestamp 1698431365
transform 1 0 5712 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[7\].div_flop_RN
timestamp 1698431365
transform 1 0 6160 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[8\].div_flop_RN
timestamp 1698431365
transform 1 0 2688 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[9\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[10\].div_flop_RN
timestamp 1698431365
transform 1 0 2240 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[11\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[12\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[13\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[14\].div_flop_RN
timestamp 1698431365
transform 1 0 2240 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[15\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[16\].div_flop_RN
timestamp 1698431365
transform 1 0 7280 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[17\].div_flop_RN
timestamp 1698431365
transform 1 0 2800 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[18\].div_flop_RN
timestamp 1698431365
transform 1 0 3360 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[19\].div_flop_RN
timestamp 1698431365
transform 1 0 3248 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[20\].div_flop_RN
timestamp 1698431365
transform 1 0 3024 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[21\].div_flop_RN
timestamp 1698431365
transform 1 0 2240 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[22\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[23\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[24\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[25\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[26\].div_flop_RN
timestamp 1698431365
transform 1 0 3696 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[27\].div_flop_RN
timestamp 1698431365
transform 1 0 6608 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[28\].div_flop_RN
timestamp 1698431365
transform 1 0 7168 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[29\].div_flop_RN
timestamp 1698431365
transform 1 0 8624 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[30\].div_flop_RN
timestamp 1698431365
transform 1 0 8848 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[31\].div_flop_RN
timestamp 1698431365
transform 1 0 9296 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[32\].div_flop_RN
timestamp 1698431365
transform 1 0 9856 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[33\].div_flop_RN
timestamp 1698431365
transform 1 0 9296 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[34\].div_flop_RN
timestamp 1698431365
transform 1 0 10976 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.slow_clock_inv_I
timestamp 1698431365
transform 1 0 8512 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__addf_1  cm_inst.cc_inst.addf_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37184 0 -1 42336
box -86 -90 3446 1098
use gf180mcu_fd_sc_mcu9t5v0__addf_2  cm_inst.cc_inst.addf_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 38304
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__addf_4  cm_inst.cc_inst.addf_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 36288
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__addh_1  cm_inst.cc_inst.addh_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 56560 0 1 20160
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__addh_2  cm_inst.cc_inst.addh_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 37184 0 -1 42336
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__addh_4  cm_inst.cc_inst.addh_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 47152 0 -1 38304
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  cm_inst.cc_inst.and2_1_inst
timestamp 1698431365
transform -1 0 33824 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_2  cm_inst.cc_inst.and2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 51744 0 -1 40320
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_4  cm_inst.cc_inst.and2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 34048 0 -1 28224
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__and3_1  cm_inst.cc_inst.and3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 51184 0 1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__and3_2  cm_inst.cc_inst.and3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 33936 0 -1 26208
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__and3_4  cm_inst.cc_inst.and3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 46928 0 -1 24192
box -86 -90 2326 1098
use gf180mcu_fd_sc_mcu9t5v0__and4_1  cm_inst.cc_inst.and4_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 49840 0 -1 16128
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__and4_2  cm_inst.cc_inst.and4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 46928 0 -1 44352
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__and4_4  cm_inst.cc_inst.and4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 30688 0 1 26208
box -86 -90 2774 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_1  cm_inst.cc_inst.aoi21_1_inst
timestamp 1698431365
transform 1 0 41440 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_2  cm_inst.cc_inst.aoi21_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 54768 0 -1 42336
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_4  cm_inst.cc_inst.aoi21_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 43680 0 -1 24192
box -86 -90 2774 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  cm_inst.cc_inst.aoi22_1_inst
timestamp 1698431365
transform -1 0 57456 0 -1 32256
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_2  cm_inst.cc_inst.aoi22_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 42560 0 -1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_4  cm_inst.cc_inst.aoi22_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 57344 0 1 24192
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  cm_inst.cc_inst.aoi211_1_inst
timestamp 1698431365
transform 1 0 54208 0 -1 14112
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_2  cm_inst.cc_inst.aoi211_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 44464 0 1 44352
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_4  cm_inst.cc_inst.aoi211_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40320 0 1 24192
box -86 -90 4118 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi221_1  cm_inst.cc_inst.aoi221_1_inst
timestamp 1698431365
transform -1 0 56224 0 1 42336
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi221_2  cm_inst.cc_inst.aoi221_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 43120 0 -1 26208
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi221_4  cm_inst.cc_inst.aoi221_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 58016 0 1 30240
box -86 -90 4566 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi222_1  cm_inst.cc_inst.aoi222_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38976 0 -1 28224
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi222_2  cm_inst.cc_inst.aoi222_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 53312 0 -1 28224
box -86 -90 2886 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi222_4  cm_inst.cc_inst.aoi222_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -90 5350 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  cm_inst.cc_inst.buf_1_inst
timestamp 1698431365
transform -1 0 35280 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_2  cm_inst.cc_inst.buf_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 57344 0 -1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_3  cm_inst.cc_inst.buf_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 33936 0 1 34272
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_4  cm_inst.cc_inst.buf_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 56784 0 1 32256
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_8  cm_inst.cc_inst.buf_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 34608 0 1 36288
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_12  cm_inst.cc_inst.buf_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 50176 0 1 24192
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_16  cm_inst.cc_inst.buf_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 54208 0 -1 14112
box -86 -90 5686 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_20  cm_inst.cc_inst.buf_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 45360 0 1 46368
box -86 -90 7030 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_1  cm_inst.cc_inst.bufz_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 27328 0 1 14112
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_2  cm_inst.cc_inst.bufz_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 16128
box -86 -90 1766 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_3  cm_inst.cc_inst.bufz_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 30912 0 -1 16128
box -86 -90 2214 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_4  cm_inst.cc_inst.bufz_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_8  cm_inst.cc_inst.bufz_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 12096
box -86 -90 3782 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_12  cm_inst.cc_inst.bufz_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 -1 16128
box -86 -90 5126 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_16  cm_inst.cc_inst.bufz_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 39312 0 -1 48384
box -86 -90 6470 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  cm_inst.cc_inst.clkbuf_1_inst
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_2  cm_inst.cc_inst.clkbuf_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 31920 0 -1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_3  cm_inst.cc_inst.clkbuf_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 26656 0 -1 40320
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_4  cm_inst.cc_inst.clkbuf_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 20944 0 -1 22176
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_8  cm_inst.cc_inst.clkbuf_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 -1 20160
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_12  cm_inst.cc_inst.clkbuf_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 30352 0 1 38304
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_16  cm_inst.cc_inst.clkbuf_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 20160
box -86 -90 5686 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_20  cm_inst.cc_inst.clkbuf_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 18144
box -86 -90 7030 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  cm_inst.cc_inst.clkinv_1_inst
timestamp 1698431365
transform 1 0 25200 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_2  cm_inst.cc_inst.clkinv_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 29680 0 1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_3  cm_inst.cc_inst.clkinv_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 28672 0 1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_4  cm_inst.cc_inst.clkinv_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 26656 0 -1 26208
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_8  cm_inst.cc_inst.clkinv_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 20160
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_12  cm_inst.cc_inst.clkinv_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 34384 0 1 40320
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_16  cm_inst.cc_inst.clkinv_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 16576 0 -1 22176
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_20  cm_inst.cc_inst.clkinv_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 20160
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnq_1  cm_inst.cc_inst.dffnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 24192
box -86 -90 3446 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnq_2  cm_inst.cc_inst.dffnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnq_4  cm_inst.cc_inst.dffnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 34384 0 -1 10080
box -86 -90 4006 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1  cm_inst.cc_inst.dffnrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2  cm_inst.cc_inst.dffnrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 1 10080
box -86 -90 4006 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4  cm_inst.cc_inst.dffnrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 1 46368
box -86 -90 4454 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1  cm_inst.cc_inst.dffnrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29232 0 1 46368
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2  cm_inst.cc_inst.dffnrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 44352
box -86 -90 4566 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4  cm_inst.cc_inst.dffnrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 16016 0 1 24192
box -86 -90 5014 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1  cm_inst.cc_inst.dffnsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40880 0 -1 14112
box -86 -90 4118 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2  cm_inst.cc_inst.dffnsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 31472 0 1 10080
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4  cm_inst.cc_inst.dffnsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 25872 0 -1 10080
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  cm_inst.cc_inst.dffq_1_inst
timestamp 1698431365
transform 1 0 19600 0 -1 12096
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_2  cm_inst.cc_inst.dffq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 1 46368
box -86 -90 3446 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_4  cm_inst.cc_inst.dffq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 27552 0 -1 48384
box -86 -90 4006 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  cm_inst.cc_inst.dffrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17360 0 1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_2  cm_inst.cc_inst.dffrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 26208
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_4  cm_inst.cc_inst.dffrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 41776 0 -1 12096
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1  cm_inst.cc_inst.dffrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 12096
box -86 -90 4230 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2  cm_inst.cc_inst.dffrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 26544 0 -1 12096
box -86 -90 4454 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4  cm_inst.cc_inst.dffrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 18368 0 -1 10080
box -86 -90 4902 1098
use gf180mcu_fd_sc_mcu9t5v0__dffsnq_1  cm_inst.cc_inst.dffsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 19264 0 -1 48384
box -86 -90 4118 1098
use gf180mcu_fd_sc_mcu9t5v0__dffsnq_2  cm_inst.cc_inst.dffsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 -1 46368
box -86 -90 4230 1098
use gf180mcu_fd_sc_mcu9t5v0__dffsnq_4  cm_inst.cc_inst.dffsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 -1 46368
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__dlya_1  cm_inst.cc_inst.dlya_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 39984 0 1 18144
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__dlya_2  cm_inst.cc_inst.dlya_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38752 0 -1 14112
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__dlya_4  cm_inst.cc_inst.dlya_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 31920 0 1 18144
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyb_1  cm_inst.cc_inst.dlyb_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 25200 0 -1 18144
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyb_2  cm_inst.cc_inst.dlyb_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 12096
box -86 -90 1766 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyb_4  cm_inst.cc_inst.dlyb_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 28896 0 -1 44352
box -86 -90 2214 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyc_1  cm_inst.cc_inst.dlyc_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 -1 42336
box -86 -90 2326 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyc_2  cm_inst.cc_inst.dlyc_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 18480 0 -1 22176
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyc_4  cm_inst.cc_inst.dlyc_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 41216 0 1 18144
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyd_1  cm_inst.cc_inst.dlyd_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37520 0 -1 12096
box -86 -90 3110 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyd_2  cm_inst.cc_inst.dlyd_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 31136 0 1 14112
box -86 -90 3334 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyd_4  cm_inst.cc_inst.dlyd_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 16128
box -86 -90 3782 1098
use gf180mcu_fd_sc_mcu9t5v0__hold  cm_inst.cc_inst.hold_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 35616 0 1 48384
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtn_1  cm_inst.cc_inst.icgtn_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21392 0 1 20160
box -86 -90 3446 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtn_2  cm_inst.cc_inst.icgtn_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtn_4  cm_inst.cc_inst.icgtn_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 23744 0 1 36288
box -86 -90 4118 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtp_2  cm_inst.cc_inst.icgtp_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 25648 0 1 22176
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtp_4  cm_inst.cc_inst.icgtp_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 28896 0 -1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  cm_inst.cc_inst.inv_1_inst
timestamp 1698431365
transform 1 0 33376 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_2  cm_inst.cc_inst.inv_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 55776 0 1 38304
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_3  cm_inst.cc_inst.inv_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 33712 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_4  cm_inst.cc_inst.inv_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 55328 0 1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_8  cm_inst.cc_inst.inv_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 38304
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_12  cm_inst.cc_inst.inv_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 46592 0 1 26208
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_16  cm_inst.cc_inst.inv_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 46592 0 1 12096
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_20  cm_inst.cc_inst.inv_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 50624 0 1 44352
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_1  cm_inst.cc_inst.invz_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 36288 0 1 44352
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_2  cm_inst.cc_inst.invz_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 26992 0 -1 42336
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_3  cm_inst.cc_inst.invz_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21504 0 -1 40320
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_4  cm_inst.cc_inst.invz_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 -1 42336
box -86 -90 2774 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_8  cm_inst.cc_inst.invz_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 25312 0 1 18144
box -86 -90 4230 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_12  cm_inst.cc_inst.invz_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 -1 18144
box -86 -90 5910 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_1  cm_inst.cc_inst.latq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 45584 0 -1 40320
box -86 -90 2326 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_2  cm_inst.cc_inst.latq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38080 0 -1 38304
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_4  cm_inst.cc_inst.latq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 48944 0 -1 38304
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__latrnq_1  cm_inst.cc_inst.latrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37296 0 -1 36288
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__latrnq_2  cm_inst.cc_inst.latrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 50400 0 -1 22176
box -86 -90 2886 1098
use gf180mcu_fd_sc_mcu9t5v0__latrnq_4  cm_inst.cc_inst.latrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__latrsnq_1  cm_inst.cc_inst.latrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 39536 0 1 10080
box -86 -90 2774 1098
use gf180mcu_fd_sc_mcu9t5v0__latrsnq_2  cm_inst.cc_inst.latrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29792 0 -1 8064
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__latrsnq_4  cm_inst.cc_inst.latrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 23184 0 1 8064
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__latsnq_1  cm_inst.cc_inst.latsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 46368
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__latsnq_2  cm_inst.cc_inst.latsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 33488 0 1 46368
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__latsnq_4  cm_inst.cc_inst.latsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 44352
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  cm_inst.cc_inst.mux2_1_inst
timestamp 1698431365
transform -1 0 52304 0 1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_2  cm_inst.cc_inst.mux2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 38976 0 1 36288
box -86 -90 1766 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_4  cm_inst.cc_inst.mux2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 1 20160
box -86 -90 2214 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  cm_inst.cc_inst.mux4_1_inst
timestamp 1698431365
transform 1 0 52528 0 -1 20160
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_2  cm_inst.cc_inst.mux4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38528 0 1 42336
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_4  cm_inst.cc_inst.mux4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 38976 0 -1 40320
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  cm_inst.cc_inst.nand2_1_inst
timestamp 1698431365
transform -1 0 53984 0 1 38304
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_2  cm_inst.cc_inst.nand2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 36512 0 1 26208
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_4  cm_inst.cc_inst.nand2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 55328 0 1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__nand3_1  cm_inst.cc_inst.nand3_1_inst
timestamp 1698431365
transform 1 0 33600 0 -1 24192
box -86 -90 870 1098
use gf180mcu_fd_sc_mcu9t5v0__nand3_2  cm_inst.cc_inst.nand3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 46256 0 -1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nand3_4  cm_inst.cc_inst.nand3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 48160 0 1 20160
box -86 -90 2886 1098
use gf180mcu_fd_sc_mcu9t5v0__nand4_1  cm_inst.cc_inst.nand4_1_inst
timestamp 1698431365
transform 1 0 40992 0 -1 46368
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__nand4_2  cm_inst.cc_inst.nand4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 46928 0 1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__nand4_4  cm_inst.cc_inst.nand4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 52752 0 -1 44352
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  cm_inst.cc_inst.nor2_1_inst
timestamp 1698431365
transform -1 0 49280 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_2  cm_inst.cc_inst.nor2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 57568 0 -1 36288
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_4  cm_inst.cc_inst.nor2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 41440 0 -1 34272
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__nor3_1  cm_inst.cc_inst.nor3_1_inst
timestamp 1698431365
transform -1 0 58240 0 1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__nor3_2  cm_inst.cc_inst.nor3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 48608 0 -1 18144
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__nor3_4  cm_inst.cc_inst.nor3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 39424 0 1 48384
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__nor4_1  cm_inst.cc_inst.nor4_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 47488 0 1 32256
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__nor4_2  cm_inst.cc_inst.nor4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 52640 0 -1 46368
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__nor4_4  cm_inst.cc_inst.nor4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 49952 0 1 30240
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  cm_inst.cc_inst.oai21_1_inst
timestamp 1698431365
transform 1 0 44688 0 1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_2  cm_inst.cc_inst.oai21_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 35056 0 1 24192
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_4  cm_inst.cc_inst.oai21_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 51520 0 -1 42336
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__oai22_1  cm_inst.cc_inst.oai22_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 37408 0 -1 26208
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__oai22_2  cm_inst.cc_inst.oai22_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 54544 0 1 32256
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__oai22_4  cm_inst.cc_inst.oai22_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 33824 0 -1 22176
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__oai31_1  cm_inst.cc_inst.oai31_1_inst
timestamp 1698431365
transform 1 0 51520 0 -1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__oai31_2  cm_inst.cc_inst.oai31_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 54768 0 1 16128
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__oai31_4  cm_inst.cc_inst.oai31_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 45920 0 -1 46368
box -86 -90 4006 1098
use gf180mcu_fd_sc_mcu9t5v0__oai32_1  cm_inst.cc_inst.oai32_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 35280 0 1 22176
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__oai32_2  cm_inst.cc_inst.oai32_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 54992 0 1 42336
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__oai32_4  cm_inst.cc_inst.oai32_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 34720 0 -1 20160
box -86 -90 4902 1098
use gf180mcu_fd_sc_mcu9t5v0__oai33_1  cm_inst.cc_inst.oai33_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 51184 0 -1 32256
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__oai33_2  cm_inst.cc_inst.oai33_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 39760 0 1 20160
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__oai33_4  cm_inst.cc_inst.oai33_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 48944 0 -1 26208
box -86 -90 5798 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  cm_inst.cc_inst.oai211_1_inst
timestamp 1698431365
transform 1 0 54768 0 1 16128
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_2  cm_inst.cc_inst.oai211_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 42336 0 1 42336
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_4  cm_inst.cc_inst.oai211_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 40432 0 1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__oai221_1  cm_inst.cc_inst.oai221_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 50064 0 -1 40320
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__oai221_2  cm_inst.cc_inst.oai221_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 44688 0 -1 36288
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__oai221_4  cm_inst.cc_inst.oai221_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 58352 0 1 36288
box -86 -90 4902 1098
use gf180mcu_fd_sc_mcu9t5v0__oai222_1  cm_inst.cc_inst.oai222_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 42784 0 -1 38304
box -86 -90 1766 1098
use gf180mcu_fd_sc_mcu9t5v0__oai222_2  cm_inst.cc_inst.oai222_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 53200 0 -1 22176
box -86 -90 3110 1098
use gf180mcu_fd_sc_mcu9t5v0__oai222_4  cm_inst.cc_inst.oai222_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 1 18144
box -86 -90 5798 1098
use gf180mcu_fd_sc_mcu9t5v0__or2_1  cm_inst.cc_inst.or2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 54544 0 1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__or2_2  cm_inst.cc_inst.or2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40992 0 -1 32256
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__or2_4  cm_inst.cc_inst.or2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 58016 0 1 22176
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__or3_1  cm_inst.cc_inst.or3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 46144 0 1 20160
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__or3_2  cm_inst.cc_inst.or3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37744 0 1 44352
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__or3_4  cm_inst.cc_inst.or3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 42448 0 -1 32256
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__or4_1  cm_inst.cc_inst.or4_1_inst
timestamp 1698431365
transform 1 0 50624 0 1 44352
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__or4_2  cm_inst.cc_inst.or4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 46256 0 1 32256
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__or4_4  cm_inst.cc_inst.or4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 49840 0 -1 36288
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffq_1  cm_inst.cc_inst.sdffq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 -1 24192
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffq_2  cm_inst.cc_inst.sdffq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 41888 0 -1 18144
box -86 -90 4566 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffq_4  cm_inst.cc_inst.sdffq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38416 0 1 12096
box -86 -90 5014 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1  cm_inst.cc_inst.sdffrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 16128
box -86 -90 4678 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2  cm_inst.cc_inst.sdffrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 24080 0 1 16128
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4  cm_inst.cc_inst.sdffrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 19600 0 -1 14112
box -86 -90 5350 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1  cm_inst.cc_inst.sdffrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -90 5238 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2  cm_inst.cc_inst.sdffrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21504 0 1 40320
box -86 -90 5462 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4  cm_inst.cc_inst.sdffrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 18928 0 -1 20160
box -86 -90 5910 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1  cm_inst.cc_inst.sdffsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 20160
box -86 -90 5014 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2  cm_inst.cc_inst.sdffsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37520 0 1 14112
box -86 -90 5126 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4  cm_inst.cc_inst.sdffsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 30800 0 1 16128
box -86 -90 5574 1098
use gf180mcu_fd_sc_mcu9t5v0__tieh  cm_inst.cc_inst.tieh_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 52080 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  cm_inst.cc_inst.tiel_inst
timestamp 1698431365
transform 1 0 50400 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_1  cm_inst.cc_inst.xnor2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37968 0 1 32256
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_2  cm_inst.cc_inst.xnor2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 50400 0 1 24192
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_4  cm_inst.cc_inst.xnor2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 46032 0 -1 20160
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor3_1  cm_inst.cc_inst.xnor3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37184 0 -1 46368
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor3_2  cm_inst.cc_inst.xnor3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 41328 0 1 30240
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor3_4  cm_inst.cc_inst.xnor3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 48832 0 -1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_1  cm_inst.cc_inst.xor2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 46480 0 -1 34272
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_2  cm_inst.cc_inst.xor2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 1 34272
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_4  cm_inst.cc_inst.xor2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38192 0 -1 32256
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__xor3_1  cm_inst.cc_inst.xor3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 50176 0 -1 24192
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__xor3_2  cm_inst.cc_inst.xor3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 53312 0 1 12096
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__xor3_4  cm_inst.cc_inst.xor3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 43120 0 -1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_0_478 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 54880 0 1 4032
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_0_494 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 56672 0 1 4032
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_0_502 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 57568 0 1 4032
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_506 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 58016 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_0_508 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 58240 0 1 4032
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 6048
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 6048
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 6048
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 6048
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698431365
transform 1 0 51856 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 6048
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 6048
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_18
timestamp 1698431365
transform 1 0 3360 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_3_20
timestamp 1698431365
transform 1 0 3584 0 -1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_3_29
timestamp 1698431365
transform 1 0 4592 0 -1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_3_61
timestamp 1698431365
transform 1 0 8176 0 -1 8064
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_3_69
timestamp 1698431365
transform 1 0 9072 0 -1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_3_174
timestamp 1698431365
transform 1 0 20832 0 -1 8064
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_182
timestamp 1698431365
transform 1 0 21728 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_3_186
timestamp 1698431365
transform 1 0 22176 0 -1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_189
timestamp 1698431365
transform 1 0 22512 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_3_193
timestamp 1698431365
transform 1 0 22960 0 -1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_3_228
timestamp 1698431365
transform 1 0 26880 0 -1 8064
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_236
timestamp 1698431365
transform 1 0 27776 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_242
timestamp 1698431365
transform 1 0 28448 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_246
timestamp 1698431365
transform 1 0 28896 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_250
timestamp 1698431365
transform 1 0 29344 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_183
timestamp 1698431365
transform 1 0 21840 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_187
timestamp 1698431365
transform 1 0 22288 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_191
timestamp 1698431365
transform 1 0 22736 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_4_226
timestamp 1698431365
transform 1 0 26656 0 1 8064
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_4_234
timestamp 1698431365
transform 1 0 27552 0 1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_237
timestamp 1698431365
transform 1 0 27888 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_4_279
timestamp 1698431365
transform 1 0 32592 0 1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_4_321
timestamp 1698431365
transform 1 0 37296 0 1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_195
timestamp 1698431365
transform 1 0 23184 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_201
timestamp 1698431365
transform 1 0 23856 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_203
timestamp 1698431365
transform 1 0 24080 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_5_261
timestamp 1698431365
transform 1 0 30576 0 -1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_277
timestamp 1698431365
transform 1 0 32368 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_286
timestamp 1698431365
transform 1 0 33376 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_289
timestamp 1698431365
transform 1 0 33712 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_293
timestamp 1698431365
transform 1 0 34160 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_5_330
timestamp 1698431365
transform 1 0 38304 0 -1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_384
timestamp 1698431365
transform 1 0 44352 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_5_387
timestamp 1698431365
transform 1 0 44688 0 -1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_419
timestamp 1698431365
transform 1 0 48272 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_6_155
timestamp 1698431365
transform 1 0 18704 0 1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_163
timestamp 1698431365
transform 1 0 19600 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_167
timestamp 1698431365
transform 1 0 20048 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_216
timestamp 1698431365
transform 1 0 25536 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_6_220
timestamp 1698431365
transform 1 0 25984 0 1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_6_236
timestamp 1698431365
transform 1 0 27776 0 1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_261
timestamp 1698431365
transform 1 0 30576 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_265
timestamp 1698431365
transform 1 0 31024 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_307
timestamp 1698431365
transform 1 0 35728 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_6_341
timestamp 1698431365
transform 1 0 39536 0 1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_349
timestamp 1698431365
transform 1 0 40432 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_353
timestamp 1698431365
transform 1 0 40880 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_357
timestamp 1698431365
transform 1 0 41328 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_361
timestamp 1698431365
transform 1 0 41776 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_6_365
timestamp 1698431365
transform 1 0 42224 0 1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_373
timestamp 1698431365
transform 1 0 43120 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_379
timestamp 1698431365
transform 1 0 43792 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_383
timestamp 1698431365
transform 1 0 44240 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_6_419
timestamp 1698431365
transform 1 0 48272 0 1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_461
timestamp 1698431365
transform 1 0 52976 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_6_464
timestamp 1698431365
transform 1 0 53312 0 1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_6_496
timestamp 1698431365
transform 1 0 56896 0 1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_504
timestamp 1698431365
transform 1 0 57792 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_508
timestamp 1698431365
transform 1 0 58240 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_158
timestamp 1698431365
transform 1 0 19040 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_160
timestamp 1698431365
transform 1 0 19264 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_191
timestamp 1698431365
transform 1 0 22736 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_195
timestamp 1698431365
transform 1 0 23184 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_7_199
timestamp 1698431365
transform 1 0 23632 0 -1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_207
timestamp 1698431365
transform 1 0 24528 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_214
timestamp 1698431365
transform 1 0 25312 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_217
timestamp 1698431365
transform 1 0 25648 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_221
timestamp 1698431365
transform 1 0 26096 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_264
timestamp 1698431365
transform 1 0 30912 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_268
timestamp 1698431365
transform 1 0 31360 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_272
timestamp 1698431365
transform 1 0 31808 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_319
timestamp 1698431365
transform 1 0 37072 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_356
timestamp 1698431365
transform 1 0 41216 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_360
timestamp 1698431365
transform 1 0 41664 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_7_399
timestamp 1698431365
transform 1 0 46032 0 -1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_415
timestamp 1698431365
transform 1 0 47824 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_419
timestamp 1698431365
transform 1 0 48272 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_7_426
timestamp 1698431365
transform 1 0 49056 0 -1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_7_442
timestamp 1698431365
transform 1 0 50848 0 -1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_450
timestamp 1698431365
transform 1 0 51744 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_454
timestamp 1698431365
transform 1 0 52192 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_457
timestamp 1698431365
transform 1 0 52528 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_461
timestamp 1698431365
transform 1 0 52976 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_463
timestamp 1698431365
transform 1 0 53200 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_466
timestamp 1698431365
transform 1 0 53536 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_7_470
timestamp 1698431365
transform 1 0 53984 0 -1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 12096
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 12096
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_139
timestamp 1698431365
transform 1 0 16912 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_141
timestamp 1698431365
transform 1 0 17136 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_192
timestamp 1698431365
transform 1 0 22848 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_194
timestamp 1698431365
transform 1 0 23072 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_226
timestamp 1698431365
transform 1 0 26656 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_8_230
timestamp 1698431365
transform 1 0 27104 0 1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_238
timestamp 1698431365
transform 1 0 28000 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_242
timestamp 1698431365
transform 1 0 28448 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_286
timestamp 1698431365
transform 1 0 33376 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_8_290
timestamp 1698431365
transform 1 0 33824 0 1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_298
timestamp 1698431365
transform 1 0 34720 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_302
timestamp 1698431365
transform 1 0 35168 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_304
timestamp 1698431365
transform 1 0 35392 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_307
timestamp 1698431365
transform 1 0 35728 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_323
timestamp 1698431365
transform 1 0 37520 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_327
timestamp 1698431365
transform 1 0 37968 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_8_375
timestamp 1698431365
transform 1 0 43344 0 1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_383
timestamp 1698431365
transform 1 0 44240 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_395
timestamp 1698431365
transform 1 0 45584 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_399
timestamp 1698431365
transform 1 0 46032 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_401
timestamp 1698431365
transform 1 0 46256 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_438
timestamp 1698431365
transform 1 0 50400 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_442
timestamp 1698431365
transform 1 0 50848 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_445
timestamp 1698431365
transform 1 0 51184 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_449
timestamp 1698431365
transform 1 0 51632 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_453
timestamp 1698431365
transform 1 0 52080 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_461
timestamp 1698431365
transform 1 0 52976 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_463
timestamp 1698431365
transform 1 0 53200 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_8_492
timestamp 1698431365
transform 1 0 56448 0 1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_508
timestamp 1698431365
transform 1 0 58240 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_224
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_9_228
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_236
timestamp 1698431365
transform 1 0 27776 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_240
timestamp 1698431365
transform 1 0 28224 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_242
timestamp 1698431365
transform 1 0 28448 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_245
timestamp 1698431365
transform 1 0 28784 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_9_249
timestamp 1698431365
transform 1 0 29232 0 -1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_257
timestamp 1698431365
transform 1 0 30128 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_261
timestamp 1698431365
transform 1 0 30576 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_263
timestamp 1698431365
transform 1 0 30800 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_9_266
timestamp 1698431365
transform 1 0 31136 0 -1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_9_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_298
timestamp 1698431365
transform 1 0 34720 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_333
timestamp 1698431365
transform 1 0 38640 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_482
timestamp 1698431365
transform 1 0 55328 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_10_139
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_155
timestamp 1698431365
transform 1 0 18704 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_161
timestamp 1698431365
transform 1 0 19376 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_165
timestamp 1698431365
transform 1 0 19824 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_169
timestamp 1698431365
transform 1 0 20272 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_173
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_181
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_222
timestamp 1698431365
transform 1 0 26208 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_228
timestamp 1698431365
transform 1 0 26880 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_259
timestamp 1698431365
transform 1 0 30352 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_263
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_295
timestamp 1698431365
transform 1 0 34384 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_299
timestamp 1698431365
transform 1 0 34832 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_303
timestamp 1698431365
transform 1 0 35280 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_307
timestamp 1698431365
transform 1 0 35728 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_10_368
timestamp 1698431365
transform 1 0 42560 0 1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_376
timestamp 1698431365
transform 1 0 43456 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_378
timestamp 1698431365
transform 1 0 43680 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_453
timestamp 1698431365
transform 1 0 52080 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_504
timestamp 1698431365
transform 1 0 57792 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_508
timestamp 1698431365
transform 1 0 58240 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_144
timestamp 1698431365
transform 1 0 17472 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_190
timestamp 1698431365
transform 1 0 22624 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_194
timestamp 1698431365
transform 1 0 23072 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_197
timestamp 1698431365
transform 1 0 23408 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_201
timestamp 1698431365
transform 1 0 23856 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_205
timestamp 1698431365
transform 1 0 24304 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_207
timestamp 1698431365
transform 1 0 24528 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_264
timestamp 1698431365
transform 1 0 30912 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_266
timestamp 1698431365
transform 1 0 31136 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_336
timestamp 1698431365
transform 1 0 38976 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_340
timestamp 1698431365
transform 1 0 39424 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_344
timestamp 1698431365
transform 1 0 39872 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_346
timestamp 1698431365
transform 1 0 40096 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_358
timestamp 1698431365
transform 1 0 41440 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_362
timestamp 1698431365
transform 1 0 41888 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_11_366
timestamp 1698431365
transform 1 0 42336 0 -1 16128
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_11_398
timestamp 1698431365
transform 1 0 45920 0 -1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_406
timestamp 1698431365
transform 1 0 46816 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_412
timestamp 1698431365
transform 1 0 47488 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_433
timestamp 1698431365
transform 1 0 49840 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_437
timestamp 1698431365
transform 1 0 50288 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_441
timestamp 1698431365
transform 1 0 50736 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_445
timestamp 1698431365
transform 1 0 51184 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_449
timestamp 1698431365
transform 1 0 51632 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_453
timestamp 1698431365
transform 1 0 52080 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_488
timestamp 1698431365
transform 1 0 56000 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 16128
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 16128
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 16128
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 16128
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_12_155
timestamp 1698431365
transform 1 0 18704 0 1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_163
timestamp 1698431365
transform 1 0 19600 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_167
timestamp 1698431365
transform 1 0 20048 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_191
timestamp 1698431365
transform 1 0 22736 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_195
timestamp 1698431365
transform 1 0 23184 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_199
timestamp 1698431365
transform 1 0 23632 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_262
timestamp 1698431365
transform 1 0 30688 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_312
timestamp 1698431365
transform 1 0 36288 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 16128
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_12_333
timestamp 1698431365
transform 1 0 38640 0 1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_12_372
timestamp 1698431365
transform 1 0 43008 0 1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_380
timestamp 1698431365
transform 1 0 43904 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_384
timestamp 1698431365
transform 1 0 44352 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_389
timestamp 1698431365
transform 1 0 44912 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_12_398
timestamp 1698431365
transform 1 0 45920 0 1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_12_412
timestamp 1698431365
transform 1 0 47488 0 1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_422
timestamp 1698431365
transform 1 0 48608 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_426
timestamp 1698431365
transform 1 0 49056 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_430
timestamp 1698431365
transform 1 0 49504 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_433
timestamp 1698431365
transform 1 0 49840 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_437
timestamp 1698431365
transform 1 0 50288 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_441
timestamp 1698431365
transform 1 0 50736 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_445
timestamp 1698431365
transform 1 0 51184 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_449
timestamp 1698431365
transform 1 0 51632 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_487
timestamp 1698431365
transform 1 0 55888 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_491
timestamp 1698431365
transform 1 0 56336 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_495
timestamp 1698431365
transform 1 0 56784 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_499
timestamp 1698431365
transform 1 0 57232 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_503
timestamp 1698431365
transform 1 0 57680 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_507
timestamp 1698431365
transform 1 0 58128 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 18144
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 18144
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_144
timestamp 1698431365
transform 1 0 17472 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_197
timestamp 1698431365
transform 1 0 23408 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_201
timestamp 1698431365
transform 1 0 23856 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_203
timestamp 1698431365
transform 1 0 24080 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_257
timestamp 1698431365
transform 1 0 30128 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_263
timestamp 1698431365
transform 1 0 30800 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_267
timestamp 1698431365
transform 1 0 31248 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_271
timestamp 1698431365
transform 1 0 31696 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_275
timestamp 1698431365
transform 1 0 32144 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_13_318
timestamp 1698431365
transform 1 0 36960 0 -1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_334
timestamp 1698431365
transform 1 0 38752 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_338
timestamp 1698431365
transform 1 0 39200 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_342
timestamp 1698431365
transform 1 0 39648 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_346
timestamp 1698431365
transform 1 0 40096 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_356
timestamp 1698431365
transform 1 0 41216 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_360
timestamp 1698431365
transform 1 0 41664 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_13_402
timestamp 1698431365
transform 1 0 46368 0 -1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_412
timestamp 1698431365
transform 1 0 47488 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_436
timestamp 1698431365
transform 1 0 50176 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_440
timestamp 1698431365
transform 1 0 50624 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_443
timestamp 1698431365
transform 1 0 50960 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_447
timestamp 1698431365
transform 1 0 51408 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_451
timestamp 1698431365
transform 1 0 51856 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_488
timestamp 1698431365
transform 1 0 56000 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 18144
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 18144
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_169
timestamp 1698431365
transform 1 0 20272 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_214
timestamp 1698431365
transform 1 0 25312 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_218
timestamp 1698431365
transform 1 0 25760 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_222
timestamp 1698431365
transform 1 0 26208 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_226
timestamp 1698431365
transform 1 0 26656 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_230
timestamp 1698431365
transform 1 0 27104 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_262
timestamp 1698431365
transform 1 0 30688 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_266
timestamp 1698431365
transform 1 0 31136 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_270
timestamp 1698431365
transform 1 0 31584 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_290
timestamp 1698431365
transform 1 0 33824 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_294
timestamp 1698431365
transform 1 0 34272 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_298
timestamp 1698431365
transform 1 0 34720 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_302
timestamp 1698431365
transform 1 0 35168 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_306
timestamp 1698431365
transform 1 0 35616 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_310
timestamp 1698431365
transform 1 0 36064 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_14_321
timestamp 1698431365
transform 1 0 37296 0 1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_329
timestamp 1698431365
transform 1 0 38192 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_335
timestamp 1698431365
transform 1 0 38864 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_382
timestamp 1698431365
transform 1 0 44128 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_397
timestamp 1698431365
transform 1 0 45808 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_401
timestamp 1698431365
transform 1 0 46256 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_405
timestamp 1698431365
transform 1 0 46704 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_437
timestamp 1698431365
transform 1 0 50288 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_441
timestamp 1698431365
transform 1 0 50736 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_445
timestamp 1698431365
transform 1 0 51184 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_449
timestamp 1698431365
transform 1 0 51632 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_453
timestamp 1698431365
transform 1 0 52080 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_508
timestamp 1698431365
transform 1 0 58240 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 20160
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_15_88
timestamp 1698431365
transform 1 0 11200 0 -1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_96
timestamp 1698431365
transform 1 0 12096 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_155
timestamp 1698431365
transform 1 0 18704 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_231
timestamp 1698431365
transform 1 0 27216 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_261
timestamp 1698431365
transform 1 0 30576 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_265
timestamp 1698431365
transform 1 0 31024 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_273
timestamp 1698431365
transform 1 0 31920 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_277
timestamp 1698431365
transform 1 0 32368 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_341
timestamp 1698431365
transform 1 0 39536 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_343
timestamp 1698431365
transform 1 0 39760 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_396
timestamp 1698431365
transform 1 0 45696 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_398
timestamp 1698431365
transform 1 0 45920 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_453
timestamp 1698431365
transform 1 0 52080 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_488
timestamp 1698431365
transform 1 0 56000 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_15_496
timestamp 1698431365
transform 1 0 56896 0 -1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_504
timestamp 1698431365
transform 1 0 57792 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_508
timestamp 1698431365
transform 1 0 58240 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 20160
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 20160
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_157
timestamp 1698431365
transform 1 0 18928 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_161
timestamp 1698431365
transform 1 0 19376 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_167
timestamp 1698431365
transform 1 0 20048 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_209
timestamp 1698431365
transform 1 0 24752 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_217
timestamp 1698431365
transform 1 0 25648 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_221
timestamp 1698431365
transform 1 0 26096 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_16_225
timestamp 1698431365
transform 1 0 26544 0 1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_16_265
timestamp 1698431365
transform 1 0 31024 0 1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_281
timestamp 1698431365
transform 1 0 32816 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_288
timestamp 1698431365
transform 1 0 33600 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_292
timestamp 1698431365
transform 1 0 34048 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_295
timestamp 1698431365
transform 1 0 34384 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_299
timestamp 1698431365
transform 1 0 34832 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_303
timestamp 1698431365
transform 1 0 35280 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_307
timestamp 1698431365
transform 1 0 35728 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_343
timestamp 1698431365
transform 1 0 39760 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_353
timestamp 1698431365
transform 1 0 40880 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_357
timestamp 1698431365
transform 1 0 41328 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_16_361
timestamp 1698431365
transform 1 0 41776 0 1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_369
timestamp 1698431365
transform 1 0 42672 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_389
timestamp 1698431365
transform 1 0 44912 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_392
timestamp 1698431365
transform 1 0 45248 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_396
timestamp 1698431365
transform 1 0 45696 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_411
timestamp 1698431365
transform 1 0 47376 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_415
timestamp 1698431365
transform 1 0 47824 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_417
timestamp 1698431365
transform 1 0 48048 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_443
timestamp 1698431365
transform 1 0 50960 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_449
timestamp 1698431365
transform 1 0 51632 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_453
timestamp 1698431365
transform 1 0 52080 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_493
timestamp 1698431365
transform 1 0 56560 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_497
timestamp 1698431365
transform 1 0 57008 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_16_501
timestamp 1698431365
transform 1 0 57456 0 1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_6
timestamp 1698431365
transform 1 0 2016 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_17_10
timestamp 1698431365
transform 1 0 2464 0 -1 22176
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_17_42
timestamp 1698431365
transform 1 0 6048 0 -1 22176
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_17_58
timestamp 1698431365
transform 1 0 7840 0 -1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 22176
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_17_88
timestamp 1698431365
transform 1 0 11200 0 -1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_96
timestamp 1698431365
transform 1 0 12096 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_100
timestamp 1698431365
transform 1 0 12544 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_149
timestamp 1698431365
transform 1 0 18032 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_189
timestamp 1698431365
transform 1 0 22512 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_193
timestamp 1698431365
transform 1 0 22960 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_197
timestamp 1698431365
transform 1 0 23408 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_199
timestamp 1698431365
transform 1 0 23632 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_202
timestamp 1698431365
transform 1 0 23968 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_225
timestamp 1698431365
transform 1 0 26544 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_17_229
timestamp 1698431365
transform 1 0 26992 0 -1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_237
timestamp 1698431365
transform 1 0 27888 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_241
timestamp 1698431365
transform 1 0 28336 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_243
timestamp 1698431365
transform 1 0 28560 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_257
timestamp 1698431365
transform 1 0 30128 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_17_261
timestamp 1698431365
transform 1 0 30576 0 -1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_269
timestamp 1698431365
transform 1 0 31472 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_273
timestamp 1698431365
transform 1 0 31920 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_286
timestamp 1698431365
transform 1 0 33376 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_324
timestamp 1698431365
transform 1 0 37632 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_328
timestamp 1698431365
transform 1 0 38080 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_336
timestamp 1698431365
transform 1 0 38976 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_342
timestamp 1698431365
transform 1 0 39648 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_356
timestamp 1698431365
transform 1 0 41216 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_363
timestamp 1698431365
transform 1 0 42000 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_367
timestamp 1698431365
transform 1 0 42448 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_17_402
timestamp 1698431365
transform 1 0 46368 0 -1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_410
timestamp 1698431365
transform 1 0 47264 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_426
timestamp 1698431365
transform 1 0 49056 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_430
timestamp 1698431365
transform 1 0 49504 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_434
timestamp 1698431365
transform 1 0 49952 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_496
timestamp 1698431365
transform 1 0 56896 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_17_500
timestamp 1698431365
transform 1 0 57344 0 -1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_41
timestamp 1698431365
transform 1 0 5936 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_18_45
timestamp 1698431365
transform 1 0 6384 0 1 22176
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_18_77
timestamp 1698431365
transform 1 0 9968 0 1 22176
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_18_93
timestamp 1698431365
transform 1 0 11760 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 22176
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_123
timestamp 1698431365
transform 1 0 15120 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_137
timestamp 1698431365
transform 1 0 16688 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_18_141
timestamp 1698431365
transform 1 0 17136 0 1 22176
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_18_157
timestamp 1698431365
transform 1 0 18928 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_165
timestamp 1698431365
transform 1 0 19824 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 22176
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_18_263
timestamp 1698431365
transform 1 0 30800 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_271
timestamp 1698431365
transform 1 0 31696 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_275
timestamp 1698431365
transform 1 0 32144 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_277
timestamp 1698431365
transform 1 0 32368 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_280
timestamp 1698431365
transform 1 0 32704 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_290
timestamp 1698431365
transform 1 0 33824 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_294
timestamp 1698431365
transform 1 0 34272 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_298
timestamp 1698431365
transform 1 0 34720 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_300
timestamp 1698431365
transform 1 0 34944 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_333
timestamp 1698431365
transform 1 0 38640 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_339
timestamp 1698431365
transform 1 0 39312 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_343
timestamp 1698431365
transform 1 0 39760 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_346
timestamp 1698431365
transform 1 0 40096 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_350
timestamp 1698431365
transform 1 0 40544 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_354
timestamp 1698431365
transform 1 0 40992 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_366
timestamp 1698431365
transform 1 0 42336 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_370
timestamp 1698431365
transform 1 0 42784 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_374
timestamp 1698431365
transform 1 0 43232 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_378
timestamp 1698431365
transform 1 0 43680 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_382
timestamp 1698431365
transform 1 0 44128 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_18_391
timestamp 1698431365
transform 1 0 45136 0 1 22176
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_423
timestamp 1698431365
transform 1 0 48720 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_427
timestamp 1698431365
transform 1 0 49168 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_429
timestamp 1698431365
transform 1 0 49392 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_432
timestamp 1698431365
transform 1 0 49728 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_436
timestamp 1698431365
transform 1 0 50176 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_440
timestamp 1698431365
transform 1 0 50624 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_444
timestamp 1698431365
transform 1 0 51072 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_447
timestamp 1698431365
transform 1 0 51408 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_506
timestamp 1698431365
transform 1 0 58016 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_508
timestamp 1698431365
transform 1 0 58240 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_19_108
timestamp 1698431365
transform 1 0 13440 0 -1 24192
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_19_124
timestamp 1698431365
transform 1 0 15232 0 -1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_132
timestamp 1698431365
transform 1 0 16128 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_144
timestamp 1698431365
transform 1 0 17472 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_187
timestamp 1698431365
transform 1 0 22288 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_191
timestamp 1698431365
transform 1 0 22736 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_195
timestamp 1698431365
transform 1 0 23184 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_199
timestamp 1698431365
transform 1 0 23632 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_205
timestamp 1698431365
transform 1 0 24304 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_230
timestamp 1698431365
transform 1 0 27104 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_234
timestamp 1698431365
transform 1 0 27552 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_238
timestamp 1698431365
transform 1 0 28000 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_242
timestamp 1698431365
transform 1 0 28448 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_278
timestamp 1698431365
transform 1 0 32480 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_286
timestamp 1698431365
transform 1 0 33376 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_337
timestamp 1698431365
transform 1 0 39088 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_341
timestamp 1698431365
transform 1 0 39536 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_345
timestamp 1698431365
transform 1 0 39984 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_378
timestamp 1698431365
transform 1 0 43680 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_382
timestamp 1698431365
transform 1 0 44128 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_386
timestamp 1698431365
transform 1 0 44576 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_407
timestamp 1698431365
transform 1 0 46928 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_411
timestamp 1698431365
transform 1 0 47376 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_415
timestamp 1698431365
transform 1 0 47824 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_419
timestamp 1698431365
transform 1 0 48272 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_426
timestamp 1698431365
transform 1 0 49056 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_432
timestamp 1698431365
transform 1 0 49728 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_496
timestamp 1698431365
transform 1 0 56896 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_19_500
timestamp 1698431365
transform 1 0 57344 0 -1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_111
timestamp 1698431365
transform 1 0 13776 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_20_115
timestamp 1698431365
transform 1 0 14224 0 1 24192
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_20_207
timestamp 1698431365
transform 1 0 24528 0 1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_227
timestamp 1698431365
transform 1 0 26768 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_237
timestamp 1698431365
transform 1 0 27888 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_20_256
timestamp 1698431365
transform 1 0 30016 0 1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_264
timestamp 1698431365
transform 1 0 30912 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_268
timestamp 1698431365
transform 1 0 31360 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_272
timestamp 1698431365
transform 1 0 31808 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_283
timestamp 1698431365
transform 1 0 33040 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_287
timestamp 1698431365
transform 1 0 33488 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_291
timestamp 1698431365
transform 1 0 33936 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_333
timestamp 1698431365
transform 1 0 38640 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_20_335
timestamp 1698431365
transform 1 0 38864 0 1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_344
timestamp 1698431365
transform 1 0 39872 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_20_384
timestamp 1698431365
transform 1 0 44352 0 1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_20_391
timestamp 1698431365
transform 1 0 45136 0 1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_394
timestamp 1698431365
transform 1 0 45472 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_436
timestamp 1698431365
transform 1 0 50176 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_461
timestamp 1698431365
transform 1 0 52976 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_465
timestamp 1698431365
transform 1 0 53424 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_20_508
timestamp 1698431365
transform 1 0 58240 0 1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_6
timestamp 1698431365
transform 1 0 2016 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_10
timestamp 1698431365
transform 1 0 2464 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_26
timestamp 1698431365
transform 1 0 4256 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_63
timestamp 1698431365
transform 1 0 8400 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_21_124
timestamp 1698431365
transform 1 0 15232 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_132
timestamp 1698431365
transform 1 0 16128 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_207
timestamp 1698431365
transform 1 0 24528 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_236
timestamp 1698431365
transform 1 0 27776 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_256
timestamp 1698431365
transform 1 0 30016 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_260
timestamp 1698431365
transform 1 0 30464 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_272
timestamp 1698431365
transform 1 0 31808 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_274
timestamp 1698431365
transform 1 0 32032 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_290
timestamp 1698431365
transform 1 0 33824 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_328
timestamp 1698431365
transform 1 0 38080 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_373
timestamp 1698431365
transform 1 0 43120 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_375
timestamp 1698431365
transform 1 0 43344 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_424
timestamp 1698431365
transform 1 0 48832 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_476
timestamp 1698431365
transform 1 0 54656 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_480
timestamp 1698431365
transform 1 0 55104 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_484
timestamp 1698431365
transform 1 0 55552 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_488
timestamp 1698431365
transform 1 0 56000 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_496
timestamp 1698431365
transform 1 0 56896 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_21_500
timestamp 1698431365
transform 1 0 57344 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 26208
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_69
timestamp 1698431365
transform 1 0 9072 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_22_139
timestamp 1698431365
transform 1 0 16912 0 1 26208
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_181
timestamp 1698431365
transform 1 0 21616 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_22_185
timestamp 1698431365
transform 1 0 22064 0 1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_193
timestamp 1698431365
transform 1 0 22960 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_208
timestamp 1698431365
transform 1 0 24640 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_22_212
timestamp 1698431365
transform 1 0 25088 0 1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_251
timestamp 1698431365
transform 1 0 29456 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_254
timestamp 1698431365
transform 1 0 29792 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_258
timestamp 1698431365
transform 1 0 30240 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_294
timestamp 1698431365
transform 1 0 34272 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_296
timestamp 1698431365
transform 1 0 34496 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_328
timestamp 1698431365
transform 1 0 38080 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_332
timestamp 1698431365
transform 1 0 38528 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_341
timestamp 1698431365
transform 1 0 39536 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_369
timestamp 1698431365
transform 1 0 42672 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_373
timestamp 1698431365
transform 1 0 43120 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_377
timestamp 1698431365
transform 1 0 43568 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_381
timestamp 1698431365
transform 1 0 44016 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_400
timestamp 1698431365
transform 1 0 46144 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_430
timestamp 1698431365
transform 1 0 49504 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_434
timestamp 1698431365
transform 1 0 49952 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_438
timestamp 1698431365
transform 1 0 50400 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_22_488
timestamp 1698431365
transform 1 0 56000 0 1 26208
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_504
timestamp 1698431365
transform 1 0 57792 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_508
timestamp 1698431365
transform 1 0 58240 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_6
timestamp 1698431365
transform 1 0 2016 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_23_46
timestamp 1698431365
transform 1 0 6496 0 -1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_23_62
timestamp 1698431365
transform 1 0 8288 0 -1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_135
timestamp 1698431365
transform 1 0 16464 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_152
timestamp 1698431365
transform 1 0 18368 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_23_166
timestamp 1698431365
transform 1 0 19936 0 -1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_23_198
timestamp 1698431365
transform 1 0 23520 0 -1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_247
timestamp 1698431365
transform 1 0 29008 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_251
timestamp 1698431365
transform 1 0 29456 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_264
timestamp 1698431365
transform 1 0 30912 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_329
timestamp 1698431365
transform 1 0 38192 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_333
timestamp 1698431365
transform 1 0 38640 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_335
timestamp 1698431365
transform 1 0 38864 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_368
timestamp 1698431365
transform 1 0 42560 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_372
timestamp 1698431365
transform 1 0 43008 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_376
timestamp 1698431365
transform 1 0 43456 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_380
timestamp 1698431365
transform 1 0 43904 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_384
timestamp 1698431365
transform 1 0 44352 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_386
timestamp 1698431365
transform 1 0 44576 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_389
timestamp 1698431365
transform 1 0 44912 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_393
timestamp 1698431365
transform 1 0 45360 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_397
timestamp 1698431365
transform 1 0 45808 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_426
timestamp 1698431365
transform 1 0 49056 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_430
timestamp 1698431365
transform 1 0 49504 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_434
timestamp 1698431365
transform 1 0 49952 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_438
timestamp 1698431365
transform 1 0 50400 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_442
timestamp 1698431365
transform 1 0 50848 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_446
timestamp 1698431365
transform 1 0 51296 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_458
timestamp 1698431365
transform 1 0 52640 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_489
timestamp 1698431365
transform 1 0 56112 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_23_496
timestamp 1698431365
transform 1 0 56896 0 -1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_504
timestamp 1698431365
transform 1 0 57792 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_508
timestamp 1698431365
transform 1 0 58240 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_24_45
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_24_77
timestamp 1698431365
transform 1 0 9968 0 1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_93
timestamp 1698431365
transform 1 0 11760 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_95
timestamp 1698431365
transform 1 0 11984 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_100
timestamp 1698431365
transform 1 0 12544 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_111
timestamp 1698431365
transform 1 0 13776 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_152
timestamp 1698431365
transform 1 0 18368 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_154
timestamp 1698431365
transform 1 0 18592 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_24_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_201
timestamp 1698431365
transform 1 0 23856 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_203
timestamp 1698431365
transform 1 0 24080 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_242
timestamp 1698431365
transform 1 0 28448 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_253
timestamp 1698431365
transform 1 0 29680 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_257
timestamp 1698431365
transform 1 0 30128 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_264
timestamp 1698431365
transform 1 0 30912 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_268
timestamp 1698431365
transform 1 0 31360 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_272
timestamp 1698431365
transform 1 0 31808 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_290
timestamp 1698431365
transform 1 0 33824 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_292
timestamp 1698431365
transform 1 0 34048 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_333
timestamp 1698431365
transform 1 0 38640 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_337
timestamp 1698431365
transform 1 0 39088 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_341
timestamp 1698431365
transform 1 0 39536 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_349
timestamp 1698431365
transform 1 0 40432 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_351
timestamp 1698431365
transform 1 0 40656 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_358
timestamp 1698431365
transform 1 0 41440 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_362
timestamp 1698431365
transform 1 0 41888 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_366
timestamp 1698431365
transform 1 0 42336 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_370
timestamp 1698431365
transform 1 0 42784 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_24_374
timestamp 1698431365
transform 1 0 43232 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_382
timestamp 1698431365
transform 1 0 44128 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_389
timestamp 1698431365
transform 1 0 44912 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_392
timestamp 1698431365
transform 1 0 45248 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_396
timestamp 1698431365
transform 1 0 45696 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_400
timestamp 1698431365
transform 1 0 46144 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_404
timestamp 1698431365
transform 1 0 46592 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_406
timestamp 1698431365
transform 1 0 46816 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_423
timestamp 1698431365
transform 1 0 48720 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_24_427
timestamp 1698431365
transform 1 0 49168 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_437
timestamp 1698431365
transform 1 0 50288 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_441
timestamp 1698431365
transform 1 0 50736 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_445
timestamp 1698431365
transform 1 0 51184 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_451
timestamp 1698431365
transform 1 0 51856 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_461
timestamp 1698431365
transform 1 0 52976 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_465
timestamp 1698431365
transform 1 0 53424 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_492
timestamp 1698431365
transform 1 0 56448 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_24_496
timestamp 1698431365
transform 1 0 56896 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_504
timestamp 1698431365
transform 1 0 57792 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_508
timestamp 1698431365
transform 1 0 58240 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_6
timestamp 1698431365
transform 1 0 2016 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_10
timestamp 1698431365
transform 1 0 2464 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_12
timestamp 1698431365
transform 1 0 2688 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_51
timestamp 1698431365
transform 1 0 7056 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_25_55
timestamp 1698431365
transform 1 0 7504 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_63
timestamp 1698431365
transform 1 0 8400 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_67
timestamp 1698431365
transform 1 0 8848 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_76
timestamp 1698431365
transform 1 0 9856 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_78
timestamp 1698431365
transform 1 0 10080 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_95
timestamp 1698431365
transform 1 0 11984 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_109
timestamp 1698431365
transform 1 0 13552 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_111
timestamp 1698431365
transform 1 0 13776 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_125
timestamp 1698431365
transform 1 0 15344 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_127
timestamp 1698431365
transform 1 0 15568 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_146
timestamp 1698431365
transform 1 0 17696 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_148
timestamp 1698431365
transform 1 0 17920 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_196
timestamp 1698431365
transform 1 0 23296 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_200
timestamp 1698431365
transform 1 0 23744 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_235
timestamp 1698431365
transform 1 0 27664 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_237
timestamp 1698431365
transform 1 0 27888 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_25_250
timestamp 1698431365
transform 1 0 29344 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_258
timestamp 1698431365
transform 1 0 30240 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_25_261
timestamp 1698431365
transform 1 0 30576 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_269
timestamp 1698431365
transform 1 0 31472 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_294
timestamp 1698431365
transform 1 0 34272 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_296
timestamp 1698431365
transform 1 0 34496 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_313
timestamp 1698431365
transform 1 0 36400 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_324
timestamp 1698431365
transform 1 0 37632 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_332
timestamp 1698431365
transform 1 0 38528 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_336
timestamp 1698431365
transform 1 0 38976 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_339
timestamp 1698431365
transform 1 0 39312 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_343
timestamp 1698431365
transform 1 0 39760 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_358
timestamp 1698431365
transform 1 0 41440 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_362
timestamp 1698431365
transform 1 0 41888 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_366
timestamp 1698431365
transform 1 0 42336 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_25_370
timestamp 1698431365
transform 1 0 42784 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_378
timestamp 1698431365
transform 1 0 43680 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_382
timestamp 1698431365
transform 1 0 44128 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_417
timestamp 1698431365
transform 1 0 48048 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_419
timestamp 1698431365
transform 1 0 48272 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_426
timestamp 1698431365
transform 1 0 49056 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_430
timestamp 1698431365
transform 1 0 49504 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_432
timestamp 1698431365
transform 1 0 49728 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_435
timestamp 1698431365
transform 1 0 50064 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_439
timestamp 1698431365
transform 1 0 50512 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_443
timestamp 1698431365
transform 1 0 50960 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_447
timestamp 1698431365
transform 1 0 51408 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_451
timestamp 1698431365
transform 1 0 51856 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_457
timestamp 1698431365
transform 1 0 52528 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 30240
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_69
timestamp 1698431365
transform 1 0 9072 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_73
timestamp 1698431365
transform 1 0 9520 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_111
timestamp 1698431365
transform 1 0 13776 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 30240
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_139
timestamp 1698431365
transform 1 0 16912 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_143
timestamp 1698431365
transform 1 0 17360 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_189
timestamp 1698431365
transform 1 0 22512 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_191
timestamp 1698431365
transform 1 0 22736 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_222
timestamp 1698431365
transform 1 0 26208 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_224
timestamp 1698431365
transform 1 0 26432 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_271
timestamp 1698431365
transform 1 0 31696 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_275
timestamp 1698431365
transform 1 0 32144 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_345
timestamp 1698431365
transform 1 0 39984 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_389
timestamp 1698431365
transform 1 0 44912 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_434
timestamp 1698431365
transform 1 0 49952 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_438
timestamp 1698431365
transform 1 0 50400 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_463
timestamp 1698431365
transform 1 0 53200 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_465
timestamp 1698431365
transform 1 0 53424 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_506
timestamp 1698431365
transform 1 0 58016 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_508
timestamp 1698431365
transform 1 0 58240 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_27_56
timestamp 1698431365
transform 1 0 7616 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_78
timestamp 1698431365
transform 1 0 10080 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_107
timestamp 1698431365
transform 1 0 13328 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_109
timestamp 1698431365
transform 1 0 13552 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_129
timestamp 1698431365
transform 1 0 15792 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_133
timestamp 1698431365
transform 1 0 16240 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_183
timestamp 1698431365
transform 1 0 21840 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_27_187
timestamp 1698431365
transform 1 0 22288 0 -1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_203
timestamp 1698431365
transform 1 0 24080 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_27_240
timestamp 1698431365
transform 1 0 28224 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_248
timestamp 1698431365
transform 1 0 29120 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_286
timestamp 1698431365
transform 1 0 33376 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_296
timestamp 1698431365
transform 1 0 34496 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_27_300
timestamp 1698431365
transform 1 0 34944 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_308
timestamp 1698431365
transform 1 0 35840 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_311
timestamp 1698431365
transform 1 0 36176 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_317
timestamp 1698431365
transform 1 0 36848 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_323
timestamp 1698431365
transform 1 0 37520 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_327
timestamp 1698431365
transform 1 0 37968 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_364
timestamp 1698431365
transform 1 0 42112 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_366
timestamp 1698431365
transform 1 0 42336 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_428
timestamp 1698431365
transform 1 0 49280 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_442
timestamp 1698431365
transform 1 0 50848 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_444
timestamp 1698431365
transform 1 0 51072 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_501
timestamp 1698431365
transform 1 0 57456 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_505
timestamp 1698431365
transform 1 0 57904 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 32256
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_28_61
timestamp 1698431365
transform 1 0 8176 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_69
timestamp 1698431365
transform 1 0 9072 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_73
timestamp 1698431365
transform 1 0 9520 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_28_115
timestamp 1698431365
transform 1 0 14224 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_123
timestamp 1698431365
transform 1 0 15120 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_183
timestamp 1698431365
transform 1 0 21840 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_28_187
timestamp 1698431365
transform 1 0 22288 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_28_221
timestamp 1698431365
transform 1 0 26096 0 1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_237
timestamp 1698431365
transform 1 0 27888 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_303
timestamp 1698431365
transform 1 0 35280 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_28_307
timestamp 1698431365
transform 1 0 35728 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_321
timestamp 1698431365
transform 1 0 37296 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_325
timestamp 1698431365
transform 1 0 37744 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_370
timestamp 1698431365
transform 1 0 42784 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_374
timestamp 1698431365
transform 1 0 43232 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_378
timestamp 1698431365
transform 1 0 43680 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_401
timestamp 1698431365
transform 1 0 46256 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_418
timestamp 1698431365
transform 1 0 48160 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_422
timestamp 1698431365
transform 1 0 48608 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_430
timestamp 1698431365
transform 1 0 49504 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_434
timestamp 1698431365
transform 1 0 49952 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_438
timestamp 1698431365
transform 1 0 50400 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_495
timestamp 1698431365
transform 1 0 56784 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_28_499
timestamp 1698431365
transform 1 0 57232 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_507
timestamp 1698431365
transform 1 0 58128 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_10
timestamp 1698431365
transform 1 0 2464 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_14
timestamp 1698431365
transform 1 0 2912 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_16
timestamp 1698431365
transform 1 0 3136 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_29_51
timestamp 1698431365
transform 1 0 7056 0 -1 34272
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 34272
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_88
timestamp 1698431365
transform 1 0 11200 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_92
timestamp 1698431365
transform 1 0 11648 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_29_98
timestamp 1698431365
transform 1 0 12320 0 -1 34272
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_130
timestamp 1698431365
transform 1 0 15904 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_144
timestamp 1698431365
transform 1 0 17472 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_160
timestamp 1698431365
transform 1 0 19264 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_166
timestamp 1698431365
transform 1 0 19936 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_170
timestamp 1698431365
transform 1 0 20384 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_172
timestamp 1698431365
transform 1 0 20608 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_193
timestamp 1698431365
transform 1 0 22960 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_221
timestamp 1698431365
transform 1 0 26096 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_223
timestamp 1698431365
transform 1 0 26320 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_29_235
timestamp 1698431365
transform 1 0 27664 0 -1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_243
timestamp 1698431365
transform 1 0 28560 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_29_247
timestamp 1698431365
transform 1 0 29008 0 -1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_255
timestamp 1698431365
transform 1 0 29904 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_257
timestamp 1698431365
transform 1 0 30128 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_260
timestamp 1698431365
transform 1 0 30464 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_277
timestamp 1698431365
transform 1 0 32368 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_322
timestamp 1698431365
transform 1 0 37408 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_326
timestamp 1698431365
transform 1 0 37856 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_29_329
timestamp 1698431365
transform 1 0 38192 0 -1 34272
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_345
timestamp 1698431365
transform 1 0 39984 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_347
timestamp 1698431365
transform 1 0 40208 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_356
timestamp 1698431365
transform 1 0 41216 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_376
timestamp 1698431365
transform 1 0 43456 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_378
timestamp 1698431365
transform 1 0 43680 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_381
timestamp 1698431365
transform 1 0 44016 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_385
timestamp 1698431365
transform 1 0 44464 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_389
timestamp 1698431365
transform 1 0 44912 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_403
timestamp 1698431365
transform 1 0 46480 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_407
timestamp 1698431365
transform 1 0 46928 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_411
timestamp 1698431365
transform 1 0 47376 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_415
timestamp 1698431365
transform 1 0 47824 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_417
timestamp 1698431365
transform 1 0 48048 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_430
timestamp 1698431365
transform 1 0 49504 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_434
timestamp 1698431365
transform 1 0 49952 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_438
timestamp 1698431365
transform 1 0 50400 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_442
timestamp 1698431365
transform 1 0 50848 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_446
timestamp 1698431365
transform 1 0 51296 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_450
timestamp 1698431365
transform 1 0 51744 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_467
timestamp 1698431365
transform 1 0 53648 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_471
timestamp 1698431365
transform 1 0 54096 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_475
timestamp 1698431365
transform 1 0 54544 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_481
timestamp 1698431365
transform 1 0 55216 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_485
timestamp 1698431365
transform 1 0 55664 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_488
timestamp 1698431365
transform 1 0 56000 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 34272
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_508
timestamp 1698431365
transform 1 0 58240 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 34272
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_30_41
timestamp 1698431365
transform 1 0 5936 0 1 34272
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_30_111
timestamp 1698431365
transform 1 0 13776 0 1 34272
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_127
timestamp 1698431365
transform 1 0 15568 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_131
timestamp 1698431365
transform 1 0 16016 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_134
timestamp 1698431365
transform 1 0 16352 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_138
timestamp 1698431365
transform 1 0 16800 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_168
timestamp 1698431365
transform 1 0 20160 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_194
timestamp 1698431365
transform 1 0 23072 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_198
timestamp 1698431365
transform 1 0 23520 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_202
timestamp 1698431365
transform 1 0 23968 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_206
timestamp 1698431365
transform 1 0 24416 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_231
timestamp 1698431365
transform 1 0 27216 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_30_253
timestamp 1698431365
transform 1 0 29680 0 1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_30_305
timestamp 1698431365
transform 1 0 35504 0 1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_313
timestamp 1698431365
transform 1 0 36400 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_322
timestamp 1698431365
transform 1 0 37408 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_326
timestamp 1698431365
transform 1 0 37856 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_337
timestamp 1698431365
transform 1 0 39088 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_347
timestamp 1698431365
transform 1 0 40208 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_353
timestamp 1698431365
transform 1 0 40880 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_359
timestamp 1698431365
transform 1 0 41552 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_363
timestamp 1698431365
transform 1 0 42000 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_367
timestamp 1698431365
transform 1 0 42448 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_375
timestamp 1698431365
transform 1 0 43344 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_379
timestamp 1698431365
transform 1 0 43792 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_383
timestamp 1698431365
transform 1 0 44240 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_391
timestamp 1698431365
transform 1 0 45136 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_395
timestamp 1698431365
transform 1 0 45584 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_399
timestamp 1698431365
transform 1 0 46032 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_30_403
timestamp 1698431365
transform 1 0 46480 0 1 34272
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_30_419
timestamp 1698431365
transform 1 0 48272 0 1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_427
timestamp 1698431365
transform 1 0 49168 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_431
timestamp 1698431365
transform 1 0 49616 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_435
timestamp 1698431365
transform 1 0 50064 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_439
timestamp 1698431365
transform 1 0 50512 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_443
timestamp 1698431365
transform 1 0 50960 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_453
timestamp 1698431365
transform 1 0 52080 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_474
timestamp 1698431365
transform 1 0 54432 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_483
timestamp 1698431365
transform 1 0 55440 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_487
timestamp 1698431365
transform 1 0 55888 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_491
timestamp 1698431365
transform 1 0 56336 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_30_495
timestamp 1698431365
transform 1 0 56784 0 1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_503
timestamp 1698431365
transform 1 0 57680 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_507
timestamp 1698431365
transform 1 0 58128 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_6
timestamp 1698431365
transform 1 0 2016 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_14
timestamp 1698431365
transform 1 0 2912 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_31_49
timestamp 1698431365
transform 1 0 6832 0 -1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_65
timestamp 1698431365
transform 1 0 8624 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_80
timestamp 1698431365
transform 1 0 10304 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_84
timestamp 1698431365
transform 1 0 10752 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698431365
transform 1 0 14784 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_128
timestamp 1698431365
transform 1 0 15680 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_132
timestamp 1698431365
transform 1 0 16128 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_178
timestamp 1698431365
transform 1 0 21280 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_214
timestamp 1698431365
transform 1 0 25312 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_256
timestamp 1698431365
transform 1 0 30016 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_264
timestamp 1698431365
transform 1 0 30912 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_274
timestamp 1698431365
transform 1 0 32032 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_278
timestamp 1698431365
transform 1 0 32480 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_290
timestamp 1698431365
transform 1 0 33824 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_31_294
timestamp 1698431365
transform 1 0 34272 0 -1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_310
timestamp 1698431365
transform 1 0 36064 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_313
timestamp 1698431365
transform 1 0 36400 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_317
timestamp 1698431365
transform 1 0 36848 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_358
timestamp 1698431365
transform 1 0 41440 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_362
timestamp 1698431365
transform 1 0 41888 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_364
timestamp 1698431365
transform 1 0 42112 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_387
timestamp 1698431365
transform 1 0 44688 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_391
timestamp 1698431365
transform 1 0 45136 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_31_395
timestamp 1698431365
transform 1 0 45584 0 -1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_411
timestamp 1698431365
transform 1 0 47376 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_419
timestamp 1698431365
transform 1 0 48272 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_424
timestamp 1698431365
transform 1 0 48832 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_427
timestamp 1698431365
transform 1 0 49168 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_431
timestamp 1698431365
transform 1 0 49616 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_502
timestamp 1698431365
transform 1 0 57568 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_506
timestamp 1698431365
transform 1 0 58016 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_32_45
timestamp 1698431365
transform 1 0 6384 0 1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_32_61
timestamp 1698431365
transform 1 0 8176 0 1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_69
timestamp 1698431365
transform 1 0 9072 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_32_111
timestamp 1698431365
transform 1 0 13776 0 1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_32_127
timestamp 1698431365
transform 1 0 15568 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_131
timestamp 1698431365
transform 1 0 16016 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_133
timestamp 1698431365
transform 1 0 16240 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_32_164
timestamp 1698431365
transform 1 0 19712 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_170
timestamp 1698431365
transform 1 0 20384 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_32_190
timestamp 1698431365
transform 1 0 22624 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_196
timestamp 1698431365
transform 1 0 23296 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_32_251
timestamp 1698431365
transform 1 0 29456 0 1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_267
timestamp 1698431365
transform 1 0 31248 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_32_297
timestamp 1698431365
transform 1 0 34608 0 1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_367
timestamp 1698431365
transform 1 0 42448 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_371
timestamp 1698431365
transform 1 0 42896 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_375
timestamp 1698431365
transform 1 0 43344 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_435
timestamp 1698431365
transform 1 0 50064 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_464
timestamp 1698431365
transform 1 0 53312 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_6
timestamp 1698431365
transform 1 0 2016 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_33_46
timestamp 1698431365
transform 1 0 6496 0 -1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_33_62
timestamp 1698431365
transform 1 0 8288 0 -1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_33_114
timestamp 1698431365
transform 1 0 14112 0 -1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_33_130
timestamp 1698431365
transform 1 0 15904 0 -1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_172
timestamp 1698431365
transform 1 0 20608 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_176
timestamp 1698431365
transform 1 0 21056 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_180
timestamp 1698431365
transform 1 0 21504 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_33_184
timestamp 1698431365
transform 1 0 21952 0 -1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_192
timestamp 1698431365
transform 1 0 22848 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_196
timestamp 1698431365
transform 1 0 23296 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_202
timestamp 1698431365
transform 1 0 23968 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_33_244
timestamp 1698431365
transform 1 0 28672 0 -1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_260
timestamp 1698431365
transform 1 0 30464 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_264
timestamp 1698431365
transform 1 0 30912 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_33_300
timestamp 1698431365
transform 1 0 34944 0 -1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_308
timestamp 1698431365
transform 1 0 35840 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_312
timestamp 1698431365
transform 1 0 36288 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_314
timestamp 1698431365
transform 1 0 36512 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_317
timestamp 1698431365
transform 1 0 36848 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_321
timestamp 1698431365
transform 1 0 37296 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_323
timestamp 1698431365
transform 1 0 37520 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_326
timestamp 1698431365
transform 1 0 37856 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_354
timestamp 1698431365
transform 1 0 40992 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_370
timestamp 1698431365
transform 1 0 42784 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_409
timestamp 1698431365
transform 1 0 47152 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_413
timestamp 1698431365
transform 1 0 47600 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_416
timestamp 1698431365
transform 1 0 47936 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_424
timestamp 1698431365
transform 1 0 48832 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_484
timestamp 1698431365
transform 1 0 55552 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_488
timestamp 1698431365
transform 1 0 56000 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_508
timestamp 1698431365
transform 1 0 58240 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_45
timestamp 1698431365
transform 1 0 6384 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_34_49
timestamp 1698431365
transform 1 0 6832 0 1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_65
timestamp 1698431365
transform 1 0 8624 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_69
timestamp 1698431365
transform 1 0 9072 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_34_111
timestamp 1698431365
transform 1 0 13776 0 1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_127
timestamp 1698431365
transform 1 0 15568 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_135
timestamp 1698431365
transform 1 0 16464 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_137
timestamp 1698431365
transform 1 0 16688 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_34_168
timestamp 1698431365
transform 1 0 20160 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_34_193
timestamp 1698431365
transform 1 0 22960 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_197
timestamp 1698431365
transform 1 0 23408 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_230
timestamp 1698431365
transform 1 0 27104 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_234
timestamp 1698431365
transform 1 0 27552 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_255
timestamp 1698431365
transform 1 0 29904 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_297
timestamp 1698431365
transform 1 0 34608 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_301
timestamp 1698431365
transform 1 0 35056 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_305
timestamp 1698431365
transform 1 0 35504 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_34_379
timestamp 1698431365
transform 1 0 43792 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_452
timestamp 1698431365
transform 1 0 51968 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_454
timestamp 1698431365
transform 1 0 52192 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_461
timestamp 1698431365
transform 1 0 52976 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_470
timestamp 1698431365
transform 1 0 53984 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_474
timestamp 1698431365
transform 1 0 54432 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_478
timestamp 1698431365
transform 1 0 54880 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_486
timestamp 1698431365
transform 1 0 55776 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_490
timestamp 1698431365
transform 1 0 56224 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_494
timestamp 1698431365
transform 1 0 56672 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_498
timestamp 1698431365
transform 1 0 57120 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_506
timestamp 1698431365
transform 1 0 58016 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_508
timestamp 1698431365
transform 1 0 58240 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_35_110
timestamp 1698431365
transform 1 0 13664 0 -1 40320
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_35_126
timestamp 1698431365
transform 1 0 15456 0 -1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_35_134
timestamp 1698431365
transform 1 0 16352 0 -1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_35_170
timestamp 1698431365
transform 1 0 20384 0 -1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_176
timestamp 1698431365
transform 1 0 21056 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_35_203
timestamp 1698431365
transform 1 0 24080 0 -1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_207
timestamp 1698431365
transform 1 0 24528 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_35_226
timestamp 1698431365
transform 1 0 26656 0 -1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_264
timestamp 1698431365
transform 1 0 30912 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_268
timestamp 1698431365
transform 1 0 31360 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_270
timestamp 1698431365
transform 1 0 31584 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_279
timestamp 1698431365
transform 1 0 32592 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_295
timestamp 1698431365
transform 1 0 34384 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_297
timestamp 1698431365
transform 1 0 34608 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_35_336
timestamp 1698431365
transform 1 0 38976 0 -1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_340
timestamp 1698431365
transform 1 0 39424 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_342
timestamp 1698431365
transform 1 0 39648 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_345
timestamp 1698431365
transform 1 0 39984 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_356
timestamp 1698431365
transform 1 0 41216 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_360
timestamp 1698431365
transform 1 0 41664 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_35_364
timestamp 1698431365
transform 1 0 42112 0 -1 40320
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_380
timestamp 1698431365
transform 1 0 43904 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_383
timestamp 1698431365
transform 1 0 44240 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_387
timestamp 1698431365
transform 1 0 44688 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_391
timestamp 1698431365
transform 1 0 45136 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_415
timestamp 1698431365
transform 1 0 47824 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_417
timestamp 1698431365
transform 1 0 48048 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_447
timestamp 1698431365
transform 1 0 51408 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_449
timestamp 1698431365
transform 1 0 51632 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_35_500
timestamp 1698431365
transform 1 0 57344 0 -1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_508
timestamp 1698431365
transform 1 0 58240 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_41
timestamp 1698431365
transform 1 0 5936 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_36_46
timestamp 1698431365
transform 1 0 6496 0 1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_54
timestamp 1698431365
transform 1 0 7392 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_56
timestamp 1698431365
transform 1 0 7616 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_61
timestamp 1698431365
transform 1 0 8176 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_99
timestamp 1698431365
transform 1 0 12432 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_103
timestamp 1698431365
transform 1 0 12880 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 40320
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_36_123
timestamp 1698431365
transform 1 0 15120 0 1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_131
timestamp 1698431365
transform 1 0 16016 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_162
timestamp 1698431365
transform 1 0 19488 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_164
timestamp 1698431365
transform 1 0 19712 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_167
timestamp 1698431365
transform 1 0 20048 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_179
timestamp 1698431365
transform 1 0 21392 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_228
timestamp 1698431365
transform 1 0 26880 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_36_232
timestamp 1698431365
transform 1 0 27328 0 1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_240
timestamp 1698431365
transform 1 0 28224 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 40320
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_263
timestamp 1698431365
transform 1 0 30800 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_295
timestamp 1698431365
transform 1 0 34384 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_299
timestamp 1698431365
transform 1 0 34832 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_303
timestamp 1698431365
transform 1 0 35280 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_307
timestamp 1698431365
transform 1 0 35728 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_36_349
timestamp 1698431365
transform 1 0 40432 0 1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_357
timestamp 1698431365
transform 1 0 41328 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_361
timestamp 1698431365
transform 1 0 41776 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_364
timestamp 1698431365
transform 1 0 42112 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_368
timestamp 1698431365
transform 1 0 42560 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_371
timestamp 1698431365
transform 1 0 42896 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_375
timestamp 1698431365
transform 1 0 43344 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_379
timestamp 1698431365
transform 1 0 43792 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_391
timestamp 1698431365
transform 1 0 45136 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_36_395
timestamp 1698431365
transform 1 0 45584 0 1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_403
timestamp 1698431365
transform 1 0 46480 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_407
timestamp 1698431365
transform 1 0 46928 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_423
timestamp 1698431365
transform 1 0 48720 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_429
timestamp 1698431365
transform 1 0 49392 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_443
timestamp 1698431365
transform 1 0 50960 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_447
timestamp 1698431365
transform 1 0 51408 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_451
timestamp 1698431365
transform 1 0 51856 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_454
timestamp 1698431365
transform 1 0 52192 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_488
timestamp 1698431365
transform 1 0 56000 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_36_492
timestamp 1698431365
transform 1 0 56448 0 1 40320
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_508
timestamp 1698431365
transform 1 0 58240 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_6
timestamp 1698431365
transform 1 0 2016 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_14
timestamp 1698431365
transform 1 0 2912 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_18
timestamp 1698431365
transform 1 0 3360 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_20
timestamp 1698431365
transform 1 0 3584 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_55
timestamp 1698431365
transform 1 0 7504 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_63
timestamp 1698431365
transform 1 0 8400 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_67
timestamp 1698431365
transform 1 0 8848 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_77
timestamp 1698431365
transform 1 0 9968 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_81
timestamp 1698431365
transform 1 0 10416 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_83
timestamp 1698431365
transform 1 0 10640 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_37_88
timestamp 1698431365
transform 1 0 11200 0 -1 42336
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_37_120
timestamp 1698431365
transform 1 0 14784 0 -1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_158
timestamp 1698431365
transform 1 0 19040 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_205
timestamp 1698431365
transform 1 0 24304 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_207
timestamp 1698431365
transform 1 0 24528 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_242
timestamp 1698431365
transform 1 0 28448 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_246
timestamp 1698431365
transform 1 0 28896 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_267
timestamp 1698431365
transform 1 0 31248 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_271
timestamp 1698431365
transform 1 0 31696 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_288
timestamp 1698431365
transform 1 0 33600 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_290
timestamp 1698431365
transform 1 0 33824 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_293
timestamp 1698431365
transform 1 0 34160 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_297
timestamp 1698431365
transform 1 0 34608 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_402
timestamp 1698431365
transform 1 0 46368 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_406
timestamp 1698431365
transform 1 0 46816 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_414
timestamp 1698431365
transform 1 0 47712 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_418
timestamp 1698431365
transform 1 0 48160 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_424
timestamp 1698431365
transform 1 0 48832 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_427
timestamp 1698431365
transform 1 0 49168 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_431
timestamp 1698431365
transform 1 0 49616 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_435
timestamp 1698431365
transform 1 0 50064 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_437
timestamp 1698431365
transform 1 0 50288 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_440
timestamp 1698431365
transform 1 0 50624 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_444
timestamp 1698431365
transform 1 0 51072 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_474
timestamp 1698431365
transform 1 0 54432 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_476
timestamp 1698431365
transform 1 0 54656 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_496
timestamp 1698431365
transform 1 0 56896 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_500
timestamp 1698431365
transform 1 0 57344 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_504
timestamp 1698431365
transform 1 0 57792 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_49
timestamp 1698431365
transform 1 0 6832 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_51
timestamp 1698431365
transform 1 0 7056 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_38_86
timestamp 1698431365
transform 1 0 10976 0 1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_102
timestamp 1698431365
transform 1 0 12768 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_38_139
timestamp 1698431365
transform 1 0 16912 0 1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_38_155
timestamp 1698431365
transform 1 0 18704 0 1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_163
timestamp 1698431365
transform 1 0 19600 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_167
timestamp 1698431365
transform 1 0 20048 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_169
timestamp 1698431365
transform 1 0 20272 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_172
timestamp 1698431365
transform 1 0 20608 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_183
timestamp 1698431365
transform 1 0 21840 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_187
timestamp 1698431365
transform 1 0 22288 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_191
timestamp 1698431365
transform 1 0 22736 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_224
timestamp 1698431365
transform 1 0 26432 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_226
timestamp 1698431365
transform 1 0 26656 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_229
timestamp 1698431365
transform 1 0 26992 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_233
timestamp 1698431365
transform 1 0 27440 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_237
timestamp 1698431365
transform 1 0 27888 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_38_293
timestamp 1698431365
transform 1 0 34160 0 1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_309
timestamp 1698431365
transform 1 0 35952 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_321
timestamp 1698431365
transform 1 0 37296 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_329
timestamp 1698431365
transform 1 0 38192 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_331
timestamp 1698431365
transform 1 0 38416 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_383
timestamp 1698431365
transform 1 0 44240 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_400
timestamp 1698431365
transform 1 0 46144 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_404
timestamp 1698431365
transform 1 0 46592 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_408
timestamp 1698431365
transform 1 0 47040 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_412
timestamp 1698431365
transform 1 0 47488 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_416
timestamp 1698431365
transform 1 0 47936 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_420
timestamp 1698431365
transform 1 0 48384 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_424
timestamp 1698431365
transform 1 0 48832 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_428
timestamp 1698431365
transform 1 0 49280 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_434
timestamp 1698431365
transform 1 0 49952 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_442
timestamp 1698431365
transform 1 0 50848 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_446
timestamp 1698431365
transform 1 0 51296 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_450
timestamp 1698431365
transform 1 0 51744 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_454
timestamp 1698431365
transform 1 0 52192 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_490
timestamp 1698431365
transform 1 0 56224 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_494
timestamp 1698431365
transform 1 0 56672 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_498
timestamp 1698431365
transform 1 0 57120 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_502
timestamp 1698431365
transform 1 0 57568 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_506
timestamp 1698431365
transform 1 0 58016 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_508
timestamp 1698431365
transform 1 0 58240 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 44352
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 44352
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 44352
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_158
timestamp 1698431365
transform 1 0 19040 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_162
timestamp 1698431365
transform 1 0 19488 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_164
timestamp 1698431365
transform 1 0 19712 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_167
timestamp 1698431365
transform 1 0 20048 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_171
timestamp 1698431365
transform 1 0 20496 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_175
timestamp 1698431365
transform 1 0 20944 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_179
timestamp 1698431365
transform 1 0 21392 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_39_183
timestamp 1698431365
transform 1 0 21840 0 -1 44352
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_199
timestamp 1698431365
transform 1 0 23632 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_203
timestamp 1698431365
transform 1 0 24080 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_216
timestamp 1698431365
transform 1 0 25536 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_219
timestamp 1698431365
transform 1 0 25872 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_39_223
timestamp 1698431365
transform 1 0 26320 0 -1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_233
timestamp 1698431365
transform 1 0 27440 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_239
timestamp 1698431365
transform 1 0 28112 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_243
timestamp 1698431365
transform 1 0 28560 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_273
timestamp 1698431365
transform 1 0 31920 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_277
timestamp 1698431365
transform 1 0 32368 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_290
timestamp 1698431365
transform 1 0 33824 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_292
timestamp 1698431365
transform 1 0 34048 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_39_295
timestamp 1698431365
transform 1 0 34384 0 -1 44352
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_39_311
timestamp 1698431365
transform 1 0 36176 0 -1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_319
timestamp 1698431365
transform 1 0 37072 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_322
timestamp 1698431365
transform 1 0 37408 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_326
timestamp 1698431365
transform 1 0 37856 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_330
timestamp 1698431365
transform 1 0 38304 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_334
timestamp 1698431365
transform 1 0 38752 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_338
timestamp 1698431365
transform 1 0 39200 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_342
timestamp 1698431365
transform 1 0 39648 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_356
timestamp 1698431365
transform 1 0 41216 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_405
timestamp 1698431365
transform 1 0 46704 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_456
timestamp 1698431365
transform 1 0 52416 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_458
timestamp 1698431365
transform 1 0 52640 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_496
timestamp 1698431365
transform 1 0 56896 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_39_500
timestamp 1698431365
transform 1 0 57344 0 -1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_508
timestamp 1698431365
transform 1 0 58240 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 44352
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_139
timestamp 1698431365
transform 1 0 16912 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_40_255
timestamp 1698431365
transform 1 0 29904 0 1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_290
timestamp 1698431365
transform 1 0 33824 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_294
timestamp 1698431365
transform 1 0 34272 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_321
timestamp 1698431365
transform 1 0 37296 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_395
timestamp 1698431365
transform 1 0 45584 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_397
timestamp 1698431365
transform 1 0 45808 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_453
timestamp 1698431365
transform 1 0 52080 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_40_488
timestamp 1698431365
transform 1 0 56000 0 1 44352
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_40_504
timestamp 1698431365
transform 1 0 57792 0 1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_508
timestamp 1698431365
transform 1 0 58240 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 46368
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 46368
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_188
timestamp 1698431365
transform 1 0 22400 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_192
timestamp 1698431365
transform 1 0 22848 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_198
timestamp 1698431365
transform 1 0 23520 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_202
timestamp 1698431365
transform 1 0 23968 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_233
timestamp 1698431365
transform 1 0 27440 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_278
timestamp 1698431365
transform 1 0 32480 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_313
timestamp 1698431365
transform 1 0 36400 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_317
timestamp 1698431365
transform 1 0 36848 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_343
timestamp 1698431365
transform 1 0 39760 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_345
timestamp 1698431365
transform 1 0 39984 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_348
timestamp 1698431365
transform 1 0 40320 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_398
timestamp 1698431365
transform 1 0 45920 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_402
timestamp 1698431365
transform 1 0 46368 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_406
timestamp 1698431365
transform 1 0 46816 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_41_410
timestamp 1698431365
transform 1 0 47264 0 -1 46368
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_453
timestamp 1698431365
transform 1 0 52080 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_457
timestamp 1698431365
transform 1 0 52528 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_476
timestamp 1698431365
transform 1 0 54656 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_480
timestamp 1698431365
transform 1 0 55104 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_484
timestamp 1698431365
transform 1 0 55552 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_488
timestamp 1698431365
transform 1 0 56000 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 46368
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 46368
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 46368
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 46368
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_139
timestamp 1698431365
transform 1 0 16912 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_183
timestamp 1698431365
transform 1 0 21840 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_226
timestamp 1698431365
transform 1 0 26656 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_42_230
timestamp 1698431365
transform 1 0 27104 0 1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_233
timestamp 1698431365
transform 1 0 27440 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_237
timestamp 1698431365
transform 1 0 27888 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_309
timestamp 1698431365
transform 1 0 35952 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_321
timestamp 1698431365
transform 1 0 37296 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_329
timestamp 1698431365
transform 1 0 38192 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_333
timestamp 1698431365
transform 1 0 38640 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_42_335
timestamp 1698431365
transform 1 0 38864 0 1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_367
timestamp 1698431365
transform 1 0 42448 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_371
timestamp 1698431365
transform 1 0 42896 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_375
timestamp 1698431365
transform 1 0 43344 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_379
timestamp 1698431365
transform 1 0 43792 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_383
timestamp 1698431365
transform 1 0 44240 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_391
timestamp 1698431365
transform 1 0 45136 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_461
timestamp 1698431365
transform 1 0 52976 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_465
timestamp 1698431365
transform 1 0 53424 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_469
timestamp 1698431365
transform 1 0 53872 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_42_473
timestamp 1698431365
transform 1 0 54320 0 1 46368
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_505
timestamp 1698431365
transform 1 0 57904 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_196
timestamp 1698431365
transform 1 0 23296 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_200
timestamp 1698431365
transform 1 0 23744 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_204
timestamp 1698431365
transform 1 0 24192 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_222
timestamp 1698431365
transform 1 0 26208 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_226
timestamp 1698431365
transform 1 0 26656 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_230
timestamp 1698431365
transform 1 0 27104 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_269
timestamp 1698431365
transform 1 0 31472 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_273
timestamp 1698431365
transform 1 0 31920 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_43_339
timestamp 1698431365
transform 1 0 39312 0 -1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_347
timestamp 1698431365
transform 1 0 40208 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_356
timestamp 1698431365
transform 1 0 41216 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_360
timestamp 1698431365
transform 1 0 41664 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_364
timestamp 1698431365
transform 1 0 42112 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_368
timestamp 1698431365
transform 1 0 42560 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_372
timestamp 1698431365
transform 1 0 43008 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_376
timestamp 1698431365
transform 1 0 43456 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_380
timestamp 1698431365
transform 1 0 43904 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_384
timestamp 1698431365
transform 1 0 44352 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_388
timestamp 1698431365
transform 1 0 44800 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_390
timestamp 1698431365
transform 1 0 45024 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_43_393
timestamp 1698431365
transform 1 0 45360 0 -1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_43_409
timestamp 1698431365
transform 1 0 47152 0 -1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_417
timestamp 1698431365
transform 1 0 48048 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_419
timestamp 1698431365
transform 1 0 48272 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_430
timestamp 1698431365
transform 1 0 49504 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_434
timestamp 1698431365
transform 1 0 49952 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_438
timestamp 1698431365
transform 1 0 50400 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_43_442
timestamp 1698431365
transform 1 0 50848 0 -1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_450
timestamp 1698431365
transform 1 0 51744 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_452
timestamp 1698431365
transform 1 0 51968 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_455
timestamp 1698431365
transform 1 0 52304 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_459
timestamp 1698431365
transform 1 0 52752 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_463
timestamp 1698431365
transform 1 0 53200 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_43_467
timestamp 1698431365
transform 1 0 53648 0 -1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_483
timestamp 1698431365
transform 1 0 55440 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_487
timestamp 1698431365
transform 1 0 55888 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_489
timestamp 1698431365
transform 1 0 56112 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_508
timestamp 1698431365
transform 1 0 58240 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 48384
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_181
timestamp 1698431365
transform 1 0 21616 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_185
timestamp 1698431365
transform 1 0 22064 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_44_189
timestamp 1698431365
transform 1 0 22512 0 1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_197
timestamp 1698431365
transform 1 0 23408 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_44_229
timestamp 1698431365
transform 1 0 26992 0 1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_44_263
timestamp 1698431365
transform 1 0 30800 0 1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_271
timestamp 1698431365
transform 1 0 31696 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_273
timestamp 1698431365
transform 1 0 31920 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_276
timestamp 1698431365
transform 1 0 32256 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_280
timestamp 1698431365
transform 1 0 32704 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_282
timestamp 1698431365
transform 1 0 32928 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_285
timestamp 1698431365
transform 1 0 33264 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_44_289
timestamp 1698431365
transform 1 0 33712 0 1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_44_306
timestamp 1698431365
transform 1 0 35616 0 1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_314
timestamp 1698431365
transform 1 0 36512 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_325
timestamp 1698431365
transform 1 0 37744 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_329
timestamp 1698431365
transform 1 0 38192 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_332
timestamp 1698431365
transform 1 0 38528 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_336
timestamp 1698431365
transform 1 0 38976 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_366
timestamp 1698431365
transform 1 0 42336 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_370
timestamp 1698431365
transform 1 0 42784 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_44_374
timestamp 1698431365
transform 1 0 43232 0 1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_382
timestamp 1698431365
transform 1 0 44128 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698431365
transform 1 0 51856 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 48384
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_44_489
timestamp 1698431365
transform 1 0 56112 0 1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_505
timestamp 1698431365
transform 1 0 57904 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_416
timestamp 1698431365
transform 1 0 47936 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698431365
transform 1 0 55776 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 50400
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_45_508
timestamp 1698431365
transform 1 0 58240 0 -1 50400
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 50400
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 50400
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698431365
transform 1 0 44016 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_451
timestamp 1698431365
transform 1 0 51856 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 50400
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_46_489
timestamp 1698431365
transform 1 0 56112 0 1 50400
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_505
timestamp 1698431365
transform 1 0 57904 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698431365
transform 1 0 55776 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 52416
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 52416
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 52416
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 52416
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698431365
transform 1 0 51856 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 52416
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_48_489
timestamp 1698431365
transform 1 0 56112 0 1 52416
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_505
timestamp 1698431365
transform 1 0 57904 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 54432
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_49_18
timestamp 1698431365
transform 1 0 3360 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_49_20
timestamp 1698431365
transform 1 0 3584 0 -1 54432
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_49_25
timestamp 1698431365
transform 1 0 4144 0 -1 54432
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_49_57
timestamp 1698431365
transform 1 0 7728 0 -1 54432
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_65
timestamp 1698431365
transform 1 0 8624 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_49_69
timestamp 1698431365
transform 1 0 9072 0 -1 54432
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_346
timestamp 1698431365
transform 1 0 40096 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_416
timestamp 1698431365
transform 1 0 47936 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 54432
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 54432
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 54432
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 54432
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698431365
transform 1 0 20496 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698431365
transform 1 0 51856 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 54432
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_50_489
timestamp 1698431365
transform 1 0 56112 0 1 54432
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_505
timestamp 1698431365
transform 1 0 57904 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_36
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_104
timestamp 1698431365
transform 1 0 12992 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_172
timestamp 1698431365
transform 1 0 20608 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_240
timestamp 1698431365
transform 1 0 28224 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_274
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_308
timestamp 1698431365
transform 1 0 35840 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_342
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_376
timestamp 1698431365
transform 1 0 43456 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_410
timestamp 1698431365
transform 1 0 47264 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_444
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_51_478
timestamp 1698431365
transform 1 0 54880 0 -1 56448
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_51_494
timestamp 1698431365
transform 1 0 56672 0 -1 56448
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_51_502
timestamp 1698431365
transform 1 0 57568 0 -1 56448
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_51_506
timestamp 1698431365
transform 1 0 58016 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 56448
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_0_Left_52 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 4032
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 4032
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_1_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_2_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_3_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_4_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_5_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_6_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_7_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_8_Left_60
timestamp 1698431365
transform 1 0 1344 0 1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_9_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_10_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_11_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_12_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_13_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_14_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_15_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_16_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_17_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_18_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_19_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_20_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_21_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_22_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_23_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_24_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_25_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_26_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_27_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_28_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_29_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_30_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_31_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 36288
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 36288
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_32_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 36288
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 36288
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_33_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 38304
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 38304
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_34_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 38304
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 38304
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_35_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 40320
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 40320
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_36_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 40320
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 40320
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_37_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_38_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_39_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 44352
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 44352
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_40_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 44352
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 44352
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_41_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 46368
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 46368
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_42_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 46368
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 46368
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_43_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 48384
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 48384
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_44_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 48384
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 48384
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_45_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 50400
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 50400
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_46_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 50400
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 50400
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_47_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 52416
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 52416
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_48_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 52416
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 52416
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_49_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 54432
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 54432
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_50_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 54432
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 54432
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_51_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtp_2  ro_inst.clock_gate
timestamp 1698431365
transform 1 0 10192 0 -1 32256
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.clock_gate_inv
timestamp 1698431365
transform -1 0 12544 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[1\].div_flop_inv
timestamp 1698431365
transform -1 0 13776 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[1\].div_flop
timestamp 1698431365
transform 1 0 11424 0 -1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[2\].div_flop_inv
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[2\].div_flop
timestamp 1698431365
transform 1 0 11648 0 -1 26208
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[3\].div_flop
timestamp 1698431365
transform 1 0 13328 0 1 26208
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[3\].div_flop_inv
timestamp 1698431365
transform -1 0 13776 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[4\].div_flop
timestamp 1698431365
transform -1 0 13104 0 1 26208
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[4\].div_flop_inv
timestamp 1698431365
transform -1 0 11648 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[5\].div_flop_inv
timestamp 1698431365
transform -1 0 11200 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[5\].div_flop
timestamp 1698431365
transform 1 0 9520 0 1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[6\].div_flop_inv
timestamp 1698431365
transform 1 0 8624 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[6\].div_flop
timestamp 1698431365
transform -1 0 9520 0 1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[7\].div_flop_inv
timestamp 1698431365
transform -1 0 8400 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[7\].div_flop
timestamp 1698431365
transform -1 0 9184 0 -1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[8\].div_flop
timestamp 1698431365
transform -1 0 7952 0 -1 26208
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[8\].div_flop_inv
timestamp 1698431365
transform 1 0 5488 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[9\].div_flop_inv
timestamp 1698431365
transform 1 0 2912 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[9\].div_flop
timestamp 1698431365
transform -1 0 5600 0 -1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[10\].div_flop_inv
timestamp 1698431365
transform -1 0 3808 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[10\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 22176
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[11\].div_flop_inv
timestamp 1698431365
transform -1 0 4256 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[11\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[12\].div_flop_inv
timestamp 1698431365
transform -1 0 2912 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[12\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 26208
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[13\].div_flop_inv
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[13\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[14\].div_flop_inv
timestamp 1698431365
transform -1 0 3472 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[14\].div_flop
timestamp 1698431365
transform -1 0 6496 0 -1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[15\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 30240
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[15\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[16\].div_flop
timestamp 1698431365
transform 1 0 5488 0 1 30240
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[16\].div_flop_inv
timestamp 1698431365
transform -1 0 7616 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[17\].div_flop_inv
timestamp 1698431365
transform 1 0 5936 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[17\].div_flop
timestamp 1698431365
transform -1 0 7056 0 -1 30240
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[18\].div_flop_inv
timestamp 1698431365
transform 1 0 5488 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[18\].div_flop
timestamp 1698431365
transform -1 0 7168 0 -1 32256
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[19\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[19\].div_flop
timestamp 1698431365
transform -1 0 7056 0 -1 34272
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[20\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[20\].div_flop
timestamp 1698431365
transform 1 0 3248 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[21\].div_flop
timestamp 1698431365
transform 1 0 2912 0 -1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[21\].div_flop_inv
timestamp 1698431365
transform -1 0 6384 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[22\].div_flop
timestamp 1698431365
transform -1 0 5264 0 1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[22\].div_flop_inv
timestamp 1698431365
transform 1 0 2464 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[23\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[23\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[24\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[24\].div_flop
timestamp 1698431365
transform 1 0 2016 0 -1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[25\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[25\].div_flop_inv
timestamp 1698431365
transform -1 0 6384 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[26\].div_flop
timestamp 1698431365
transform 1 0 3920 0 -1 42336
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[26\].div_flop_inv
timestamp 1698431365
transform -1 0 6496 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[27\].div_flop_inv
timestamp 1698431365
transform -1 0 8176 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[27\].div_flop
timestamp 1698431365
transform 1 0 5600 0 -1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[28\].div_flop
timestamp 1698431365
transform 1 0 7392 0 1 42336
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[28\].div_flop_inv
timestamp 1698431365
transform -1 0 9968 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[29\].div_flop_inv
timestamp 1698431365
transform -1 0 11200 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[29\].div_flop
timestamp 1698431365
transform 1 0 8848 0 1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[30\].div_flop_inv
timestamp 1698431365
transform -1 0 13664 0 -1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[30\].div_flop
timestamp 1698431365
transform 1 0 9632 0 -1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[31\].div_flop_inv
timestamp 1698431365
transform -1 0 13776 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[31\].div_flop
timestamp 1698431365
transform 1 0 9520 0 1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[32\].div_flop
timestamp 1698431365
transform 1 0 10080 0 -1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[32\].div_flop_inv
timestamp 1698431365
transform -1 0 14112 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[33\].div_flop
timestamp 1698431365
transform 1 0 9520 0 1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[33\].div_flop_inv
timestamp 1698431365
transform -1 0 13776 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[34\].div_flop
timestamp 1698431365
transform 1 0 11200 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[34\].div_flop_inv
timestamp 1698431365
transform -1 0 13776 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  ro_inst.ring_osc_0
timestamp 1698431365
transform 1 0 11760 0 -1 34272
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.ring_osc_1
timestamp 1698431365
transform -1 0 14224 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.ring_osc_2
timestamp 1698431365
transform 1 0 11536 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_1  ro_inst.sig_cmp
timestamp 1698431365
transform -1 0 11536 0 -1 30240
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_1  ro_inst.sig_latch
timestamp 1698431365
transform 1 0 9744 0 1 30240
box -86 -90 2326 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.slow_clock_inv
timestamp 1698431365
transform 1 0 8736 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_104 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 8960 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 12768 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 16576 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 20384 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 24192 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 28000 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 31808 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 35616 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 39424 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 43232 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 47040 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 50848 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 54656 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_118
timestamp 1698431365
transform 1 0 9184 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_119
timestamp 1698431365
transform 1 0 17024 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_120
timestamp 1698431365
transform 1 0 24864 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_121
timestamp 1698431365
transform 1 0 32704 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_122
timestamp 1698431365
transform 1 0 40544 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_123
timestamp 1698431365
transform 1 0 48384 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_124
timestamp 1698431365
transform 1 0 56224 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_125
timestamp 1698431365
transform 1 0 5264 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_126
timestamp 1698431365
transform 1 0 13104 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 20944 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_128
timestamp 1698431365
transform 1 0 28784 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_129
timestamp 1698431365
transform 1 0 36624 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_130
timestamp 1698431365
transform 1 0 44464 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_131
timestamp 1698431365
transform 1 0 52304 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_132
timestamp 1698431365
transform 1 0 9184 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_133
timestamp 1698431365
transform 1 0 17024 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_134
timestamp 1698431365
transform 1 0 24864 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_135
timestamp 1698431365
transform 1 0 32704 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_136
timestamp 1698431365
transform 1 0 40544 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_137
timestamp 1698431365
transform 1 0 48384 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_138
timestamp 1698431365
transform 1 0 56224 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_139
timestamp 1698431365
transform 1 0 5264 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_140
timestamp 1698431365
transform 1 0 13104 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_141
timestamp 1698431365
transform 1 0 20944 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_142
timestamp 1698431365
transform 1 0 28784 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_143
timestamp 1698431365
transform 1 0 36624 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_144
timestamp 1698431365
transform 1 0 44464 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_145
timestamp 1698431365
transform 1 0 52304 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_146
timestamp 1698431365
transform 1 0 9184 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_147
timestamp 1698431365
transform 1 0 17024 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_148
timestamp 1698431365
transform 1 0 24864 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_149
timestamp 1698431365
transform 1 0 32704 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_150
timestamp 1698431365
transform 1 0 40544 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_151
timestamp 1698431365
transform 1 0 48384 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_152
timestamp 1698431365
transform 1 0 56224 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_153
timestamp 1698431365
transform 1 0 5264 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_154
timestamp 1698431365
transform 1 0 13104 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_155
timestamp 1698431365
transform 1 0 20944 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_156
timestamp 1698431365
transform 1 0 28784 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_157
timestamp 1698431365
transform 1 0 36624 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_158
timestamp 1698431365
transform 1 0 44464 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_159
timestamp 1698431365
transform 1 0 52304 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_160
timestamp 1698431365
transform 1 0 9184 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_161
timestamp 1698431365
transform 1 0 17024 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_162
timestamp 1698431365
transform 1 0 24864 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_163
timestamp 1698431365
transform 1 0 32704 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_164
timestamp 1698431365
transform 1 0 40544 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_165
timestamp 1698431365
transform 1 0 48384 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_166
timestamp 1698431365
transform 1 0 56224 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_167
timestamp 1698431365
transform 1 0 5264 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_168
timestamp 1698431365
transform 1 0 13104 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_169
timestamp 1698431365
transform 1 0 20944 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_170
timestamp 1698431365
transform 1 0 28784 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_171
timestamp 1698431365
transform 1 0 36624 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_172
timestamp 1698431365
transform 1 0 44464 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_173
timestamp 1698431365
transform 1 0 52304 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_174
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_175
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_176
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_177
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_178
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_179
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_180
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_181
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_182
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_183
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_184
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_185
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_186
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_187
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_188
timestamp 1698431365
transform 1 0 9184 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_189
timestamp 1698431365
transform 1 0 17024 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_190
timestamp 1698431365
transform 1 0 24864 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_191
timestamp 1698431365
transform 1 0 32704 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_192
timestamp 1698431365
transform 1 0 40544 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_193
timestamp 1698431365
transform 1 0 48384 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_194
timestamp 1698431365
transform 1 0 56224 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_195
timestamp 1698431365
transform 1 0 5264 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_196
timestamp 1698431365
transform 1 0 13104 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_197
timestamp 1698431365
transform 1 0 20944 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_198
timestamp 1698431365
transform 1 0 28784 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_199
timestamp 1698431365
transform 1 0 36624 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_200
timestamp 1698431365
transform 1 0 44464 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_201
timestamp 1698431365
transform 1 0 52304 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_202
timestamp 1698431365
transform 1 0 9184 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_203
timestamp 1698431365
transform 1 0 17024 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_204
timestamp 1698431365
transform 1 0 24864 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_205
timestamp 1698431365
transform 1 0 32704 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_206
timestamp 1698431365
transform 1 0 40544 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_207
timestamp 1698431365
transform 1 0 48384 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_208
timestamp 1698431365
transform 1 0 56224 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_209
timestamp 1698431365
transform 1 0 5264 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_210
timestamp 1698431365
transform 1 0 13104 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_211
timestamp 1698431365
transform 1 0 20944 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_212
timestamp 1698431365
transform 1 0 28784 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_213
timestamp 1698431365
transform 1 0 36624 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_214
timestamp 1698431365
transform 1 0 44464 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_215
timestamp 1698431365
transform 1 0 52304 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_216
timestamp 1698431365
transform 1 0 9184 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_217
timestamp 1698431365
transform 1 0 17024 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_218
timestamp 1698431365
transform 1 0 24864 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_219
timestamp 1698431365
transform 1 0 32704 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_220
timestamp 1698431365
transform 1 0 40544 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_221
timestamp 1698431365
transform 1 0 48384 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_222
timestamp 1698431365
transform 1 0 56224 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_223
timestamp 1698431365
transform 1 0 5264 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_224
timestamp 1698431365
transform 1 0 13104 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_225
timestamp 1698431365
transform 1 0 20944 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_226
timestamp 1698431365
transform 1 0 28784 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_227
timestamp 1698431365
transform 1 0 36624 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_228
timestamp 1698431365
transform 1 0 44464 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_229
timestamp 1698431365
transform 1 0 52304 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_230
timestamp 1698431365
transform 1 0 9184 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_231
timestamp 1698431365
transform 1 0 17024 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_232
timestamp 1698431365
transform 1 0 24864 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_233
timestamp 1698431365
transform 1 0 32704 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_234
timestamp 1698431365
transform 1 0 40544 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_235
timestamp 1698431365
transform 1 0 48384 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_236
timestamp 1698431365
transform 1 0 56224 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_237
timestamp 1698431365
transform 1 0 5264 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_238
timestamp 1698431365
transform 1 0 13104 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_239
timestamp 1698431365
transform 1 0 20944 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_240
timestamp 1698431365
transform 1 0 28784 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_241
timestamp 1698431365
transform 1 0 36624 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_242
timestamp 1698431365
transform 1 0 44464 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_243
timestamp 1698431365
transform 1 0 52304 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_244
timestamp 1698431365
transform 1 0 9184 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_245
timestamp 1698431365
transform 1 0 17024 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_246
timestamp 1698431365
transform 1 0 24864 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_247
timestamp 1698431365
transform 1 0 32704 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_248
timestamp 1698431365
transform 1 0 40544 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_249
timestamp 1698431365
transform 1 0 48384 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_250
timestamp 1698431365
transform 1 0 56224 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_251
timestamp 1698431365
transform 1 0 5264 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_252
timestamp 1698431365
transform 1 0 13104 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_253
timestamp 1698431365
transform 1 0 20944 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_254
timestamp 1698431365
transform 1 0 28784 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_255
timestamp 1698431365
transform 1 0 36624 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_256
timestamp 1698431365
transform 1 0 44464 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_257
timestamp 1698431365
transform 1 0 52304 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_258
timestamp 1698431365
transform 1 0 9184 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_259
timestamp 1698431365
transform 1 0 17024 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_260
timestamp 1698431365
transform 1 0 24864 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_261
timestamp 1698431365
transform 1 0 32704 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_262
timestamp 1698431365
transform 1 0 40544 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_263
timestamp 1698431365
transform 1 0 48384 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_264
timestamp 1698431365
transform 1 0 56224 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_265
timestamp 1698431365
transform 1 0 5264 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_266
timestamp 1698431365
transform 1 0 13104 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_267
timestamp 1698431365
transform 1 0 20944 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_268
timestamp 1698431365
transform 1 0 28784 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_269
timestamp 1698431365
transform 1 0 36624 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_270
timestamp 1698431365
transform 1 0 44464 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_271
timestamp 1698431365
transform 1 0 52304 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_272
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_273
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_274
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_275
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_276
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_277
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_278
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_279
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_280
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_281
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_282
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_283
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_284
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_285
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_286
timestamp 1698431365
transform 1 0 9184 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_287
timestamp 1698431365
transform 1 0 17024 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_288
timestamp 1698431365
transform 1 0 24864 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_289
timestamp 1698431365
transform 1 0 32704 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_290
timestamp 1698431365
transform 1 0 40544 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_291
timestamp 1698431365
transform 1 0 48384 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_292
timestamp 1698431365
transform 1 0 56224 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_293
timestamp 1698431365
transform 1 0 5264 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_294
timestamp 1698431365
transform 1 0 13104 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_295
timestamp 1698431365
transform 1 0 20944 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_296
timestamp 1698431365
transform 1 0 28784 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_297
timestamp 1698431365
transform 1 0 36624 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_298
timestamp 1698431365
transform 1 0 44464 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_299
timestamp 1698431365
transform 1 0 52304 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_300
timestamp 1698431365
transform 1 0 9184 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_301
timestamp 1698431365
transform 1 0 17024 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_302
timestamp 1698431365
transform 1 0 24864 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_303
timestamp 1698431365
transform 1 0 32704 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_304
timestamp 1698431365
transform 1 0 40544 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_305
timestamp 1698431365
transform 1 0 48384 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_306
timestamp 1698431365
transform 1 0 56224 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_307
timestamp 1698431365
transform 1 0 5264 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_308
timestamp 1698431365
transform 1 0 13104 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_309
timestamp 1698431365
transform 1 0 20944 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_310
timestamp 1698431365
transform 1 0 28784 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_311
timestamp 1698431365
transform 1 0 36624 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_312
timestamp 1698431365
transform 1 0 44464 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_313
timestamp 1698431365
transform 1 0 52304 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_314
timestamp 1698431365
transform 1 0 9184 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_315
timestamp 1698431365
transform 1 0 17024 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_316
timestamp 1698431365
transform 1 0 24864 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_317
timestamp 1698431365
transform 1 0 32704 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_318
timestamp 1698431365
transform 1 0 40544 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_319
timestamp 1698431365
transform 1 0 48384 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_320
timestamp 1698431365
transform 1 0 56224 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_321
timestamp 1698431365
transform 1 0 5264 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_322
timestamp 1698431365
transform 1 0 13104 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_323
timestamp 1698431365
transform 1 0 20944 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_324
timestamp 1698431365
transform 1 0 28784 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_325
timestamp 1698431365
transform 1 0 36624 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_326
timestamp 1698431365
transform 1 0 44464 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_327
timestamp 1698431365
transform 1 0 52304 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_328
timestamp 1698431365
transform 1 0 9184 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_329
timestamp 1698431365
transform 1 0 17024 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_330
timestamp 1698431365
transform 1 0 24864 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_331
timestamp 1698431365
transform 1 0 32704 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_332
timestamp 1698431365
transform 1 0 40544 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_333
timestamp 1698431365
transform 1 0 48384 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_334
timestamp 1698431365
transform 1 0 56224 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_335
timestamp 1698431365
transform 1 0 5264 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_336
timestamp 1698431365
transform 1 0 13104 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_337
timestamp 1698431365
transform 1 0 20944 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_338
timestamp 1698431365
transform 1 0 28784 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_339
timestamp 1698431365
transform 1 0 36624 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_340
timestamp 1698431365
transform 1 0 44464 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_341
timestamp 1698431365
transform 1 0 52304 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_342
timestamp 1698431365
transform 1 0 9184 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_343
timestamp 1698431365
transform 1 0 17024 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_344
timestamp 1698431365
transform 1 0 24864 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_345
timestamp 1698431365
transform 1 0 32704 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_346
timestamp 1698431365
transform 1 0 40544 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_347
timestamp 1698431365
transform 1 0 48384 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_348
timestamp 1698431365
transform 1 0 56224 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_349
timestamp 1698431365
transform 1 0 5264 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_350
timestamp 1698431365
transform 1 0 13104 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_351
timestamp 1698431365
transform 1 0 20944 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_352
timestamp 1698431365
transform 1 0 28784 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_353
timestamp 1698431365
transform 1 0 36624 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_354
timestamp 1698431365
transform 1 0 44464 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_355
timestamp 1698431365
transform 1 0 52304 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_356
timestamp 1698431365
transform 1 0 9184 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_357
timestamp 1698431365
transform 1 0 17024 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_358
timestamp 1698431365
transform 1 0 24864 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_359
timestamp 1698431365
transform 1 0 32704 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_360
timestamp 1698431365
transform 1 0 40544 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_361
timestamp 1698431365
transform 1 0 48384 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_362
timestamp 1698431365
transform 1 0 56224 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_363
timestamp 1698431365
transform 1 0 5264 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_364
timestamp 1698431365
transform 1 0 13104 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_365
timestamp 1698431365
transform 1 0 20944 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_366
timestamp 1698431365
transform 1 0 28784 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_367
timestamp 1698431365
transform 1 0 36624 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_368
timestamp 1698431365
transform 1 0 44464 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_369
timestamp 1698431365
transform 1 0 52304 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_370
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_371
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_372
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_373
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_374
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_375
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_376
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_377
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_378
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_379
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_380
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_381
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_382
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_383
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_384
timestamp 1698431365
transform 1 0 9184 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_385
timestamp 1698431365
transform 1 0 17024 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_386
timestamp 1698431365
transform 1 0 24864 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_387
timestamp 1698431365
transform 1 0 32704 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_388
timestamp 1698431365
transform 1 0 40544 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_389
timestamp 1698431365
transform 1 0 48384 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_390
timestamp 1698431365
transform 1 0 56224 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_391
timestamp 1698431365
transform 1 0 5264 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_392
timestamp 1698431365
transform 1 0 13104 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_393
timestamp 1698431365
transform 1 0 20944 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_394
timestamp 1698431365
transform 1 0 28784 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_395
timestamp 1698431365
transform 1 0 36624 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_396
timestamp 1698431365
transform 1 0 44464 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_397
timestamp 1698431365
transform 1 0 52304 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_398
timestamp 1698431365
transform 1 0 9184 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_399
timestamp 1698431365
transform 1 0 17024 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_400
timestamp 1698431365
transform 1 0 24864 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_401
timestamp 1698431365
transform 1 0 32704 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_402
timestamp 1698431365
transform 1 0 40544 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_403
timestamp 1698431365
transform 1 0 48384 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_404
timestamp 1698431365
transform 1 0 56224 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_405
timestamp 1698431365
transform 1 0 5264 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_406
timestamp 1698431365
transform 1 0 13104 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_407
timestamp 1698431365
transform 1 0 20944 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_408
timestamp 1698431365
transform 1 0 28784 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_409
timestamp 1698431365
transform 1 0 36624 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_410
timestamp 1698431365
transform 1 0 44464 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_411
timestamp 1698431365
transform 1 0 52304 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_412
timestamp 1698431365
transform 1 0 9184 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_413
timestamp 1698431365
transform 1 0 17024 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_414
timestamp 1698431365
transform 1 0 24864 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_415
timestamp 1698431365
transform 1 0 32704 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_416
timestamp 1698431365
transform 1 0 40544 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_417
timestamp 1698431365
transform 1 0 48384 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_418
timestamp 1698431365
transform 1 0 56224 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_419
timestamp 1698431365
transform 1 0 5264 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_420
timestamp 1698431365
transform 1 0 13104 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_421
timestamp 1698431365
transform 1 0 20944 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_422
timestamp 1698431365
transform 1 0 28784 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_423
timestamp 1698431365
transform 1 0 36624 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_424
timestamp 1698431365
transform 1 0 44464 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_425
timestamp 1698431365
transform 1 0 52304 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_426
timestamp 1698431365
transform 1 0 9184 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_427
timestamp 1698431365
transform 1 0 17024 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_428
timestamp 1698431365
transform 1 0 24864 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_429
timestamp 1698431365
transform 1 0 32704 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_430
timestamp 1698431365
transform 1 0 40544 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_431
timestamp 1698431365
transform 1 0 48384 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_432
timestamp 1698431365
transform 1 0 56224 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_433
timestamp 1698431365
transform 1 0 5264 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_434
timestamp 1698431365
transform 1 0 13104 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_435
timestamp 1698431365
transform 1 0 20944 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_436
timestamp 1698431365
transform 1 0 28784 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_437
timestamp 1698431365
transform 1 0 36624 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_438
timestamp 1698431365
transform 1 0 44464 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_439
timestamp 1698431365
transform 1 0 52304 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_440
timestamp 1698431365
transform 1 0 9184 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_441
timestamp 1698431365
transform 1 0 17024 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_442
timestamp 1698431365
transform 1 0 24864 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_443
timestamp 1698431365
transform 1 0 32704 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_444
timestamp 1698431365
transform 1 0 40544 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_445
timestamp 1698431365
transform 1 0 48384 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_446
timestamp 1698431365
transform 1 0 56224 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_447
timestamp 1698431365
transform 1 0 5264 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_448
timestamp 1698431365
transform 1 0 13104 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_449
timestamp 1698431365
transform 1 0 20944 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_450
timestamp 1698431365
transform 1 0 28784 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_451
timestamp 1698431365
transform 1 0 36624 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_452
timestamp 1698431365
transform 1 0 44464 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_453
timestamp 1698431365
transform 1 0 52304 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_454
timestamp 1698431365
transform 1 0 9184 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_455
timestamp 1698431365
transform 1 0 17024 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_456
timestamp 1698431365
transform 1 0 24864 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_457
timestamp 1698431365
transform 1 0 32704 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_458
timestamp 1698431365
transform 1 0 40544 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_459
timestamp 1698431365
transform 1 0 48384 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_460
timestamp 1698431365
transform 1 0 56224 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_461
timestamp 1698431365
transform 1 0 5264 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_462
timestamp 1698431365
transform 1 0 13104 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_463
timestamp 1698431365
transform 1 0 20944 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_464
timestamp 1698431365
transform 1 0 28784 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_465
timestamp 1698431365
transform 1 0 36624 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_466
timestamp 1698431365
transform 1 0 44464 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_467
timestamp 1698431365
transform 1 0 52304 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_468
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_469
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_470
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_471
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_472
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_473
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_474
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_475
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_476
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_477
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_478
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_479
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_480
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_481
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -90 310 1098
<< labels >>
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 in[0]
port 1 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 in[10]
port 2 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 in[11]
port 3 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 in[12]
port 4 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 in[13]
port 5 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 in[14]
port 6 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 in[15]
port 7 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 in[16]
port 8 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 in[17]
port 9 nsew signal input
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 in[1]
port 10 nsew signal input
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 in[2]
port 11 nsew signal input
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 in[3]
port 12 nsew signal input
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 in[4]
port 13 nsew signal input
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 in[5]
port 14 nsew signal input
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 in[6]
port 15 nsew signal input
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 in[7]
port 16 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 in[8]
port 17 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 in[9]
port 18 nsew signal input
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 out[0]
port 19 nsew signal tristate
flabel metal3 s 0 53760 800 53872 0 FreeSans 448 0 0 0 out[10]
port 20 nsew signal tristate
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 out[11]
port 21 nsew signal tristate
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 out[1]
port 22 nsew signal tristate
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 out[2]
port 23 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 out[3]
port 24 nsew signal tristate
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 out[4]
port 25 nsew signal tristate
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 out[5]
port 26 nsew signal tristate
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 out[6]
port 27 nsew signal tristate
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 out[7]
port 28 nsew signal tristate
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 out[8]
port 29 nsew signal tristate
flabel metal3 s 59200 53760 60000 53872 0 FreeSans 448 0 0 0 out[9]
port 30 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 rst_n
port 31 nsew signal input
flabel metal4 s 4448 3972 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 35168 3972 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 19808 3972 20128 56508 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
flabel metal4 s 50528 3972 50848 56508 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
rlabel metal1 29960 55440 29960 55440 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 27160 35504 27160 35504 0 _000_
rlabel metal2 31416 32648 31416 32648 0 _001_
rlabel metal2 32312 34328 32312 34328 0 _002_
rlabel metal2 25592 33208 25592 33208 0 _003_
rlabel metal2 26040 32256 26040 32256 0 _004_
rlabel metal2 23968 30632 23968 30632 0 _005_
rlabel metal2 23464 35000 23464 35000 0 _006_
rlabel metal3 19992 36568 19992 36568 0 _007_
rlabel metal2 17304 37856 17304 37856 0 _008_
rlabel metal2 18760 35728 18760 35728 0 _009_
rlabel metal2 17976 39928 17976 39928 0 _010_
rlabel metal3 18816 36120 18816 36120 0 _011_
rlabel metal3 12208 32536 12208 32536 0 _012_
rlabel metal2 20496 29960 20496 29960 0 _013_
rlabel metal2 18200 32200 18200 32200 0 _014_
rlabel metal2 16408 33152 16408 33152 0 _015_
rlabel metal2 17752 30352 17752 30352 0 _016_
rlabel metal3 36736 28616 36736 28616 0 _017_
rlabel metal2 27832 28224 27832 28224 0 _018_
rlabel metal2 40264 28784 40264 28784 0 _019_
rlabel metal2 45248 16632 45248 16632 0 _020_
rlabel metal2 53032 16688 53032 16688 0 _021_
rlabel metal2 39088 30632 39088 30632 0 _022_
rlabel metal2 46984 15120 46984 15120 0 _023_
rlabel metal2 54264 16688 54264 16688 0 _024_
rlabel metal3 52640 17864 52640 17864 0 _025_
rlabel metal2 53648 15848 53648 15848 0 _026_
rlabel metal2 47992 19152 47992 19152 0 _027_
rlabel metal2 49336 15680 49336 15680 0 _028_
rlabel metal2 45080 30632 45080 30632 0 _029_
rlabel metal2 48216 29176 48216 29176 0 _030_
rlabel metal2 47880 26992 47880 26992 0 _031_
rlabel metal2 40880 30632 40880 30632 0 _032_
rlabel metal3 49056 31752 49056 31752 0 _033_
rlabel metal2 47432 25536 47432 25536 0 _034_
rlabel metal3 49168 19880 49168 19880 0 _035_
rlabel metal2 34888 24976 34888 24976 0 _036_
rlabel metal2 29792 24696 29792 24696 0 _037_
rlabel metal3 30996 26712 30996 26712 0 _038_
rlabel metal2 26712 35224 26712 35224 0 _039_
rlabel metal2 29176 24752 29176 24752 0 _040_
rlabel metal2 26264 21504 26264 21504 0 _041_
rlabel metal2 30072 23128 30072 23128 0 _042_
rlabel metal2 29512 25088 29512 25088 0 _043_
rlabel metal2 32368 25704 32368 25704 0 _044_
rlabel metal2 37576 26600 37576 26600 0 _045_
rlabel via1 28392 25709 28392 25709 0 _046_
rlabel metal2 28336 26600 28336 26600 0 _047_
rlabel metal3 42056 20888 42056 20888 0 _048_
rlabel metal2 44072 21112 44072 21112 0 _049_
rlabel metal2 46200 16184 46200 16184 0 _050_
rlabel metal2 43736 20552 43736 20552 0 _051_
rlabel metal3 42448 21000 42448 21000 0 _052_
rlabel metal2 29400 22680 29400 22680 0 _053_
rlabel metal2 26488 27496 26488 27496 0 _054_
rlabel metal2 24584 30800 24584 30800 0 _055_
rlabel metal2 21280 28728 21280 28728 0 _056_
rlabel metal2 15064 30240 15064 30240 0 _057_
rlabel metal2 24248 29232 24248 29232 0 _058_
rlabel metal3 32424 30632 32424 30632 0 _059_
rlabel metal2 41272 29176 41272 29176 0 _060_
rlabel metal2 39816 29792 39816 29792 0 _061_
rlabel metal3 42952 42728 42952 42728 0 _062_
rlabel metal3 53032 32648 53032 32648 0 _063_
rlabel metal2 54152 45080 54152 45080 0 _064_
rlabel metal2 44072 42392 44072 42392 0 _065_
rlabel metal2 50680 40600 50680 40600 0 _066_
rlabel metal2 42392 42224 42392 42224 0 _067_
rlabel metal2 42616 44632 42616 44632 0 _068_
rlabel metal2 52696 31024 52696 31024 0 _069_
rlabel metal2 53032 45080 53032 45080 0 _070_
rlabel metal2 42168 44688 42168 44688 0 _071_
rlabel metal2 41888 41944 41888 41944 0 _072_
rlabel metal3 38136 41496 38136 41496 0 _073_
rlabel metal2 25928 29904 25928 29904 0 _074_
rlabel metal2 26712 26712 26712 26712 0 _075_
rlabel metal3 26936 26488 26936 26488 0 _076_
rlabel metal2 38584 16072 38584 16072 0 _077_
rlabel metal2 28392 17808 28392 17808 0 _078_
rlabel metal2 36344 14728 36344 14728 0 _079_
rlabel metal2 27944 26096 27944 26096 0 _080_
rlabel metal2 32872 22456 32872 22456 0 _081_
rlabel metal2 38920 22848 38920 22848 0 _082_
rlabel metal3 36960 25816 36960 25816 0 _083_
rlabel metal2 31416 25312 31416 25312 0 _084_
rlabel metal2 37352 39256 37352 39256 0 _085_
rlabel metal2 32760 39480 32760 39480 0 _086_
rlabel metal2 31808 25704 31808 25704 0 _087_
rlabel metal2 31416 26208 31416 26208 0 _088_
rlabel metal2 25144 31808 25144 31808 0 _089_
rlabel metal2 27160 26376 27160 26376 0 _090_
rlabel metal3 20328 28616 20328 28616 0 _091_
rlabel metal2 32200 16688 32200 16688 0 _092_
rlabel metal2 31304 24192 31304 24192 0 _093_
rlabel metal2 27160 18256 27160 18256 0 _094_
rlabel metal2 31640 12656 31640 12656 0 _095_
rlabel metal2 31080 12152 31080 12152 0 _096_
rlabel metal2 26936 21924 26936 21924 0 _097_
rlabel metal2 22792 24136 22792 24136 0 _098_
rlabel metal3 25592 23800 25592 23800 0 _099_
rlabel metal2 26152 23016 26152 23016 0 _100_
rlabel metal2 26544 23912 26544 23912 0 _101_
rlabel metal2 26376 24920 26376 24920 0 _102_
rlabel metal2 34440 23352 34440 23352 0 _103_
rlabel metal2 37632 23912 37632 23912 0 _104_
rlabel metal2 36008 25928 36008 25928 0 _105_
rlabel metal2 37464 25200 37464 25200 0 _106_
rlabel metal2 38696 25872 38696 25872 0 _107_
rlabel metal2 23912 22624 23912 22624 0 _108_
rlabel metal2 39144 25032 39144 25032 0 _109_
rlabel metal2 39256 25368 39256 25368 0 _110_
rlabel metal2 36904 33936 36904 33936 0 _111_
rlabel metal2 37240 33936 37240 33936 0 _112_
rlabel metal2 38864 30968 38864 30968 0 _113_
rlabel metal2 38024 37744 38024 37744 0 _114_
rlabel metal2 37352 28616 37352 28616 0 _115_
rlabel metal2 35672 28392 35672 28392 0 _116_
rlabel metal2 33544 27328 33544 27328 0 _117_
rlabel metal2 34552 28672 34552 28672 0 _118_
rlabel metal2 33320 45864 33320 45864 0 _119_
rlabel metal2 33096 32088 33096 32088 0 _120_
rlabel metal2 23464 27048 23464 27048 0 _121_
rlabel metal3 33656 28728 33656 28728 0 _122_
rlabel metal2 45136 29736 45136 29736 0 _123_
rlabel metal3 52472 30408 52472 30408 0 _124_
rlabel metal2 37912 30296 37912 30296 0 _125_
rlabel metal2 35000 28952 35000 28952 0 _126_
rlabel metal2 35112 28840 35112 28840 0 _127_
rlabel metal2 27160 28000 27160 28000 0 _128_
rlabel metal2 26320 29736 26320 29736 0 _129_
rlabel metal2 19432 27608 19432 27608 0 _130_
rlabel metal2 26824 18816 26824 18816 0 _131_
rlabel metal2 24360 16128 24360 16128 0 _132_
rlabel metal2 28168 24976 28168 24976 0 _133_
rlabel metal2 25592 20776 25592 20776 0 _134_
rlabel metal2 24920 20888 24920 20888 0 _135_
rlabel metal2 25256 23800 25256 23800 0 _136_
rlabel metal2 49672 39368 49672 39368 0 _137_
rlabel metal2 54320 39928 54320 39928 0 _138_
rlabel metal2 49112 40264 49112 40264 0 _139_
rlabel metal2 48664 40208 48664 40208 0 _140_
rlabel metal2 50568 41440 50568 41440 0 _141_
rlabel metal2 53256 31892 53256 31892 0 _142_
rlabel metal2 50008 40376 50008 40376 0 _143_
rlabel metal3 48664 40712 48664 40712 0 _144_
rlabel metal2 47320 36736 47320 36736 0 _145_
rlabel metal2 25816 29456 25816 29456 0 _146_
rlabel metal2 18984 28112 18984 28112 0 _147_
rlabel metal2 14448 30520 14448 30520 0 _148_
rlabel metal2 23968 24472 23968 24472 0 _149_
rlabel metal2 24080 48776 24080 48776 0 _150_
rlabel metal3 27440 43400 27440 43400 0 _151_
rlabel metal2 25592 25032 25592 25032 0 _152_
rlabel metal2 26040 24024 26040 24024 0 _153_
rlabel metal2 25144 22008 25144 22008 0 _154_
rlabel metal3 26376 24472 26376 24472 0 _155_
rlabel metal2 25648 23912 25648 23912 0 _156_
rlabel metal2 37912 23016 37912 23016 0 _157_
rlabel metal2 37352 25368 37352 25368 0 _158_
rlabel metal2 38920 26040 38920 26040 0 _159_
rlabel metal2 38808 26320 38808 26320 0 _160_
rlabel metal2 38920 35616 38920 35616 0 _161_
rlabel metal2 38696 30324 38696 30324 0 _162_
rlabel metal2 37240 28336 37240 28336 0 _163_
rlabel metal2 35448 26936 35448 26936 0 _164_
rlabel metal2 35728 29736 35728 29736 0 _165_
rlabel metal2 34328 32592 34328 32592 0 _166_
rlabel metal2 35448 29960 35448 29960 0 _167_
rlabel metal2 38472 31248 38472 31248 0 _168_
rlabel metal2 36176 29736 36176 29736 0 _169_
rlabel metal2 36904 29008 36904 29008 0 _170_
rlabel metal2 28056 28728 28056 28728 0 _171_
rlabel metal2 15064 28672 15064 28672 0 _172_
rlabel metal2 25480 34216 25480 34216 0 _173_
rlabel metal2 31528 44156 31528 44156 0 _174_
rlabel metal2 33992 45864 33992 45864 0 _175_
rlabel metal2 29792 41496 29792 41496 0 _176_
rlabel metal2 27048 34048 27048 34048 0 _177_
rlabel metal2 27440 30744 27440 30744 0 _178_
rlabel metal2 51800 33936 51800 33936 0 _179_
rlabel metal2 54376 23240 54376 23240 0 _180_
rlabel metal3 52696 31752 52696 31752 0 _181_
rlabel metal2 50456 31892 50456 31892 0 _182_
rlabel metal2 53144 34832 53144 34832 0 _183_
rlabel metal2 53256 30128 53256 30128 0 _184_
rlabel metal2 53872 29960 53872 29960 0 _185_
rlabel metal3 51072 33432 51072 33432 0 _186_
rlabel metal2 49448 30856 49448 30856 0 _187_
rlabel metal2 27048 30744 27048 30744 0 _188_
rlabel metal3 21896 29960 21896 29960 0 _189_
rlabel metal2 24808 39592 24808 39592 0 _190_
rlabel metal3 25816 41944 25816 41944 0 _191_
rlabel metal2 26992 41496 26992 41496 0 _192_
rlabel metal2 25144 35056 25144 35056 0 _193_
rlabel metal2 26600 30968 26600 30968 0 _194_
rlabel metal3 36400 22904 36400 22904 0 _195_
rlabel metal2 36400 27160 36400 27160 0 _196_
rlabel metal2 39592 26712 39592 26712 0 _197_
rlabel metal2 39032 26880 39032 26880 0 _198_
rlabel metal2 40152 36064 40152 36064 0 _199_
rlabel metal2 37352 30016 37352 30016 0 _200_
rlabel metal3 35336 29624 35336 29624 0 _201_
rlabel metal2 35112 24640 35112 24640 0 _202_
rlabel metal2 35224 30072 35224 30072 0 _203_
rlabel metal2 33432 34104 33432 34104 0 _204_
rlabel metal2 35000 30800 35000 30800 0 _205_
rlabel metal2 37352 32200 37352 32200 0 _206_
rlabel metal2 35672 31136 35672 31136 0 _207_
rlabel metal2 34216 30128 34216 30128 0 _208_
rlabel metal3 30520 29848 30520 29848 0 _209_
rlabel metal2 19656 29232 19656 29232 0 _210_
rlabel metal2 53592 22680 53592 22680 0 _211_
rlabel metal3 52528 26712 52528 26712 0 _212_
rlabel metal3 48272 26600 48272 26600 0 _213_
rlabel metal3 44744 25816 44744 25816 0 _214_
rlabel metal3 45248 25704 45248 25704 0 _215_
rlabel metal2 44856 26320 44856 26320 0 _216_
rlabel metal3 28504 26768 28504 26768 0 _217_
rlabel metal2 24696 28112 24696 28112 0 _218_
rlabel metal2 22344 23576 22344 23576 0 _219_
rlabel metal2 22232 26264 22232 26264 0 _220_
rlabel metal3 25144 27720 25144 27720 0 _221_
rlabel metal2 25984 25928 25984 25928 0 _222_
rlabel metal3 25144 28056 25144 28056 0 _223_
rlabel metal2 13160 29512 13160 29512 0 _224_
rlabel metal2 20664 30352 20664 30352 0 _225_
rlabel metal3 24640 29736 24640 29736 0 _226_
rlabel metal2 21784 29064 21784 29064 0 _227_
rlabel metal2 21672 29792 21672 29792 0 _228_
rlabel metal3 20552 30072 20552 30072 0 _229_
rlabel metal2 18536 28504 18536 28504 0 _230_
rlabel metal2 18760 29400 18760 29400 0 _231_
rlabel metal3 15568 30744 15568 30744 0 _232_
rlabel metal2 22344 34440 22344 34440 0 _233_
rlabel metal2 22456 33208 22456 33208 0 _234_
rlabel metal3 21840 33880 21840 33880 0 _235_
rlabel metal2 22232 33152 22232 33152 0 _236_
rlabel metal2 26040 34216 26040 34216 0 _237_
rlabel metal2 20720 35784 20720 35784 0 _238_
rlabel metal2 24136 33712 24136 33712 0 _239_
rlabel metal2 20776 36456 20776 36456 0 _240_
rlabel metal2 13608 32592 13608 32592 0 _241_
rlabel metal2 21448 33320 21448 33320 0 _242_
rlabel metal2 10360 31892 10360 31892 0 _243_
rlabel metal2 30408 7672 30408 7672 0 cm_inst.cc_inst.in\[0\]
rlabel metal3 29904 7672 29904 7672 0 cm_inst.cc_inst.in\[1\]
rlabel metal3 31024 7560 31024 7560 0 cm_inst.cc_inst.in\[2\]
rlabel metal3 21840 7784 21840 7784 0 cm_inst.cc_inst.in\[3\]
rlabel metal2 51576 31808 51576 31808 0 cm_inst.cc_inst.in\[4\]
rlabel metal3 27664 20216 27664 20216 0 cm_inst.cc_inst.in\[5\]
rlabel metal2 51128 14560 51128 14560 0 cm_inst.cc_inst.out_notouch_\[0\]
rlabel metal2 43400 37100 43400 37100 0 cm_inst.cc_inst.out_notouch_\[100\]
rlabel metal2 55048 37464 55048 37464 0 cm_inst.cc_inst.out_notouch_\[101\]
rlabel metal2 41944 37128 41944 37128 0 cm_inst.cc_inst.out_notouch_\[102\]
rlabel metal2 55160 21896 55160 21896 0 cm_inst.cc_inst.out_notouch_\[103\]
rlabel metal2 54824 18312 54824 18312 0 cm_inst.cc_inst.out_notouch_\[104\]
rlabel metal2 40376 42448 40376 42448 0 cm_inst.cc_inst.out_notouch_\[105\]
rlabel metal2 37240 40208 37240 40208 0 cm_inst.cc_inst.out_notouch_\[106\]
rlabel metal3 49504 38696 49504 38696 0 cm_inst.cc_inst.out_notouch_\[107\]
rlabel metal3 43792 38696 43792 38696 0 cm_inst.cc_inst.out_notouch_\[108\]
rlabel metal2 49112 36848 49112 36848 0 cm_inst.cc_inst.out_notouch_\[109\]
rlabel metal2 33656 34664 33656 34664 0 cm_inst.cc_inst.out_notouch_\[10\]
rlabel metal3 43232 36680 43232 36680 0 cm_inst.cc_inst.out_notouch_\[110\]
rlabel metal2 54824 21784 54824 21784 0 cm_inst.cc_inst.out_notouch_\[111\]
rlabel metal2 52752 17752 52752 17752 0 cm_inst.cc_inst.out_notouch_\[112\]
rlabel metal2 36904 42448 36904 42448 0 cm_inst.cc_inst.out_notouch_\[113\]
rlabel metal2 37016 39536 37016 39536 0 cm_inst.cc_inst.out_notouch_\[114\]
rlabel metal3 46648 38808 46648 38808 0 cm_inst.cc_inst.out_notouch_\[115\]
rlabel metal3 41888 37912 41888 37912 0 cm_inst.cc_inst.out_notouch_\[116\]
rlabel metal2 52248 37464 52248 37464 0 cm_inst.cc_inst.out_notouch_\[117\]
rlabel metal2 38920 36680 38920 36680 0 cm_inst.cc_inst.out_notouch_\[118\]
rlabel metal2 52864 20664 52864 20664 0 cm_inst.cc_inst.out_notouch_\[119\]
rlabel metal2 55384 39424 55384 39424 0 cm_inst.cc_inst.out_notouch_\[11\]
rlabel metal2 53368 18200 53368 18200 0 cm_inst.cc_inst.out_notouch_\[120\]
rlabel metal2 39816 43848 39816 43848 0 cm_inst.cc_inst.out_notouch_\[121\]
rlabel metal2 37688 39368 37688 39368 0 cm_inst.cc_inst.out_notouch_\[122\]
rlabel metal2 49336 39200 49336 39200 0 cm_inst.cc_inst.out_notouch_\[123\]
rlabel metal3 40712 38696 40712 38696 0 cm_inst.cc_inst.out_notouch_\[124\]
rlabel metal3 52248 37800 52248 37800 0 cm_inst.cc_inst.out_notouch_\[125\]
rlabel metal2 39760 36008 39760 36008 0 cm_inst.cc_inst.out_notouch_\[126\]
rlabel metal2 53032 21896 53032 21896 0 cm_inst.cc_inst.out_notouch_\[127\]
rlabel metal2 47880 12264 47880 12264 0 cm_inst.cc_inst.out_notouch_\[128\]
rlabel metal2 37016 12376 37016 12376 0 cm_inst.cc_inst.out_notouch_\[129\]
rlabel metal2 34440 32872 34440 32872 0 cm_inst.cc_inst.out_notouch_\[12\]
rlabel metal2 32312 8092 32312 8092 0 cm_inst.cc_inst.out_notouch_\[130\]
rlabel metal2 26152 10640 26152 10640 0 cm_inst.cc_inst.out_notouch_\[131\]
rlabel metal2 27216 46088 27216 46088 0 cm_inst.cc_inst.out_notouch_\[132\]
rlabel metal2 35896 46312 35896 46312 0 cm_inst.cc_inst.out_notouch_\[133\]
rlabel metal2 26040 44156 26040 44156 0 cm_inst.cc_inst.out_notouch_\[134\]
rlabel metal2 24136 25312 24136 25312 0 cm_inst.cc_inst.out_notouch_\[135\]
rlabel metal2 47208 14112 47208 14112 0 cm_inst.cc_inst.out_notouch_\[136\]
rlabel metal2 37464 11536 37464 11536 0 cm_inst.cc_inst.out_notouch_\[137\]
rlabel metal2 32200 10640 32200 10640 0 cm_inst.cc_inst.out_notouch_\[138\]
rlabel metal2 25312 12488 25312 12488 0 cm_inst.cc_inst.out_notouch_\[139\]
rlabel metal2 55048 29400 55048 29400 0 cm_inst.cc_inst.out_notouch_\[13\]
rlabel metal2 25928 47880 25928 47880 0 cm_inst.cc_inst.out_notouch_\[140\]
rlabel metal2 35224 46312 35224 46312 0 cm_inst.cc_inst.out_notouch_\[141\]
rlabel metal2 25312 42840 25312 42840 0 cm_inst.cc_inst.out_notouch_\[142\]
rlabel metal2 23352 25480 23352 25480 0 cm_inst.cc_inst.out_notouch_\[143\]
rlabel metal2 45080 13552 45080 13552 0 cm_inst.cc_inst.out_notouch_\[144\]
rlabel metal2 35336 10864 35336 10864 0 cm_inst.cc_inst.out_notouch_\[145\]
rlabel metal2 30128 12488 30128 12488 0 cm_inst.cc_inst.out_notouch_\[146\]
rlabel metal2 22568 11760 22568 11760 0 cm_inst.cc_inst.out_notouch_\[147\]
rlabel metal2 20608 46648 20608 46648 0 cm_inst.cc_inst.out_notouch_\[148\]
rlabel metal2 31080 46816 31080 46816 0 cm_inst.cc_inst.out_notouch_\[149\]
rlabel metal2 32200 37968 32200 37968 0 cm_inst.cc_inst.out_notouch_\[14\]
rlabel metal3 21896 42840 21896 42840 0 cm_inst.cc_inst.out_notouch_\[150\]
rlabel metal2 21000 25704 21000 25704 0 cm_inst.cc_inst.out_notouch_\[151\]
rlabel metal2 45696 11480 45696 11480 0 cm_inst.cc_inst.out_notouch_\[152\]
rlabel metal2 36792 12152 36792 12152 0 cm_inst.cc_inst.out_notouch_\[153\]
rlabel metal2 30688 11816 30688 11816 0 cm_inst.cc_inst.out_notouch_\[154\]
rlabel metal2 22904 10360 22904 10360 0 cm_inst.cc_inst.out_notouch_\[155\]
rlabel metal2 23128 48440 23128 48440 0 cm_inst.cc_inst.out_notouch_\[156\]
rlabel metal3 32648 45864 32648 45864 0 cm_inst.cc_inst.out_notouch_\[157\]
rlabel metal3 22792 44632 22792 44632 0 cm_inst.cc_inst.out_notouch_\[158\]
rlabel metal2 21392 23912 21392 23912 0 cm_inst.cc_inst.out_notouch_\[159\]
rlabel metal2 47208 26096 47208 26096 0 cm_inst.cc_inst.out_notouch_\[15\]
rlabel metal2 45976 17864 45976 17864 0 cm_inst.cc_inst.out_notouch_\[160\]
rlabel metal2 42560 12824 42560 12824 0 cm_inst.cc_inst.out_notouch_\[161\]
rlabel metal3 36568 15848 36568 15848 0 cm_inst.cc_inst.out_notouch_\[162\]
rlabel metal2 28504 17248 28504 17248 0 cm_inst.cc_inst.out_notouch_\[163\]
rlabel metal3 25088 13832 25088 13832 0 cm_inst.cc_inst.out_notouch_\[164\]
rlabel metal3 33656 43064 33656 43064 0 cm_inst.cc_inst.out_notouch_\[165\]
rlabel metal2 26600 39592 26600 39592 0 cm_inst.cc_inst.out_notouch_\[166\]
rlabel metal2 24136 21308 24136 21308 0 cm_inst.cc_inst.out_notouch_\[167\]
rlabel metal2 45192 20916 45192 20916 0 cm_inst.cc_inst.out_notouch_\[168\]
rlabel metal2 42112 14840 42112 14840 0 cm_inst.cc_inst.out_notouch_\[169\]
rlabel metal2 48328 13608 48328 13608 0 cm_inst.cc_inst.out_notouch_\[16\]
rlabel metal2 35336 17472 35336 17472 0 cm_inst.cc_inst.out_notouch_\[170\]
rlabel metal2 28952 14952 28952 14952 0 cm_inst.cc_inst.out_notouch_\[171\]
rlabel metal2 20216 15120 20216 15120 0 cm_inst.cc_inst.out_notouch_\[172\]
rlabel metal2 35560 48384 35560 48384 0 cm_inst.cc_inst.out_notouch_\[173\]
rlabel metal2 23688 39424 23688 39424 0 cm_inst.cc_inst.out_notouch_\[174\]
rlabel metal1 23072 22008 23072 22008 0 cm_inst.cc_inst.out_notouch_\[175\]
rlabel metal3 42168 21672 42168 21672 0 cm_inst.cc_inst.out_notouch_\[176\]
rlabel metal2 39816 15008 39816 15008 0 cm_inst.cc_inst.out_notouch_\[177\]
rlabel metal2 33208 18256 33208 18256 0 cm_inst.cc_inst.out_notouch_\[178\]
rlabel metal2 26488 17584 26488 17584 0 cm_inst.cc_inst.out_notouch_\[179\]
rlabel metal2 48720 45864 48720 45864 0 cm_inst.cc_inst.out_notouch_\[17\]
rlabel metal2 22904 13608 22904 13608 0 cm_inst.cc_inst.out_notouch_\[180\]
rlabel metal2 30520 44408 30520 44408 0 cm_inst.cc_inst.out_notouch_\[181\]
rlabel metal2 23800 39424 23800 39424 0 cm_inst.cc_inst.out_notouch_\[182\]
rlabel metal2 21336 22232 21336 22232 0 cm_inst.cc_inst.out_notouch_\[183\]
rlabel metal2 43680 21672 43680 21672 0 cm_inst.cc_inst.out_notouch_\[184\]
rlabel metal2 40488 14112 40488 14112 0 cm_inst.cc_inst.out_notouch_\[185\]
rlabel metal2 33880 16296 33880 16296 0 cm_inst.cc_inst.out_notouch_\[186\]
rlabel metal2 28056 16128 28056 16128 0 cm_inst.cc_inst.out_notouch_\[187\]
rlabel metal2 23576 14448 23576 14448 0 cm_inst.cc_inst.out_notouch_\[188\]
rlabel metal2 31248 44184 31248 44184 0 cm_inst.cc_inst.out_notouch_\[189\]
rlabel metal2 33096 28168 33096 28168 0 cm_inst.cc_inst.out_notouch_\[18\]
rlabel metal2 24472 39256 24472 39256 0 cm_inst.cc_inst.out_notouch_\[190\]
rlabel metal2 22064 21896 22064 21896 0 cm_inst.cc_inst.out_notouch_\[191\]
rlabel metal2 29232 21784 29232 21784 0 cm_inst.cc_inst.out_notouch_\[192\]
rlabel metal2 33880 39256 33880 39256 0 cm_inst.cc_inst.out_notouch_\[193\]
rlabel metal2 16296 21672 16296 21672 0 cm_inst.cc_inst.out_notouch_\[194\]
rlabel metal2 17752 19264 17752 19264 0 cm_inst.cc_inst.out_notouch_\[195\]
rlabel metal2 25480 21056 25480 21056 0 cm_inst.cc_inst.out_notouch_\[196\]
rlabel metal2 28392 34608 28392 34608 0 cm_inst.cc_inst.out_notouch_\[197\]
rlabel metal2 26488 36176 26488 36176 0 cm_inst.cc_inst.out_notouch_\[198\]
rlabel metal2 26264 25592 26264 25592 0 cm_inst.cc_inst.out_notouch_\[199\]
rlabel metal2 52696 39816 52696 39816 0 cm_inst.cc_inst.out_notouch_\[19\]
rlabel metal1 51128 43176 51128 43176 0 cm_inst.cc_inst.out_notouch_\[1\]
rlabel metal2 29624 21336 29624 21336 0 cm_inst.cc_inst.out_notouch_\[200\]
rlabel metal2 33432 40264 33432 40264 0 cm_inst.cc_inst.out_notouch_\[201\]
rlabel metal2 15736 22232 15736 22232 0 cm_inst.cc_inst.out_notouch_\[202\]
rlabel metal2 18200 19824 18200 19824 0 cm_inst.cc_inst.out_notouch_\[203\]
rlabel metal2 24584 21280 24584 21280 0 cm_inst.cc_inst.out_notouch_\[204\]
rlabel metal2 27832 35224 27832 35224 0 cm_inst.cc_inst.out_notouch_\[205\]
rlabel metal2 25928 36232 25928 36232 0 cm_inst.cc_inst.out_notouch_\[206\]
rlabel metal2 28392 23688 28392 23688 0 cm_inst.cc_inst.out_notouch_\[208\]
rlabel metal2 32144 24024 32144 24024 0 cm_inst.cc_inst.out_notouch_\[209\]
rlabel metal2 35784 27832 35784 27832 0 cm_inst.cc_inst.out_notouch_\[20\]
rlabel metal2 52920 29960 52920 29960 0 cm_inst.cc_inst.out_notouch_\[21\]
rlabel metal2 35056 25704 35056 25704 0 cm_inst.cc_inst.out_notouch_\[22\]
rlabel metal2 45080 24808 45080 24808 0 cm_inst.cc_inst.out_notouch_\[23\]
rlabel metal2 49000 14784 49000 14784 0 cm_inst.cc_inst.out_notouch_\[24\]
rlabel metal2 48104 44968 48104 44968 0 cm_inst.cc_inst.out_notouch_\[25\]
rlabel metal3 33432 26712 33432 26712 0 cm_inst.cc_inst.out_notouch_\[26\]
rlabel metal2 53480 39424 53480 39424 0 cm_inst.cc_inst.out_notouch_\[27\]
rlabel metal2 35392 26712 35392 26712 0 cm_inst.cc_inst.out_notouch_\[28\]
rlabel metal2 53592 29400 53592 29400 0 cm_inst.cc_inst.out_notouch_\[29\]
rlabel metal2 34328 33880 34328 33880 0 cm_inst.cc_inst.out_notouch_\[2\]
rlabel metal2 34552 23912 34552 23912 0 cm_inst.cc_inst.out_notouch_\[30\]
rlabel metal2 45752 26320 45752 26320 0 cm_inst.cc_inst.out_notouch_\[31\]
rlabel metal2 50008 21000 50008 21000 0 cm_inst.cc_inst.out_notouch_\[32\]
rlabel metal2 41944 46424 41944 46424 0 cm_inst.cc_inst.out_notouch_\[33\]
rlabel metal2 47544 29120 47544 29120 0 cm_inst.cc_inst.out_notouch_\[34\]
rlabel metal2 55496 44352 55496 44352 0 cm_inst.cc_inst.out_notouch_\[35\]
rlabel metal2 47880 31752 47880 31752 0 cm_inst.cc_inst.out_notouch_\[36\]
rlabel metal2 55832 36008 55832 36008 0 cm_inst.cc_inst.out_notouch_\[37\]
rlabel metal2 42224 32648 42224 32648 0 cm_inst.cc_inst.out_notouch_\[38\]
rlabel metal2 55720 24136 55720 24136 0 cm_inst.cc_inst.out_notouch_\[39\]
rlabel metal2 55720 39536 55720 39536 0 cm_inst.cc_inst.out_notouch_\[3\]
rlabel metal2 49112 18256 49112 18256 0 cm_inst.cc_inst.out_notouch_\[40\]
rlabel metal2 41272 47768 41272 47768 0 cm_inst.cc_inst.out_notouch_\[41\]
rlabel metal2 46872 31192 46872 31192 0 cm_inst.cc_inst.out_notouch_\[42\]
rlabel metal3 54264 44856 54264 44856 0 cm_inst.cc_inst.out_notouch_\[43\]
rlabel metal2 47208 31080 47208 31080 0 cm_inst.cc_inst.out_notouch_\[44\]
rlabel metal2 55048 35168 55048 35168 0 cm_inst.cc_inst.out_notouch_\[45\]
rlabel metal2 41720 32368 41720 32368 0 cm_inst.cc_inst.out_notouch_\[46\]
rlabel metal2 55048 23072 55048 23072 0 cm_inst.cc_inst.out_notouch_\[47\]
rlabel metal2 47208 20244 47208 20244 0 cm_inst.cc_inst.out_notouch_\[48\]
rlabel metal2 38696 45976 38696 45976 0 cm_inst.cc_inst.out_notouch_\[49\]
rlabel metal2 35560 34272 35560 34272 0 cm_inst.cc_inst.out_notouch_\[4\]
rlabel metal2 44744 30352 44744 30352 0 cm_inst.cc_inst.out_notouch_\[50\]
rlabel metal3 52304 44744 52304 44744 0 cm_inst.cc_inst.out_notouch_\[51\]
rlabel metal2 45080 32368 45080 32368 0 cm_inst.cc_inst.out_notouch_\[52\]
rlabel metal2 52248 35784 52248 35784 0 cm_inst.cc_inst.out_notouch_\[53\]
rlabel metal2 39312 32648 39312 32648 0 cm_inst.cc_inst.out_notouch_\[54\]
rlabel metal2 52920 24136 52920 24136 0 cm_inst.cc_inst.out_notouch_\[55\]
rlabel metal2 47656 19096 47656 19096 0 cm_inst.cc_inst.out_notouch_\[56\]
rlabel metal2 39592 46424 39592 46424 0 cm_inst.cc_inst.out_notouch_\[57\]
rlabel metal3 44912 29848 44912 29848 0 cm_inst.cc_inst.out_notouch_\[58\]
rlabel metal3 52640 43960 52640 43960 0 cm_inst.cc_inst.out_notouch_\[59\]
rlabel metal2 55664 29960 55664 29960 0 cm_inst.cc_inst.out_notouch_\[5\]
rlabel metal2 45752 31892 45752 31892 0 cm_inst.cc_inst.out_notouch_\[60\]
rlabel metal2 53592 35168 53592 35168 0 cm_inst.cc_inst.out_notouch_\[61\]
rlabel metal2 40152 32256 40152 32256 0 cm_inst.cc_inst.out_notouch_\[62\]
rlabel metal2 53592 24080 53592 24080 0 cm_inst.cc_inst.out_notouch_\[63\]
rlabel metal2 55944 14280 55944 14280 0 cm_inst.cc_inst.out_notouch_\[64\]
rlabel metal2 45920 41944 45920 41944 0 cm_inst.cc_inst.out_notouch_\[65\]
rlabel metal2 40152 25256 40152 25256 0 cm_inst.cc_inst.out_notouch_\[66\]
rlabel metal2 55496 41160 55496 41160 0 cm_inst.cc_inst.out_notouch_\[67\]
rlabel metal2 42280 25200 42280 25200 0 cm_inst.cc_inst.out_notouch_\[68\]
rlabel metal2 56728 31640 56728 31640 0 cm_inst.cc_inst.out_notouch_\[69\]
rlabel metal2 31752 37408 31752 37408 0 cm_inst.cc_inst.out_notouch_\[6\]
rlabel metal2 40824 27048 40824 27048 0 cm_inst.cc_inst.out_notouch_\[70\]
rlabel metal2 55384 25088 55384 25088 0 cm_inst.cc_inst.out_notouch_\[71\]
rlabel metal2 54824 14784 54824 14784 0 cm_inst.cc_inst.out_notouch_\[72\]
rlabel metal2 45248 41944 45248 41944 0 cm_inst.cc_inst.out_notouch_\[73\]
rlabel metal2 39592 25424 39592 25424 0 cm_inst.cc_inst.out_notouch_\[74\]
rlabel metal2 54880 40824 54880 40824 0 cm_inst.cc_inst.out_notouch_\[75\]
rlabel metal2 41720 26096 41720 26096 0 cm_inst.cc_inst.out_notouch_\[76\]
rlabel metal2 55048 31136 55048 31136 0 cm_inst.cc_inst.out_notouch_\[77\]
rlabel metal2 40264 27160 40264 27160 0 cm_inst.cc_inst.out_notouch_\[78\]
rlabel metal2 54824 27328 54824 27328 0 cm_inst.cc_inst.out_notouch_\[79\]
rlabel metal2 47880 25312 47880 25312 0 cm_inst.cc_inst.out_notouch_\[7\]
rlabel metal2 52696 15176 52696 15176 0 cm_inst.cc_inst.out_notouch_\[80\]
rlabel metal2 43064 42616 43064 42616 0 cm_inst.cc_inst.out_notouch_\[81\]
rlabel metal2 36904 24808 36904 24808 0 cm_inst.cc_inst.out_notouch_\[82\]
rlabel metal2 52696 41440 52696 41440 0 cm_inst.cc_inst.out_notouch_\[83\]
rlabel metal2 36624 23800 36624 23800 0 cm_inst.cc_inst.out_notouch_\[84\]
rlabel metal2 52920 32200 52920 32200 0 cm_inst.cc_inst.out_notouch_\[85\]
rlabel metal2 36344 23240 36344 23240 0 cm_inst.cc_inst.out_notouch_\[86\]
rlabel metal2 52696 26768 52696 26768 0 cm_inst.cc_inst.out_notouch_\[87\]
rlabel metal2 53424 15736 53424 15736 0 cm_inst.cc_inst.out_notouch_\[88\]
rlabel metal2 43792 41944 43792 41944 0 cm_inst.cc_inst.out_notouch_\[89\]
rlabel metal2 50456 14112 50456 14112 0 cm_inst.cc_inst.out_notouch_\[8\]
rlabel metal2 36232 23184 36232 23184 0 cm_inst.cc_inst.out_notouch_\[90\]
rlabel metal2 53368 41720 53368 41720 0 cm_inst.cc_inst.out_notouch_\[91\]
rlabel metal2 38136 21420 38136 21420 0 cm_inst.cc_inst.out_notouch_\[92\]
rlabel metal2 53592 31696 53592 31696 0 cm_inst.cc_inst.out_notouch_\[93\]
rlabel metal2 37352 21560 37352 21560 0 cm_inst.cc_inst.out_notouch_\[94\]
rlabel metal2 53368 26264 53368 26264 0 cm_inst.cc_inst.out_notouch_\[95\]
rlabel metal2 55720 17360 55720 17360 0 cm_inst.cc_inst.out_notouch_\[96\]
rlabel metal2 42056 43792 42056 43792 0 cm_inst.cc_inst.out_notouch_\[97\]
rlabel metal2 39816 39088 39816 39088 0 cm_inst.cc_inst.out_notouch_\[98\]
rlabel metal2 51464 39088 51464 39088 0 cm_inst.cc_inst.out_notouch_\[99\]
rlabel metal2 50904 46256 50904 46256 0 cm_inst.cc_inst.out_notouch_\[9\]
rlabel metal3 40824 35784 40824 35784 0 cm_inst.page\[0\]
rlabel metal2 49392 32648 49392 32648 0 cm_inst.page\[1\]
rlabel metal3 34496 34776 34496 34776 0 cm_inst.page\[2\]
rlabel metal2 36456 30688 36456 30688 0 cm_inst.page\[3\]
rlabel metal2 28616 31136 28616 31136 0 cm_inst.page\[4\]
rlabel metal2 26040 31360 26040 31360 0 cm_inst.page\[5\]
rlabel metal2 8344 30800 8344 30800 0 in[0]
rlabel metal3 854 34328 854 34328 0 in[1]
rlabel metal3 4158 32312 4158 32312 0 in[2]
rlabel metal2 21952 37688 21952 37688 0 in[3]
rlabel metal3 7938 33656 7938 33656 0 in[4]
rlabel metal3 2478 36344 2478 36344 0 in[5]
rlabel metal2 18648 35784 18648 35784 0 in[6]
rlabel metal3 14168 35056 14168 35056 0 in[7]
rlabel metal3 4578 30296 4578 30296 0 out[0]
rlabel metal3 2310 53816 2310 53816 0 out[10]
rlabel metal3 2534 7448 2534 7448 0 out[11]
rlabel metal2 15512 29344 15512 29344 0 out[1]
rlabel metal3 8862 28952 8862 28952 0 out[2]
rlabel metal2 15064 27160 15064 27160 0 out[3]
rlabel metal3 3766 27608 3766 27608 0 out[4]
rlabel metal2 13944 28840 13944 28840 0 out[5]
rlabel metal3 7574 31640 7574 31640 0 out[6]
rlabel metal3 11088 30072 11088 30072 0 out[7]
rlabel metal3 2310 6776 2310 6776 0 out[8]
rlabel metal2 56112 54152 56112 54152 0 out[9]
rlabel metal2 12936 30912 12936 30912 0 ro_inst.counter\[0\]
rlabel metal2 4984 23520 4984 23520 0 ro_inst.counter\[10\]
rlabel metal2 4984 25312 4984 25312 0 ro_inst.counter\[11\]
rlabel metal3 3864 26824 3864 26824 0 ro_inst.counter\[12\]
rlabel metal3 5544 28616 5544 28616 0 ro_inst.counter\[13\]
rlabel metal2 3248 27944 3248 27944 0 ro_inst.counter\[14\]
rlabel metal2 5768 29120 5768 29120 0 ro_inst.counter\[15\]
rlabel metal2 8792 31360 8792 31360 0 ro_inst.counter\[16\]
rlabel metal2 3752 30352 3752 30352 0 ro_inst.counter\[17\]
rlabel metal3 4760 32536 4760 32536 0 ro_inst.counter\[18\]
rlabel metal2 3752 34272 3752 34272 0 ro_inst.counter\[19\]
rlabel metal2 14728 28280 14728 28280 0 ro_inst.counter\[1\]
rlabel metal2 6328 35784 6328 35784 0 ro_inst.counter\[20\]
rlabel metal2 6216 37184 6216 37184 0 ro_inst.counter\[21\]
rlabel metal2 1960 37296 1960 37296 0 ro_inst.counter\[22\]
rlabel metal3 5376 38696 5376 38696 0 ro_inst.counter\[23\]
rlabel metal2 5320 40096 5320 40096 0 ro_inst.counter\[24\]
rlabel metal2 6216 39200 6216 39200 0 ro_inst.counter\[25\]
rlabel metal2 6328 41216 6328 41216 0 ro_inst.counter\[26\]
rlabel metal2 8008 40320 8008 40320 0 ro_inst.counter\[27\]
rlabel metal2 9800 42280 9800 42280 0 ro_inst.counter\[28\]
rlabel metal2 12152 41440 12152 41440 0 ro_inst.counter\[29\]
rlabel metal2 12936 28896 12936 28896 0 ro_inst.counter\[2\]
rlabel metal2 13216 39816 13216 39816 0 ro_inst.counter\[30\]
rlabel metal3 13216 38696 13216 38696 0 ro_inst.counter\[31\]
rlabel metal2 13664 37800 13664 37800 0 ro_inst.counter\[32\]
rlabel metal3 13216 36568 13216 36568 0 ro_inst.counter\[33\]
rlabel metal2 14840 31892 14840 31892 0 ro_inst.counter\[34\]
rlabel metal3 15120 26488 15120 26488 0 ro_inst.counter\[3\]
rlabel metal2 11480 26264 11480 26264 0 ro_inst.counter\[4\]
rlabel metal2 12824 25648 12824 25648 0 ro_inst.counter\[5\]
rlabel metal2 6216 25256 6216 25256 0 ro_inst.counter\[6\]
rlabel metal2 5880 24584 5880 24584 0 ro_inst.counter\[7\]
rlabel metal3 5264 24696 5264 24696 0 ro_inst.counter\[8\]
rlabel metal2 2296 24136 2296 24136 0 ro_inst.counter\[9\]
rlabel metal2 11592 28168 11592 28168 0 ro_inst.counter_n\[0\]
rlabel metal2 1848 25032 1848 25032 0 ro_inst.counter_n\[10\]
rlabel metal2 2352 24696 2352 24696 0 ro_inst.counter_n\[11\]
rlabel metal2 2520 28056 2520 28056 0 ro_inst.counter_n\[12\]
rlabel metal2 6216 28672 6216 28672 0 ro_inst.counter_n\[13\]
rlabel metal2 3192 28952 3192 28952 0 ro_inst.counter_n\[14\]
rlabel metal2 5656 30688 5656 30688 0 ro_inst.counter_n\[15\]
rlabel metal2 6216 31080 6216 31080 0 ro_inst.counter_n\[16\]
rlabel metal3 6664 31752 6664 31752 0 ro_inst.counter_n\[17\]
rlabel metal2 5768 33432 5768 33432 0 ro_inst.counter_n\[18\]
rlabel metal3 4536 35112 4536 35112 0 ro_inst.counter_n\[19\]
rlabel metal2 12320 27720 12320 27720 0 ro_inst.counter_n\[1\]
rlabel metal2 3976 36232 3976 36232 0 ro_inst.counter_n\[20\]
rlabel metal3 4368 36792 4368 36792 0 ro_inst.counter_n\[21\]
rlabel metal2 2744 37184 2744 37184 0 ro_inst.counter_n\[22\]
rlabel metal2 2408 38864 2408 38864 0 ro_inst.counter_n\[23\]
rlabel metal2 2744 40152 2744 40152 0 ro_inst.counter_n\[24\]
rlabel metal2 4088 41104 4088 41104 0 ro_inst.counter_n\[25\]
rlabel metal2 6216 41496 6216 41496 0 ro_inst.counter_n\[26\]
rlabel metal3 7112 40488 7112 40488 0 ro_inst.counter_n\[27\]
rlabel metal2 8120 42392 8120 42392 0 ro_inst.counter_n\[28\]
rlabel metal2 9576 41160 9576 41160 0 ro_inst.counter_n\[29\]
rlabel metal2 13496 26768 13496 26768 0 ro_inst.counter_n\[2\]
rlabel metal2 10360 39704 10360 39704 0 ro_inst.counter_n\[30\]
rlabel metal2 10248 38864 10248 38864 0 ro_inst.counter_n\[31\]
rlabel metal2 10808 37688 10808 37688 0 ro_inst.counter_n\[32\]
rlabel metal2 11368 36120 11368 36120 0 ro_inst.counter_n\[33\]
rlabel metal3 12712 35112 12712 35112 0 ro_inst.counter_n\[34\]
rlabel metal2 12936 26320 12936 26320 0 ro_inst.counter_n\[3\]
rlabel metal3 10528 25368 10528 25368 0 ro_inst.counter_n\[4\]
rlabel metal3 10584 24696 10584 24696 0 ro_inst.counter_n\[5\]
rlabel metal2 8848 24696 8848 24696 0 ro_inst.counter_n\[6\]
rlabel metal2 8120 24528 8120 24528 0 ro_inst.counter_n\[7\]
rlabel metal2 5768 25368 5768 25368 0 ro_inst.counter_n\[8\]
rlabel metal2 4872 23632 4872 23632 0 ro_inst.counter_n\[9\]
rlabel metal2 14056 30576 14056 30576 0 ro_inst.enable
rlabel metal2 12264 31892 12264 31892 0 ro_inst.ring\[0\]
rlabel metal2 14056 33152 14056 33152 0 ro_inst.ring\[1\]
rlabel metal2 11704 30072 11704 30072 0 ro_inst.ring\[2\]
rlabel metal2 10472 30744 10472 30744 0 ro_inst.running
rlabel metal2 11648 30408 11648 30408 0 ro_inst.saved_signal
rlabel metal3 11368 30520 11368 30520 0 ro_inst.signal
rlabel metal2 9912 31080 9912 31080 0 ro_inst.slow_clk_n
rlabel metal3 21672 28728 21672 28728 0 ro_sel\[0\]
rlabel via2 19096 31640 19096 31640 0 ro_sel\[1\]
rlabel metal2 18424 32648 18424 32648 0 ro_sel\[2\]
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
