`default_nettype none

(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__addf_1(input A, B, CI, output CO, S); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__addf_2(input A, B, CI, output CO, S); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__addf_4(input A, B, CI, output CO, S); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__addh_1(input A, B, output CO, S); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__addh_2(input A, B, output CO, S); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__addh_4(input A, B, output CO, S); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__and2_1(input A1, A2, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__and2_2(input A1, A2, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__and2_4(input A1, A2, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__and3_1(input A1, A2, A3, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__and3_2(input A1, A2, A3, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__and3_4(input A1, A2, A3, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__and4_1(input A1, A2, A3, A4, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__and4_2(input A1, A2, A3, A4, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__and4_4(input A1, A2, A3, A4, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__antenna(input I); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi21_1(input A1, A2, B, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi21_2(input A1, A2, B, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi21_4(input A1, A2, B, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi22_1(input A1, A2, B1, B2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi22_2(input A1, A2, B1, B2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi22_4(input A1, A2, B1, B2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi211_1(input A1, A2, B, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi211_2(input A1, A2, B, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi211_4(input A1, A2, B, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi221_1(input A1, A2, B1, B2, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi221_2(input A1, A2, B1, B2, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi221_4(input A1, A2, B1, B2, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi222_1(input A1, A2, B1, B2, C1, C2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi222_2(input A1, A2, B1, B2, C1, C2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__aoi222_4(input A1, A2, B1, B2, C1, C2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__buf_1(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__buf_2(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__buf_3(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__buf_4(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__buf_8(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__buf_12(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__buf_16(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__buf_20(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__bufz_1(input EN, I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__bufz_2(input EN, I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__bufz_3(input EN, I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__bufz_4(input EN, I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__bufz_8(input EN, I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__bufz_12(input EN, I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__bufz_16(input EN, I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkbuf_1(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkbuf_2(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkbuf_3(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkbuf_4(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkbuf_8(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkbuf_12(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkbuf_16(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkbuf_20(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkinv_1(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkinv_2(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkinv_3(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkinv_4(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkinv_8(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkinv_12(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkinv_16(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__clkinv_20(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnq_1(input CLKN, D, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnq_2(input CLKN, D, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnq_4(input CLKN, D, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1(input CLKN, D, RN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2(input CLKN, D, RN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4(input CLKN, D, RN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1(input CLKN, D, RN, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2(input CLKN, D, RN, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4(input CLKN, D, RN, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1(input CLKN, D, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2(input CLKN, D, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4(input CLKN, D, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffq_1(input CLK, D, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffq_2(input CLK, D, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffq_4(input CLK, D, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffrnq_1(input CLK, D, RN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffrnq_2(input CLK, D, RN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffrnq_4(input CLK, D, RN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1(input CLK, D, RN, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2(input CLK, D, RN, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4(input CLK, D, RN, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffsnq_1(input CLK, D, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffsnq_2(input CLK, D, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dffsnq_4(input CLK, D, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlya_1(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlya_2(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlya_4(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlyb_1(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlyb_2(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlyb_4(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlyc_1(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlyc_2(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlyc_4(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlyd_1(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlyd_2(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__dlyd_4(input I, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__endcap(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fill_1(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fill_2(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fill_4(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fill_8(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fill_16(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fill_32(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fill_64(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fillcap_4(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fillcap_8(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fillcap_16(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fillcap_32(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__fillcap_64(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__filltie(); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__hold(inout Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__icgtn_1(input CLKN, E, TE, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__icgtn_2(input CLKN, E, TE, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__icgtn_4(input CLKN, E, TE, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__icgtp_1(input CLK, E, TE, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__icgtp_2(input CLK, E, TE, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__icgtp_4(input CLK, E, TE, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__inv_1(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__inv_2(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__inv_3(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__inv_4(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__inv_8(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__inv_12(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__inv_16(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__inv_20(input I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__invz_1(input EN, I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__invz_2(input EN, I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__invz_3(input EN, I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__invz_4(input EN, I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__invz_8(input EN, I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__invz_12(input EN, I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__invz_16(input EN, I, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latq_1(input D, E, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latq_2(input D, E, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latq_4(input D, E, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latrnq_1(input D, E, RN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latrnq_2(input D, E, RN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latrnq_4(input D, E, RN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latrsnq_1(input D, E, RN, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latrsnq_2(input D, E, RN, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latrsnq_4(input D, E, RN, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latsnq_1(input D, E, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latsnq_2(input D, E, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__latsnq_4(input D, E, SETN, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__mux2_1(input I0, I1, S, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__mux2_2(input I0, I1, S, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__mux2_4(input I0, I1, S, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__mux4_1(input I0, I1, I2, I3, S0, S1, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__mux4_2(input I0, I1, I2, I3, S0, S1, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__mux4_4(input I0, I1, I2, I3, S0, S1, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nand2_1(input A1, A2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nand2_2(input A1, A2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nand2_4(input A1, A2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nand3_1(input A1, A2, A3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nand3_2(input A1, A2, A3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nand3_4(input A1, A2, A3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nand4_1(input A1, A2, A3, A4, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nand4_2(input A1, A2, A3, A4, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nand4_4(input A1, A2, A3, A4, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nor2_1(input A1, A2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nor2_2(input A1, A2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nor2_4(input A1, A2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nor3_1(input A1, A2, A3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nor3_2(input A1, A2, A3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nor3_4(input A1, A2, A3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nor4_1(input A1, A2, A3, A4, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nor4_2(input A1, A2, A3, A4, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__nor4_4(input A1, A2, A3, A4, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai21_1(input A1, A2, B, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai21_2(input A1, A2, B, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai21_4(input A1, A2, B, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai22_1(input A1, A2, B1, B2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai22_2(input A1, A2, B1, B2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai22_4(input A1, A2, B1, B2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai31_1(input A1, A2, A3, B, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai31_2(input A1, A2, A3, B, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai31_4(input A1, A2, A3, B, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai32_1(input A1, A2, A3, B1, B2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai32_2(input A1, A2, A3, B1, B2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai32_4(input A1, A2, A3, B1, B2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai33_1(input A1, A2, A3, B1, B2, B3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai33_2(input A1, A2, A3, B1, B2, B3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai33_4(input A1, A2, A3, B1, B2, B3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai211_1(input A1, A2, B, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai211_2(input A1, A2, B, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai211_4(input A1, A2, B, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai221_1(input A1, A2, B1, B2, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai221_2(input A1, A2, B1, B2, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai221_4(input A1, A2, B1, B2, C, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai222_1(input A1, A2, B1, B2, C1, C2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai222_2(input A1, A2, B1, B2, C1, C2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__oai222_4(input A1, A2, B1, B2, C1, C2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__or2_1(input A1, A2, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__or2_2(input A1, A2, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__or2_4(input A1, A2, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__or3_1(input A1, A2, A3, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__or3_2(input A1, A2, A3, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__or3_4(input A1, A2, A3, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__or4_1(input A1, A2, A3, A4, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__or4_2(input A1, A2, A3, A4, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__or4_4(input A1, A2, A3, A4, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffq_1(input CLK, D, SE, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffq_2(input CLK, D, SE, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffq_4(input CLK, D, SE, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1(input CLK, D, RN, SE, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2(input CLK, D, RN, SE, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4(input CLK, D, RN, SE, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1(input CLK, D, RN, SE, SETN, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2(input CLK, D, RN, SE, SETN, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4(input CLK, D, RN, SE, SETN, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1(input CLK, D, SE, SETN, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2(input CLK, D, SE, SETN, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4(input CLK, D, SE, SETN, SI, output Q); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__tieh(output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__tiel(output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xnor2_1(input A1, A2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xnor2_2(input A1, A2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xnor2_4(input A1, A2, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xnor3_1(input A1, A2, A3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xnor3_2(input A1, A2, A3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xnor3_4(input A1, A2, A3, output ZN); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xor2_1(input A1, A2, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xor2_2(input A1, A2, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xor2_4(input A1, A2, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xor3_1(input A1, A2, A3, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xor3_2(input A1, A2, A3, output Z); endmodule
(* blackbox *) module gf180mcu_fd_sc_mcu9t5v0__xor3_4(input A1, A2, A3, output Z); endmodule

