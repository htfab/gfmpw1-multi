* NGSPICE file created from rotfpga2a.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_2 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_4 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_1 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

.subckt rotfpga2a clk in[0] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17]
+ in[18] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] out[0] out[10] out[11]
+ out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] rst_n vdd vss
X_2106_ _1593_ _1570_ _1571_ _1578_ _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2037_ _1525_ _1526_ _1527_ _1528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_37_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3155_ _0609_ _0590_ _0602_ _0782_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__3691__A2 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3086_ _0518_ _0521_ g.g_y\[3\].g_x\[2\].t.r_h _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3752__CLK net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3988_ net42 _3988_/E g.g_y\[1\].g_x\[7\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2939_ g.g_y\[4\].g_x\[7\].t.r_v _0197_ _0580_ g.g_y\[3\].g_x\[7\].t.r_v _0581_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_9_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1996__A2 _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3842_ g.g_y\[5\].g_x\[4\].t.w_si net119 g.g_y\[5\].g_x\[4\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_42_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3911_ net61 _3911_/E g.g_y\[3\].g_x\[6\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3773_ net98 _3773_/E g.g_y\[7\].g_x\[2\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2655_ g.g_y\[5\].g_x\[3\].t.r_h _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2724_ _0377_ _0378_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout127 net132 net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout105 g.g_y\[7\].g_x\[5\].t.out_sc net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout116 net117 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2586_ g.g_y\[4\].g_x\[5\].t.out_sc _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3553__B _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3207_ _0639_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3069_ _0688_ _0703_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3138_ _0762_ _0764_ _0766_ _0768_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_37_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3352__A1 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout106_I net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ _1727_ _1713_ _1719_ _0112_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_3_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2371_ _0026_ _0035_ _0044_ _0046_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_4041_ net32 _4041_/E g.g_y\[0\].g_x\[4\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_19_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3825_ net83 _3825_/E g.g_y\[5\].g_x\[7\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3756_ g.g_y\[7\].g_x\[5\].t.w_si net131 g.g_y\[7\].g_x\[5\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3582__A1 _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2137__A2 _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2707_ _0319_ _0105_ _0108_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_42_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2569_ g.g_y\[4\].g_x\[5\].t.r_d _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2638_ g.bi_l\[36\]\[0\] g.g_y\[4\].g_x\[4\].t.r_h _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_6_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3687_ _0923_ _1248_ _0695_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3640__C _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1871_ _1365_ _1349_ _1350_ _1357_ _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1940_ _1431_ _1434_ g.g_y\[7\].g_x\[6\].t.r_h _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3610_ _0146_ _1181_ _1182_ _1186_ g.g_y\[6\].g_x\[0\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3472_ _1764_ _1766_ _1072_ _1069_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__2498__I _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2423_ _0093_ _0094_ _0095_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3316__A1 _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ _0955_ _0958_ g.g_y\[1\].g_x\[0\].t.r_v _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2285_ _1405_ net106 _1765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3619__A2 _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2354_ g.bi_l\[36\]\[1\] net69 _0029_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4024_ net35 _4024_/E g.g_y\[1\].g_x\[0\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3808_ net89 _3808_/E g.g_y\[6\].g_x\[3\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XTAP_TAPCELL_ROW_50_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3739_ _1127_ _1119_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1802__A1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3836__CLK net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3986__CLK net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2070_ net102 _1445_ _1560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_64_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2972_ _0581_ _0612_ _0613_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1854_ net92 g.bi_l\[54\]\[1\] g.g_y\[6\].g_x\[6\].t.r_d _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1923_ net108 g.bi_l\[63\]\[1\] g.g_y\[7\].g_x\[7\].t.r_d _1418_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2406_ _0075_ _0077_ _0078_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3524_ _1699_ _1685_ _1692_ _1118_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3455_ _1745_ _1057_ _1058_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3386_ g.g_y\[1\].g_x\[5\].t.r_d _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2337_ _1507_ _0010_ _0012_ _0014_ g.g_y\[6\].g_x\[6\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2268_ _1359_ _1746_ _1750_ g.g_y\[7\].g_x\[0\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2199_ g.g_y\[0\].g_x\[1\].t.r_v _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_4007_ net38 _4007_/E g.g_y\[1\].g_x\[3\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_47_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_10_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2267__A1 _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3240_ _0839_ _0857_ _0863_ _0444_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2053_ _1538_ _1543_ g.g_y\[7\].g_x\[4\].t.r_h _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2122_ _1607_ _1609_ _1601_ _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3171_ g.g_y\[1\].g_x\[5\].t.r_h _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_29_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2955_ _0596_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1837_ _1313_ _1315_ _1317_ _1325_ _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1906_ _1393_ _1388_ _1400_ _1376_ _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_3507_ _1090_ _1092_ _1094_ _1468_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2886_ _1565_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_32_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3438_ _1684_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3369_ _0813_ _0816_ g.g_y\[1\].g_x\[6\].t.r_h _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_67_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2972__A2 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput20 net20 out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2671_ _0328_ _0329_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2740_ _0392_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3376__B _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3140__A2 _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3223_ net38 g.bi_l\[11\]\[1\] g.g_y\[1\].g_x\[3\].t.r_d _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2105_ _1569_ _1593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2036_ g.bi_l\[4\]\[0\] g.g_y\[0\].g_x\[4\].t.r_v _1527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_37_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3154_ _0609_ _0603_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3085_ _0520_ _0505_ _0513_ _0719_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_9_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2938_ g.g_y\[4\].g_x\[7\].t.r_v _0200_ _0204_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3987_ net43 _3987_/E g.g_y\[1\].g_x\[7\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XANTENNA__2651__A1 _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2869_ _0496_ _0505_ _0513_ _0515_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_13_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3772_ g.g_y\[7\].g_x\[2\].t.w_si net127 g.g_y\[7\].g_x\[2\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3841_ g.g_y\[5\].g_x\[4\].t.out_sc _3841_/E g.g_y\[5\].g_x\[4\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XTAP_TAPCELL_ROW_42_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2723_ _0174_ _0182_ _0199_ _0203_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3910_ g.g_y\[3\].g_x\[7\].t.w_na _3910_/E _3910_/RN g.bi_l\[31\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__2936__A2 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2654_ _0283_ _0313_ _0314_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2585_ _0245_ _0247_ _0248_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout106 net107 net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout128 net129 net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout117 net120 net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3206_ _0653_ _0652_ _0660_ _0640_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_10_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3137_ _0732_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2019_ _1491_ _1510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3068_ net48 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3352__A2 _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ _0026_ _0045_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4040_ g.g_y\[0\].g_x\[4\].t.w_si net130 g.g_y\[0\].g_x\[4\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2854__A1 _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3755_ net104 _3755_/E g.g_y\[7\].g_x\[5\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XANTENNA__3582__A2 _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3824_ g.g_y\[6\].g_x\[0\].t.w_na _3824_/E _3824_/RN g.bi_l\[48\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2706_ g.g_y\[5\].g_x\[1\].t.r_h _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3686_ _0878_ _0871_ _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2499_ _0163_ net16 _0165_ _0161_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2568_ _0231_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2637_ _0295_ _0296_ _0297_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2073__A2 _1528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2836__A1 _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1870_ _1348_ _1365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3540_ g.g_y\[0\].g_x\[0\].t.r_v _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_16_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3471_ _1431_ _1434_ g.g_y\[7\].g_x\[6\].t.r_v _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2422_ g.bi_l\[41\]\[0\] g.g_y\[5\].g_x\[1\].t.r_h _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2353_ g.g_y\[4\].g_x\[4\].t.r_d _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2284_ g.g_y\[7\].g_x\[6\].t.r_v _1764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4023_ net35 _4023_/E g.g_y\[1\].g_x\[0\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_59_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2463__B _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1802__A2 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1999_ g.g_y\[6\].g_x\[5\].t.r_d _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3807_ net89 _3807_/E g.g_y\[6\].g_x\[3\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_42_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3738_ _1638_ _1287_ _1290_ _1291_ g.g_y\[0\].g_x\[2\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3555__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3669_ _0616_ _0618_ _0765_ _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1869__A2 _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3307__A2 _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3491__A1 _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3546__A2 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2820__C _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1922_ g.g_y\[7\].g_x\[7\].t.r_h _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_64_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2971_ _0177_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_29_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1853_ g.g_y\[6\].g_x\[6\].t.r_h _1348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3523_ _1693_ _1699_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2336_ _1763_ _0006_ _0008_ _0013_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2405_ _0075_ _1659_ _1662_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3385_ _0993_ _0996_ _0997_ g.g_y\[1\].g_x\[6\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3454_ _0977_ _0941_ _0954_ _0957_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2276__A2 _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2267_ _1747_ _1748_ _1749_ _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2198_ _1680_ _1681_ _1682_ _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4006_ g.g_y\[1\].g_x\[3\].t.w_si net125 g.g_y\[1\].g_x\[3\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3464__A1 _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3170_ _0793_ _0795_ _0796_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2052_ _1539_ _1541_ _1542_ _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2121_ _1569_ _1570_ _1608_ _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__3455__A1 _1745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1905_ _1389_ _1390_ _1391_ _1393_ _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_32_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2954_ g.g_y\[2\].g_x\[0\].t.r_h _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3058__I1 _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2885_ _0491_ _0494_ _0524_ _0531_ g.g_y\[4\].g_x\[2\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1836_ _1311_ _1310_ _1330_ _1300_ _1331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3506_ _1096_ _1103_ g.g_y\[0\].g_x\[4\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2319_ _1790_ _1789_ _1797_ _1798_ _1799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__3826__CLK net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3368_ _0815_ _0797_ _0808_ _0983_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_3299_ _0754_ _0740_ _0746_ _0919_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3437_ _0733_ _0749_ _1042_ _1679_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_67_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3976__CLK net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input11_I in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput21 net21 out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__3221__I1 _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3437__A1 _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout129_I net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2670_ _0091_ _0090_ _0104_ _0107_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_34_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input3_I in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2104_ _1568_ _1579_ _1589_ _1591_ _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3153_ _0607_ _0610_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3222_ g.g_y\[1\].g_x\[3\].t.r_h _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_37_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2035_ g.bi_l\[4\]\[1\] net31 g.g_y\[0\].g_x\[4\].t.r_d _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3084_ _0520_ _0514_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3986_ g.g_y\[1\].g_x\[7\].t.w_si net124 g.g_y\[1\].g_x\[7\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2937_ _0481_ _0577_ _0578_ _0579_ g.g_y\[4\].g_x\[0\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_20_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2868_ _0496_ _0514_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1914__A1 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1819_ g.g_y\[0\].g_x\[6\].t.r_d _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2799_ g.bi_l\[36\]\[0\] g.g_y\[4\].g_x\[4\].t.r_v _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2890__A2 _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Left_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3658__A1 _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_57_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3771_ net99 _3771_/E g.g_y\[7\].g_x\[2\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_54_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3840_ g.g_y\[5\].g_x\[5\].t.w_na _3840_/E _3840_/RN g.bi_l\[45\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XTAP_TAPCELL_ROW_42_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2722_ _0376_ _0192_ _0202_ _0175_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xfanout107 g.g_y\[7\].g_x\[6\].t.out_sc net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout129 net132 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout118 net119 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2653_ _0037_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2584_ g.g_y\[4\].g_x\[5\].t.r_h _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3205_ _0655_ _0532_ _0829_ _0830_ g.g_y\[2\].g_x\[6\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3067_ _0698_ _0700_ _0701_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3136_ _0732_ _0761_ _0767_ g.g_y\[3\].g_x\[1\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2018_ _1490_ _1498_ _1506_ _1508_ _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_18_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3969_ net46 _3969_/E g.g_y\[2\].g_x\[2\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2130__I g.g_y\[6\].g_x\[3\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2854__A2 _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3823_ g.g_y\[6\].g_x\[0\].t.w_dh _3823_/E _3823_/RN g.bi_l\[48\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_19_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3754_ net107 _3754_/E g.g_y\[7\].g_x\[6\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_54_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _0360_ _0362_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2636_ g.bi_l\[34\]\[0\] g.g_y\[4\].g_x\[2\].t.r_h _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3685_ g.g_y\[2\].g_x\[1\].t.r_h _0920_ _0921_ _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2498_ _1440_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2567_ g.g_y\[4\].g_x\[5\].t.r_v _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_65_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3098__A2 _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3119_ _0739_ _0738_ _0750_ _0734_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__3645__I1 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout111_I net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2283_ g.g_y\[6\].g_x\[6\].t.r_d _1763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2352_ _0027_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2421_ net74 g.bi_l\[41\]\[1\] g.g_y\[5\].g_x\[1\].t.r_d _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3470_ _0790_ _0811_ _1070_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_24_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_67_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4022_ g.g_y\[1\].g_x\[0\].t.w_si net114 g.g_y\[1\].g_x\[0\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3806_ g.g_y\[6\].g_x\[3\].t.w_si net116 g.g_y\[6\].g_x\[3\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3599_ g.g_y\[6\].g_x\[1\].t.r_h _0113_ _0114_ _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1998_ _1488_ _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2619_ net77 _0072_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3737_ _1111_ _1113_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3555__A3 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3668_ _0306_ _1230_ _1232_ _1233_ g.g_y\[3\].g_x\[3\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1823__B _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1852_ _1344_ _1346_ _1337_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1921_ _1409_ _1415_ g.g_y\[7\].g_x\[6\].t.r_v _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2970_ _0583_ _0605_ _0611_ _0198_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_21_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__I0 _1528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3522_ _1111_ _1113_ _1115_ _1116_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3453_ _0938_ _0945_ _0956_ _0939_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2404_ _1654_ _1648_ _1653_ _0076_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2266_ _1375_ _1381_ _1398_ _1376_ _1749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2335_ _1564_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3384_ net40 _0883_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2197_ g.bi_l\[9\]\[0\] _1679_ _1682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4005_ net39 _4005_/E g.g_y\[1\].g_x\[3\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_47_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2736__A1 _1773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3161__A1 _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2727__A1 _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2120_ g.bi_l\[59\]\[0\] g.g_y\[7\].g_x\[3\].t.r_v _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4060__CLK net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3662__C _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3152__A1 _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2051_ g.bi_l\[59\]\[0\] g.g_y\[7\].g_x\[3\].t.r_h _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_72_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1835_ _1301_ _1304_ _1305_ _1311_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_60_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1904_ _1374_ _1381_ _1398_ _1395_ _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_2953_ _0592_ _0593_ _0594_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2884_ _0528_ _0530_ _0491_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3505_ _1468_ _1100_ _1102_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3143__A1 _1745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3436_ g.g_y\[2\].g_x\[1\].t.r_v _0752_ _0756_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2318_ g.g_y\[5\].g_x\[6\].t.r_d _1798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2249_ g.g_y\[7\].g_x\[1\].t.r_h _1734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3367_ _0815_ _0809_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3298_ _0754_ _0747_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput22 net22 out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__3437__A2 _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3657__C _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2103_ _1590_ _1568_ _1591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3152_ _0774_ _0779_ _0780_ g.g_y\[2\].g_x\[7\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3221_ _0842_ _0844_ _0838_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3083_ g.g_y\[3\].g_x\[2\].t.r_h _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3428__A2 _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2034_ g.g_y\[0\].g_x\[4\].t.r_v _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3985_ net42 _3985_/E g.g_y\[1\].g_x\[7\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_72_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3600__A2 _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1818_ g.g_y\[0\].g_x\[6\].t.r_h _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2936_ net62 _0274_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_20_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2798_ _0444_ _0446_ _0447_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2867_ net55 _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3667__A2 _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3419_ _0914_ _0908_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3658__A2 _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3816__CLK net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3770_ g.g_y\[7\].g_x\[3\].t.w_na _3770_/E _3770_/RN g.bi_l\[59\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XTAP_TAPCELL_ROW_42_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2652_ _0285_ _0305_ _0312_ _1623_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2721_ _0193_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout108 net109 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout119 net120 net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2583_ _0184_ _0185_ _0246_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3204_ _0785_ _0824_ _0826_ _0432_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3966__CLK net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2017_ _1490_ _1507_ _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3066_ g.g_y\[2\].g_x\[3\].t.r_h _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3135_ _0762_ _0764_ _0766_ _0732_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3968_ g.g_y\[2\].g_x\[3\].t.out_sc _3968_/E g.g_y\[2\].g_x\[3\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2919_ g.g_y\[3\].g_x\[0\].t.r_h _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3899_ net65 _3899_/E g.g_y\[4\].g_x\[0\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_5_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3822_ net85 _3822_/E g.g_y\[6\].g_x\[0\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3753_ net106 _3753_/E g.g_y\[7\].g_x\[6\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2704_ _0125_ _1722_ _0361_ _1707_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3684_ _0444_ _1243_ _1245_ _1246_ g.g_y\[2\].g_x\[4\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2635_ net66 g.bi_l\[34\]\[1\] g.g_y\[4\].g_x\[2\].t.r_d _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2566_ g.g_y\[6\].g_x\[5\].t.r_v _1509_ _0229_ g.g_y\[5\].g_x\[5\].t.r_v _0230_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2497_ _0162_ _0166_ g.g_y\[6\].g_x\[0\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_53_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3049_ g.g_y\[4\].g_x\[3\].t.r_v _0308_ _0311_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_2_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3118_ _1680_ _1681_ _0735_ _0739_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_52_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2387__B _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2297__A1 _1773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout90 net91 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2420_ g.g_y\[5\].g_x\[1\].t.r_h _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_36_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2282_ _1762_ net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2351_ g.g_y\[4\].g_x\[4\].t.r_v _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_19_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4021_ g.g_y\[1\].g_x\[0\].t.out_sc _4021_/E g.g_y\[1\].g_x\[0\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_59_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1997_ g.g_y\[6\].g_x\[5\].t.r_v _1488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3805_ g.g_y\[6\].g_x\[3\].t.out_sc _3805_/E g.g_y\[6\].g_x\[3\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_3736_ _1288_ _1289_ _1583_ _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2549_ _1798_ _1781_ _1791_ _0216_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3598_ _1530_ _1173_ _1175_ _1176_ g.g_y\[6\].g_x\[4\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2618_ _0278_ _0279_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3667_ g.g_y\[4\].g_x\[3\].t.r_v _0305_ _0684_ _0306_ _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_29_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1851_ _1301_ _1304_ _1345_ _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1920_ _1411_ _1412_ _1414_ _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2403_ _1637_ net98 _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2745__A2 _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3521_ _1581_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3383_ _0994_ _0995_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3452_ _0724_ _1053_ _1055_ _1056_ g.g_y\[1\].g_x\[1\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2334_ _1413_ _1768_ _0011_ g.g_y\[6\].g_x\[6\].t.r_d _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2265_ _1393_ _1388_ _1400_ _1395_ _1748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4004_ g.g_y\[1\].g_x\[4\].t.out_sc _4004_/E g.g_y\[1\].g_x\[4\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_2196_ g.bi_l\[9\]\[1\] net36 g.g_y\[1\].g_x\[1\].t.r_d _1681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_63_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2736__A2 _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2984__A2 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3719_ _1274_ _1275_ _1679_ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3161__A2 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ net100 g.bi_l\[59\]\[1\] _1540_ _1541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2952_ g.bi_l\[22\]\[0\] g.g_y\[2\].g_x\[6\].t.r_h _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2415__A1 _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1834_ _1300_ _1312_ _1326_ _1328_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_1903_ net17 g.g_y\[7\].g_x\[0\].t.r_h _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2883_ _0486_ _0477_ _0529_ _0295_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3504_ _1085_ _1077_ _1101_ _1467_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3366_ g.g_y\[1\].g_x\[6\].t.r_h _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3435_ g.g_y\[1\].g_x\[1\].t.r_d _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2317_ _1782_ _1783_ _1784_ _1790_ _1797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2179_ _1600_ _1630_ _1540_ _1666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2248_ _1702_ _1731_ _1732_ _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3297_ _0889_ _0917_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput23 net23 out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_31_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3220_ _0443_ _0446_ _0843_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2033_ g.g_y\[7\].g_x\[4\].t.r_d _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2102_ g.g_y\[0\].g_x\[3\].t.out_sc _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3151_ net51 _0682_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3082_ _0670_ _0672_ _0716_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_11_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2935_ _0543_ _0570_ _0142_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_20_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3984_ g.g_y\[2\].g_x\[0\].t.w_na _3984_/E _3984_/RN g.bi_l\[16\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__2939__A2 _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1817_ _1306_ _1310_ _1311_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2797_ g.bi_l\[20\]\[0\] g.g_y\[2\].g_x\[4\].t.r_v _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2866_ _0509_ _0511_ _0512_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3349_ _0962_ _0966_ g.g_y\[2\].g_x\[0\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3418_ g.g_y\[1\].g_x\[2\].t.r_h _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4050__CLK net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3594__A2 _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2582_ g.bi_l\[38\]\[0\] g.g_y\[4\].g_x\[6\].t.r_h _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2720_ _0195_ _1746_ _0375_ g.g_y\[5\].g_x\[0\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2651_ _0285_ _0308_ _0311_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xfanout109 net26 net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3203_ _0789_ _0787_ _0828_ g.g_y\[2\].g_x\[6\].t.r_d _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_1_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2016_ g.g_y\[6\].g_x\[5\].t.out_sc _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3065_ _0647_ _0648_ _0699_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3134_ _0616_ _0618_ _0765_ _0762_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3898_ g.g_y\[4\].g_x\[1\].t.out_sc _3898_/E g.g_y\[4\].g_x\[1\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_18_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2632__I1 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3967_ net48 _3967_/E g.g_y\[2\].g_x\[3\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2918_ _0546_ _0550_ _0559_ _0561_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_2849_ g.g_y\[3\].g_x\[2\].t.r_d _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3752_ g.g_y\[7\].g_x\[6\].t.w_si net131 g.g_y\[7\].g_x\[6\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3821_ net86 _3821_/E g.g_y\[6\].g_x\[0\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3567__A2 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2565_ g.g_y\[6\].g_x\[5\].t.r_v _1512_ _1515_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2703_ _1725_ _1729_ _1704_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2634_ _0294_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3683_ g.g_y\[3\].g_x\[4\].t.r_v _0463_ _0836_ _0444_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2496_ _0163_ net16 _0165_ _1385_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3117_ _0734_ _0740_ _0746_ _0748_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_TAPCELL_ROW_18_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3255__A1 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3048_ _0485_ _0681_ _0683_ g.g_y\[3\].g_x\[4\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1837__B _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3558__A2 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3806__CLK net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2297__A2 _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3956__CLK net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout91 g.g_y\[6\].g_x\[4\].t.out_sc net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout80 g.g_y\[5\].g_x\[5\].t.out_sc net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3549__A2 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2281_ _1759_ _1761_ g.g_y\[6\].g_x\[7\].t.r_h _1762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2350_ g.g_y\[5\].g_x\[4\].t.r_d _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_19_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4020_ g.g_y\[1\].g_x\[1\].t.w_na _4020_/E _4020_/RN g.bi_l\[9\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_35_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3804_ g.g_y\[6\].g_x\[4\].t.w_na _3804_/E _3804_/RN g.bi_l\[52\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_1996_ _1454_ _1479_ _1486_ g.g_y\[7\].g_x\[5\].t.r_v _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_50_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2212__A2 _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2332__I _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3735_ g.g_y\[0\].g_x\[1\].t.r_h _1119_ _1120_ _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2548_ _1798_ _1792_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3597_ _0019_ _0021_ _0022_ _1530_ _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2617_ _0025_ _0034_ _0048_ _0051_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_7_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3666_ _0717_ _1231_ _0715_ _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2279__A2 _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2479_ _0145_ _0148_ _0134_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1850_ g.bi_l\[63\]\[0\] g.g_y\[7\].g_x\[7\].t.r_v _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3520_ _0075_ _0077_ _1114_ _1111_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_21_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1953__A1 _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2333_ _1770_ _1794_ _1800_ _1413_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2402_ g.g_y\[7\].g_x\[2\].t.r_v _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3382_ _0796_ _0795_ _0812_ _0815_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3451_ net35 _1747_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2264_ _1742_ _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2195_ _1679_ _1680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_4003_ g.g_y\[1\].g_x\[4\].t.out_sc _4003_/E g.g_y\[1\].g_x\[4\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_63_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ g.g_y\[0\].g_x\[4\].t.r_h _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3649_ _0354_ _0358_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3718_ _1044_ _1695_ _1045_ _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2672__A2 _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3621__A1 _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2112__A1 _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2415__A2 _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1902_ _1376_ _1383_ _1394_ _1396_ _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2951_ net52 g.bi_l\[22\]\[1\] g.g_y\[2\].g_x\[6\].t.r_d _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1833_ _1327_ _1300_ _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3503_ _1482_ _1485_ _1085_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2882_ _0308_ _0311_ _0486_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2316_ _1780_ _1779_ _1795_ _1771_ _1796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3296_ _0890_ _0910_ _0916_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3365_ _0977_ _0979_ _0980_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3434_ _0993_ _1038_ _1040_ g.g_y\[1\].g_x\[2\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2178_ _1632_ _1665_ g.g_y\[7\].g_x\[3\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2247_ _1378_ _1732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput24 net24 out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_31_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2590__A1 _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3150_ _0776_ _0778_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2032_ g.g_y\[7\].g_x\[4\].t.r_h _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2101_ _1585_ _1587_ _1588_ _1589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3081_ _0670_ _0465_ _0468_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_45_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2934_ _0573_ net14 _0575_ _0571_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_20_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3983_ g.g_y\[2\].g_x\[0\].t.w_dh _3983_/E _3983_/RN g.bi_l\[16\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2865_ g.g_y\[3\].g_x\[2\].t.r_h _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_60_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1816_ g.g_y\[0\].g_x\[7\].t.r_v _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2796_ g.bi_l\[20\]\[1\] net49 _0445_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3417_ _1006_ _1008_ _1025_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_0_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3348_ _0963_ net12 _0965_ _0552_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3279_ net36 g.bi_l\[9\]\[1\] g.g_y\[1\].g_x\[1\].t.r_d _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2315__A1 _1773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_59_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout127_I net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2581_ _0242_ _0243_ _0244_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2650_ _0301_ _0300_ _0309_ _0310_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_10_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3202_ _0790_ _0811_ _0817_ _0789_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3133_ _0563_ _0565_ _0568_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2015_ _1502_ _1504_ _1505_ _1506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3064_ g.bi_l\[20\]\[0\] g.g_y\[2\].g_x\[4\].t.r_h _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3966_ g.g_y\[2\].g_x\[3\].t.w_si net125 g.g_y\[2\].g_x\[3\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2917_ _0546_ _0560_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2848_ g.g_y\[3\].g_x\[2\].t.r_v _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3897_ g.g_y\[4\].g_x\[1\].t.out_sc _3897_/E g.g_y\[4\].g_x\[1\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_60_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2779_ _1775_ _0388_ _0430_ g.g_y\[4\].g_x\[6\].t.r_d _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_13_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3751_ net106 _3751_/E g.g_y\[7\].g_x\[6\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_3820_ g.g_y\[6\].g_x\[0\].t.w_si net116 g.g_y\[6\].g_x\[0\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2702_ g.g_y\[4\].g_x\[1\].t.r_v _0351_ _0359_ g.g_y\[5\].g_x\[1\].t.r_v _0360_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3682_ _0869_ _1244_ _0867_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2564_ _1751_ _0227_ _0228_ g.g_y\[5\].g_x\[6\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2495_ _0123_ _0113_ _0164_ _1353_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_50_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2633_ g.g_y\[4\].g_x\[2\].t.r_h _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_2_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4040__CLK net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3116_ _0734_ _0747_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3047_ net57 _0682_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3949_ net51 _3949_/E g.g_y\[2\].g_x\[6\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_68_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout92 g.g_y\[6\].g_x\[6\].t.out_sc net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout81 g.g_y\[5\].g_x\[5\].t.out_sc net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout70 g.g_y\[4\].g_x\[4\].t.out_sc net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2280_ _1367_ _1347_ _1358_ _1760_ _1761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__3485__A2 _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3803_ g.g_y\[6\].g_x\[4\].t.w_dh _3803_/E _3803_/RN g.bi_l\[52\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_59_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2996__A1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1995_ g.g_y\[0\].g_x\[5\].t.r_v _1482_ _1485_ _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2616_ _0043_ _0042_ _0050_ _0026_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3734_ _1106_ _1098_ _1122_ _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3645__S _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3665_ _0718_ _0720_ _0721_ _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_15_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2547_ g.g_y\[5\].g_x\[6\].t.r_h _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3596_ _0059_ _1174_ _0057_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2478_ _0146_ _1386_ _0147_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_7_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2401_ g.g_y\[6\].g_x\[2\].t.r_d _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2332_ _1565_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3381_ _0807_ _0806_ _0814_ _0791_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3450_ _0901_ _1049_ _1051_ _1054_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3458__A2 _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2263_ _1745_ _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2194_ g.g_y\[1\].g_x\[1\].t.r_v _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4002_ g.g_y\[1\].g_x\[4\].t.w_si net125 g.g_y\[1\].g_x\[4\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_63_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3579_ _1602_ _1622_ _1629_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ net31 g.bi_l\[4\]\[1\] _1468_ _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3648_ g.g_y\[5\].g_x\[0\].t.r_v _0152_ _0542_ _0556_ _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1944__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3717_ _0733_ _0749_ _1042_ _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3621__A2 _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3385__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2112__A2 _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1901_ net94 _1395_ _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1832_ g.g_y\[0\].g_x\[7\].t.out_sc _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_32_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2950_ _0591_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2881_ g.g_y\[4\].g_x\[1\].t.r_h _0526_ _0527_ g.g_y\[4\].g_x\[2\].t.r_h _0528_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__1935__C _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3502_ g.g_y\[0\].g_x\[3\].t.r_h _1098_ _1099_ _1470_ _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3433_ net37 _1039_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2315_ _1773_ _1774_ _1776_ _1780_ _1795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2246_ _1704_ _1722_ _1730_ _1674_ _1731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3295_ _0912_ _0915_ g.g_y\[1\].g_x\[2\].t.r_v _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3364_ _0955_ _0958_ _0953_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2177_ _1633_ _1635_ _1664_ _1540_ _1665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_31_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput25 net25 out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2100_ g.g_y\[0\].g_x\[3\].t.r_h _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3080_ g.g_y\[3\].g_x\[3\].t.r_h _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2031_ _1404_ _1428_ _1521_ _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3982_ net44 _3982_/E g.g_y\[2\].g_x\[0\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XANTENNA__3597__A1 _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1815_ _1307_ _1308_ _1309_ _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2933_ _0572_ _0576_ g.g_y\[4\].g_x\[0\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2795_ g.g_y\[2\].g_x\[4\].t.r_d _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_20_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2864_ _0452_ _0454_ _0510_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_40_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3416_ _1006_ _0859_ _0862_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_4_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2229_ g.bi_l\[48\]\[0\] g.g_y\[6\].g_x\[0\].t.r_h _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3347_ _0930_ _0920_ _0964_ _0597_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3278_ _0898_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2563__A2 _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2315__A2 _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3579__A1 _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2580_ g.bi_l\[36\]\[0\] g.g_y\[4\].g_x\[4\].t.r_h _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3201_ _0785_ _0788_ _0819_ _0827_ g.g_y\[2\].g_x\[6\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3063_ _0695_ _0696_ _0697_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3132_ _0718_ _0720_ _0763_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2014_ g.g_y\[6\].g_x\[5\].t.r_h _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_54_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3965_ net48 _3965_/E g.g_y\[2\].g_x\[3\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_72_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2778_ _0390_ _0413_ _0419_ _1775_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3896_ g.g_y\[4\].g_x\[1\].t.w_si net110 g.g_y\[4\].g_x\[1\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2916_ g.g_y\[3\].g_x\[0\].t.out_sc _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2847_ _0084_ _0493_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3742__A1 _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2784__A2 _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1831__I1 _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2536__A2 _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3750_ g.g_y\[7\].g_x\[7\].t.w_na _3750_/E _3750_/RN g.bi_l\[63\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2701_ _0354_ _0358_ g.g_y\[4\].g_x\[1\].t.r_v _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2632_ _0290_ _0292_ _0284_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3681_ g.g_y\[2\].g_x\[3\].t.r_h _0871_ _0872_ _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2563_ net80 _0072_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2494_ _1724_ _1728_ _0123_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3046_ _1444_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3115_ g.g_y\[2\].g_x\[1\].t.out_sc _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2463__A1 _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3948_ g.g_y\[2\].g_x\[7\].t.out_sc _3948_/E g.g_y\[2\].g_x\[7\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_18_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_36_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3879_ net69 _3879_/E g.g_y\[4\].g_x\[4\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XTAP_TAPCELL_ROW_69_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Left_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3126__B _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xfanout93 g.g_y\[6\].g_x\[6\].t.out_sc net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout82 g.g_y\[5\].g_x\[6\].t.out_sc net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3852__CLK net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout71 net72 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout60 g.g_y\[3\].g_x\[5\].t.out_sc net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_72_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3802_ net91 _3802_/E g.g_y\[6\].g_x\[4\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_1994_ _1475_ _1474_ _1483_ _1484_ _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2996__A2 _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3595_ g.g_y\[6\].g_x\[3\].t.r_h _0061_ _0062_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3733_ _0075_ _0077_ _1114_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2615_ _0276_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3664_ _0880_ _0705_ _0711_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2477_ g.bi_l\[48\]\[0\] g.g_y\[6\].g_x\[0\].t.r_v _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2546_ _0210_ _0212_ _0213_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3029_ g.g_y\[3\].g_x\[5\].t.r_h _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2987__A2 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_72_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4030__CLK net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2400_ _1751_ _0071_ _0073_ g.g_y\[6\].g_x\[3\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2331_ _1763_ _1769_ _0001_ _0009_ g.g_y\[6\].g_x\[6\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_46_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2262_ _1439_ _1745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3380_ _0276_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4001_ g.g_y\[1\].g_x\[4\].t.out_sc _4001_/E g.g_y\[1\].g_x\[4\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_2193_ _1674_ _1675_ _1677_ _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ g.g_y\[0\].g_x\[4\].t.r_d _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3716_ _0899_ _1049_ _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3578_ _1480_ _1157_ _1159_ _1160_ g.g_y\[7\].g_x\[5\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_43_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2529_ _0175_ _0183_ _0194_ _0196_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_30_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3647_ _0545_ _0562_ _0569_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ _1318_ _1324_ _1325_ _1326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1900_ g.g_y\[7\].g_x\[0\].t.r_d _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2880_ _0354_ _0358_ g.g_y\[4\].g_x\[1\].t.r_h _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3501_ _1595_ _1598_ g.g_y\[0\].g_x\[3\].t.r_h _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3432_ _1444_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3363_ _0957_ _0943_ _0949_ _0978_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2314_ _1771_ _1781_ _1791_ _1793_ _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2176_ _1636_ _1656_ _1663_ _1633_ _1664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2245_ _1704_ _1725_ _1729_ _1730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_20_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3294_ _0906_ _0905_ _0913_ _0914_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_23_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput26 net109 out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3119__A2 _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3309__B _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2030_ _1404_ _1431_ _1434_ _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_27_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3597__A2 _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2932_ _0573_ net14 _0575_ _0142_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3981_ net44 _3981_/E g.g_y\[2\].g_x\[0\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA__3936__CLK net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2021__A2 _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1814_ g.bi_l\[15\]\[0\] g.g_y\[1\].g_x\[7\].t.r_v _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_20_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2794_ _0443_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2863_ g.bi_l\[27\]\[0\] g.g_y\[3\].g_x\[3\].t.r_h _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3415_ _1021_ _1023_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3346_ _0751_ _0755_ _0930_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2159_ _1643_ _1644_ _1646_ _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2228_ _1710_ _1712_ _1703_ _1713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3277_ g.g_y\[1\].g_x\[1\].t.r_h _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2260__A2 _1743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3512__A2 _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3579__A2 _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3200_ _0824_ _0826_ _0785_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2013_ _1348_ _1349_ _1503_ _1504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__1801__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3062_ g.bi_l\[18\]\[0\] g.g_y\[2\].g_x\[2\].t.r_h _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3267__A1 _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3131_ _0718_ _0518_ _0521_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3964_ g.g_y\[2\].g_x\[4\].t.w_na _3964_/E _3964_/RN g.bi_l\[20\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3895_ g.g_y\[4\].g_x\[1\].t.out_sc _3895_/E g.g_y\[4\].g_x\[1\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_2915_ _0555_ _0558_ _0544_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2846_ _0081_ _0103_ _0492_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__3742__A2 _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2777_ _0386_ _0389_ _0421_ _0429_ g.g_y\[4\].g_x\[6\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_5_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3329_ g.bi_l\[16\]\[0\] g.g_y\[2\].g_x\[0\].t.r_v _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3412__B _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2970__C _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout132_I net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2562_ _0225_ _0226_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2631_ _1604_ _1605_ _0291_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2700_ _0357_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3680_ _0839_ _0857_ _0863_ _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2493_ _1353_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2463__A2 _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3114_ _0742_ _0744_ _0745_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3045_ _0679_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3878_ g.g_y\[4\].g_x\[5\].t.out_sc _3878_/E g.g_y\[4\].g_x\[5\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_3947_ g.g_y\[2\].g_x\[7\].t.out_sc _3947_/E g.g_y\[2\].g_x\[7\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_18_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3412__A1 _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2829_ g.g_y\[4\].g_x\[3\].t.r_h _0477_ _0478_ _0473_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_69_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout83 g.g_y\[5\].g_x\[7\].t.out_sc net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout94 g.g_y\[7\].g_x\[0\].t.out_sc net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 net73 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout50 g.g_y\[2\].g_x\[4\].t.out_sc net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout61 g.g_y\[3\].g_x\[6\].t.out_sc net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3317__B g.g_y\[3\].g_x\[0\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2142__A1 _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3801_ net90 _3801_/E g.g_y\[6\].g_x\[4\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1993_ g.g_y\[0\].g_x\[5\].t.r_d _1484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3732_ _1525_ _1282_ _1285_ _1286_ g.g_y\[0\].g_x\[4\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_70_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3594_ _0025_ _0047_ _0053_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2545_ _0155_ _0158_ _0153_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2614_ _1439_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3663_ _0253_ _1226_ _1228_ _1229_ g.g_y\[3\].g_x\[5\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_2_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2476_ _1384_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3028_ _0637_ _0664_ _0665_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2330_ _0006_ _0008_ _1763_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2261_ _1557_ _1740_ _1741_ _1744_ g.g_y\[7\].g_x\[1\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2192_ g.bi_l\[57\]\[0\] _1676_ _1677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4000_ g.g_y\[1\].g_x\[5\].t.w_na _4000_/E _4000_/RN g.bi_l\[13\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_20_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3091__A2 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ g.g_y\[0\].g_x\[4\].t.r_h _1467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_28_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3715_ _0977_ _0979_ _1050_ _0899_ _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3577_ _1454_ _1479_ _1486_ _1480_ _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2528_ _0175_ _0195_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3646_ _0295_ _1212_ _1214_ _1215_ g.g_y\[4\].g_x\[2\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3842__CLK net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2459_ g.g_y\[7\].g_x\[0\].t.r_v _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3992__CLK net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2896__A2 _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ g.g_y\[0\].g_x\[7\].t.r_h _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_52_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3500_ _1597_ _1579_ _1589_ _1097_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_2313_ _1771_ _1792_ _1793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3362_ _0957_ _0950_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3431_ _1036_ _1037_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2244_ _1728_ _1729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2175_ _1659_ _1662_ g.g_y\[7\].g_x\[2\].t.r_h _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3293_ g.g_y\[1\].g_x\[2\].t.r_d _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_63_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3629_ _0125_ _1722_ _0361_ _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1959_ _1297_ net2 _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3678__I1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3602__I1 _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2931_ _0536_ _0526_ _0574_ _0189_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3980_ g.g_y\[2\].g_x\[0\].t.w_si net114 g.g_y\[2\].g_x\[0\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2557__A1 _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1813_ g.bi_l\[15\]\[1\] net42 g.g_y\[1\].g_x\[7\].t.r_d _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2793_ g.g_y\[2\].g_x\[4\].t.r_v _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_20_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2862_ _0506_ _0507_ _0508_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3276_ _0893_ _0895_ _0896_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3345_ _0597_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3414_ _0880_ _0705_ _1022_ _1573_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2158_ g.bi_l\[50\]\[0\] _1645_ _1646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2227_ _1674_ _1675_ _1711_ _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2089_ _1573_ _1574_ _1576_ _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2787__A1 _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3028__A2 _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3130_ g.g_y\[3\].g_x\[1\].t.r_h _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2012_ g.bi_l\[54\]\[0\] g.g_y\[6\].g_x\[6\].t.r_h _1503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3061_ net46 g.bi_l\[18\]\[1\] g.g_y\[2\].g_x\[2\].t.r_d _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3267__A2 _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2845_ _0081_ _0105_ _0108_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_33_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3894_ g.g_y\[4\].g_x\[2\].t.w_na _3894_/E _3894_/RN g.bi_l\[34\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3963_ g.g_y\[2\].g_x\[4\].t.w_dh _3963_/E _3963_/RN g.bi_l\[20\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2914_ _0556_ _0143_ _0557_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2776_ _0426_ _0428_ _0386_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3328_ _0551_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3259_ _0880_ _0692_ _0706_ _0709_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_8_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3926__CLK net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2561_ _1780_ _1779_ _1795_ _1798_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2630_ g.bi_l\[43\]\[0\] g.g_y\[5\].g_x\[3\].t.r_v _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2492_ _0133_ _0160_ _0161_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2889__B _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout125_I net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3185__A1 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3113_ g.g_y\[2\].g_x\[1\].t.r_h _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3044_ _0441_ _0450_ _0464_ _0467_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_18_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3877_ g.g_y\[4\].g_x\[5\].t.out_sc _3877_/E g.g_y\[4\].g_x\[5\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2828_ _0308_ _0311_ g.g_y\[4\].g_x\[3\].t.r_h _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3946_ g.g_y\[2\].g_x\[7\].t.w_si net123 g.g_y\[2\].g_x\[7\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3412__A2 _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2759_ _0391_ _0411_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2526__I1 _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout73 g.g_y\[4\].g_x\[6\].t.out_sc net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout62 g.g_y\[3\].g_x\[7\].t.out_sc net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout51 g.g_y\[2\].g_x\[6\].t.out_sc net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout40 g.g_y\[1\].g_x\[5\].t.out_sc net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout84 g.g_y\[5\].g_x\[7\].t.out_sc net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout95 g.g_y\[7\].g_x\[0\].t.out_sc net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2142__A2 _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3800_ g.g_y\[6\].g_x\[4\].t.w_si net127 g.g_y\[6\].g_x\[4\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1992_ _1467_ _1469_ _1471_ _1475_ _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3731_ _1090_ _1092_ _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3662_ g.g_y\[4\].g_x\[5\].t.r_v _0252_ _0636_ _0253_ _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3593_ _1365_ _1169_ _1171_ _1172_ g.g_y\[6\].g_x\[6\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2613_ _0167_ _0272_ _0273_ _0275_ g.g_y\[5\].g_x\[5\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3508__B _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2544_ _0157_ _0140_ _0149_ _0211_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2475_ _0141_ _0143_ _0144_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_66_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3027_ _0235_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3929_ g.g_y\[3\].g_x\[3\].t.w_dh _3929_/E _3929_/RN g.bi_l\[27\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__2372__A2 _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3624__A2 _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3388__A1 _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1874__A1 _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2260_ net94 _1743_ _1744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2191_ g.g_y\[7\].g_x\[1\].t.r_v _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2142__B _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1975_ _1460_ _1464_ _1465_ _1466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3714_ _1575_ _1267_ _1269_ _1271_ g.g_y\[1\].g_x\[3\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3645_ _0523_ _0493_ _0084_ _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3576_ _1522_ _1158_ _1520_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2458_ _0127_ _0128_ g.g_y\[6\].g_x\[1\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2527_ g.g_y\[4\].g_x\[7\].t.out_sc _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2389_ _0056_ _0064_ g.g_y\[6\].g_x\[4\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4059_ net28 _4059_/E g.g_y\[0\].g_x\[0\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_61_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3611__B _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2312_ net82 _1792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3361_ _0953_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3292_ _0899_ _0900_ _0902_ _0906_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3430_ _0896_ _0895_ _0911_ _0914_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_69_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2174_ _1660_ _1650_ _1661_ _1637_ _1662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2243_ _1718_ _1717_ _1726_ _1727_ _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__3240__C _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2272__A1 _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1958_ _1448_ _1449_ _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1889_ g.g_y\[6\].g_x\[0\].t.r_v _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_43_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3628_ g.g_y\[4\].g_x\[1\].t.r_v _0351_ _0359_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3559_ _1147_ net7 _1148_ _3559_/ZN vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2566__A2 _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3515__A1 _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1852__I1 _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2930_ _0353_ _0357_ _0536_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2861_ g.bi_l\[25\]\[0\] g.g_y\[3\].g_x\[1\].t.r_h _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3832__CLK net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1812_ g.g_y\[1\].g_x\[7\].t.r_v _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_25_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2792_ g.g_y\[3\].g_x\[4\].t.r_d _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3413_ _0707_ _0710_ _0687_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2226_ g.bi_l\[57\]\[0\] g.g_y\[7\].g_x\[1\].t.r_v _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3344_ _0936_ _0960_ _0961_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3275_ g.g_y\[1\].g_x\[2\].t.r_v _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_67_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2245__A1 _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2157_ g.g_y\[6\].g_x\[2\].t.r_v _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2088_ g.bi_l\[11\]\[0\] _1575_ _1576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3678__S _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2548__A2 _1792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2720__A2 _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3060_ _0694_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2011_ _1499_ _1500_ _1501_ _1502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_58_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3727__A1 _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2913_ g.bi_l\[32\]\[0\] g.g_y\[4\].g_x\[0\].t.r_v _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3962_ net50 _3962_/E g.g_y\[2\].g_x\[4\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3893_ g.g_y\[4\].g_x\[2\].t.w_dh _3893_/E _3893_/RN g.bi_l\[34\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__2415__B _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2844_ g.g_y\[4\].g_x\[2\].t.r_d _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2775_ _0376_ _0384_ _0427_ _0201_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2209_ _1693_ _1673_ _1694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3327_ _1389_ _1390_ _0944_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3189_ _0807_ _0806_ _0814_ _0815_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3258_ _0687_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3718__A1 _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout118_I net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2560_ _1790_ _1789_ _1797_ _1771_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2491_ _1385_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3112_ _0694_ _0696_ _0743_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3043_ _0459_ _0458_ _0466_ _0442_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3945_ g.g_y\[2\].g_x\[7\].t.out_sc _3945_/E g.g_y\[2\].g_x\[7\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XANTENNA__2999__A2 _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2620__A1 _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3876_ g.g_y\[4\].g_x\[5\].t.w_si net113 g.g_y\[4\].g_x\[5\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2758_ net61 _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2827_ _0310_ _0293_ _0302_ _0476_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_18_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2689_ g.g_y\[4\].g_x\[1\].t.r_h _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_69_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4056__CLK net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout85 g.g_y\[6\].g_x\[0\].t.out_sc net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout96 g.g_y\[7\].g_x\[1\].t.out_sc net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout30 g.g_y\[0\].g_x\[2\].t.out_sc net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout52 g.g_y\[2\].g_x\[6\].t.out_sc net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout74 net75 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout41 g.g_y\[1\].g_x\[5\].t.out_sc net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout63 g.g_y\[3\].g_x\[7\].t.out_sc net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3987__D net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3592_ _0000_ _1768_ _1411_ _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2612_ net79 _0274_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1991_ _1465_ _1464_ _1481_ _1455_ _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3730_ _1283_ _1284_ _1470_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_41_Left_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3661_ _0669_ _1227_ _0667_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2543_ _0157_ _0150_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2474_ g.bi_l\[32\]\[0\] g.g_y\[4\].g_x\[0\].t.r_v _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_11_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3026_ _0639_ _0657_ _0663_ _0253_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__3094__A1 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3928_ net56 _3928_/E g.g_y\[3\].g_x\[3\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3859_ g.g_y\[5\].g_x\[1\].t.w_dh _3859_/E _3859_/RN g.bi_l\[41\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__3149__A2 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3388__A2 _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3560__A2 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2190_ g.bi_l\[57\]\[1\] net96 g.g_y\[7\].g_x\[1\].t.r_d _1675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1974_ g.g_y\[0\].g_x\[5\].t.r_v _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3575_ _1523_ _1547_ _1554_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3644_ _0529_ _1213_ _0295_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3713_ _1270_ _1026_ _0846_ _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2388_ _0057_ _0059_ _0063_ _1531_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_53_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2457_ net85 _1757_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2526_ _0187_ _0192_ _0193_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1865__A2 _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4058_ g.g_y\[0\].g_x\[1\].t.out_sc _4058_/E g.g_y\[0\].g_x\[1\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XTAP_TAPCELL_ROW_26_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3009_ g.g_y\[2\].g_x\[4\].t.r_h _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_69_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2311_ _1785_ _1789_ _1790_ _1791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3533__A2 _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2242_ g.g_y\[6\].g_x\[1\].t.r_d _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_3360_ g.g_y\[1\].g_x\[7\].t.r_h _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3291_ _0896_ _0895_ _0911_ _0891_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2173_ _1377_ _1379_ _1651_ _1660_ _1661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_25_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2272__A2 _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1957_ _1429_ _1409_ _1430_ _1405_ _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_28_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput18 net18 out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1888_ _1381_ _1382_ g.g_y\[7\].g_x\[0\].t.r_h _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3627_ _0366_ _1199_ _0364_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3558_ _1297_ net6 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2509_ g.g_y\[3\].g_x\[7\].t.r_d _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3489_ _1086_ _1087_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1811_ _1302_ _1304_ _1305_ _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2791_ _0440_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2860_ net53 g.bi_l\[25\]\[1\] g.g_y\[3\].g_x\[1\].t.r_d _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2801__I1 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3412_ _1567_ _1592_ _1020_ _1575_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_13_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3532__B _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2225_ _1707_ _1708_ _1709_ _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3343_ _0552_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3274_ _0497_ _0499_ _0894_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2156_ g.bi_l\[50\]\[1\] net88 g.g_y\[6\].g_x\[2\].t.r_d _1644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2087_ g.g_y\[1\].g_x\[3\].t.r_v _1575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2989_ net61 _0629_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2837__I _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ g.bi_l\[52\]\[0\] g.g_y\[6\].g_x\[4\].t.r_h _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3961_ net49 _3961_/E g.g_y\[2\].g_x\[4\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2912_ _0141_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3727__A2 _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2774_ _0200_ _0204_ _0376_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2843_ _0485_ _0489_ _0490_ g.g_y\[4\].g_x\[3\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3892_ net67 _3892_/E g.g_y\[4\].g_x\[2\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3326_ g.bi_l\[0\]\[0\] g.g_y\[0\].g_x\[0\].t.r_v _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2431__B _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2139_ g.g_y\[6\].g_x\[3\].t.r_d _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2208_ g.g_y\[0\].g_x\[1\].t.out_sc _1693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3188_ g.g_y\[1\].g_x\[6\].t.r_d _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__3663__A1 _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3257_ _0878_ _0700_ _0708_ _0688_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_48_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3718__A2 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2457__A2 _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2393__A1 _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2490_ _0135_ _0152_ _0159_ _0146_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2448__A2 _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3042_ _0481_ _0676_ _0677_ _0678_ g.g_y\[3\].g_x\[5\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3111_ g.bi_l\[18\]\[0\] g.g_y\[2\].g_x\[2\].t.r_h _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3875_ g.g_y\[4\].g_x\[5\].t.out_sc _3875_/E g.g_y\[4\].g_x\[5\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3944_ g.g_y\[3\].g_x\[0\].t.out_sc _3944_/E g.g_y\[3\].g_x\[0\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_2757_ _0404_ _0408_ _0409_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2826_ _0310_ _0303_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2688_ _0294_ _0296_ _0345_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_14_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3309_ _0885_ _0922_ _0924_ _0928_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2336__B _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout86 g.g_y\[6\].g_x\[0\].t.out_sc net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout97 g.g_y\[7\].g_x\[1\].t.out_sc net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout31 g.g_y\[0\].g_x\[4\].t.out_sc net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout42 net43 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout75 g.g_y\[5\].g_x\[1\].t.out_sc net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout64 net65 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout53 net54 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2246__B _1730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1990_ _1480_ _1458_ _1459_ _1465_ _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_15_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout130_I net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3591_ _0007_ _1170_ _1365_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2611_ _1742_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2542_ _0153_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3660_ _0670_ _0672_ _0673_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2473_ g.bi_l\[32\]\[1\] net64 _0142_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3025_ _0639_ _0659_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3858_ net74 _3858_/E g.g_y\[5\].g_x\[1\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3927_ net56 _3927_/E g.g_y\[3\].g_x\[3\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3789_ net92 _3789_/E g.g_y\[6\].g_x\[6\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_41_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2809_ g.g_y\[3\].g_x\[4\].t.r_h _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1973_ _1461_ _1462_ _1463_ _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_EDGE_ROW_23_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3712_ _1027_ _1029_ _1030_ _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2339__A1 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3574_ _1489_ _1509_ _1516_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4046__CLK net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2525_ g.g_y\[4\].g_x\[7\].t.r_h _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3643_ _0486_ _0477_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2387_ g.g_y\[6\].g_x\[3\].t.r_h _0061_ _0062_ _0057_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2456_ _0122_ _0124_ _0126_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4057_ g.g_y\[0\].g_x\[1\].t.out_sc _4057_/E g.g_y\[0\].g_x\[1\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3008_ _0643_ _0645_ _0638_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2502__A1 _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2310_ g.g_y\[5\].g_x\[6\].t.r_h _1790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2241_ _1352_ _1354_ _1714_ _1718_ _1726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2172_ g.g_y\[7\].g_x\[2\].t.r_h _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3290_ _1638_ _1639_ _0892_ _0896_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1956_ _1432_ _1420_ _1433_ _1426_ _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1887_ net17 _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3488_ _1465_ _1464_ _1481_ _1484_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3626_ _0210_ _0212_ _0367_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput19 net19 out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_3557_ net8 _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2508_ g.g_y\[3\].g_x\[7\].t.r_v _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2439_ _1727_ _1720_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2723__A1 _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3451__A2 _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1810_ g.bi_l\[63\]\[0\] g.g_y\[7\].g_x\[7\].t.r_v _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3203__A2 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2790_ g.g_y\[3\].g_x\[4\].t.r_v _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_4_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3411_ _1595_ _1598_ g.g_y\[0\].g_x\[3\].t.r_v _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_40_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3342_ _0938_ _0952_ _0959_ _0946_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2155_ _1642_ _1643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2224_ g.bi_l\[41\]\[0\] g.g_y\[5\].g_x\[1\].t.r_v _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3273_ g.bi_l\[18\]\[0\] _0889_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_36_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2086_ g.bi_l\[11\]\[1\] net38 g.g_y\[1\].g_x\[3\].t.r_d _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1939_ _1432_ _1420_ _1433_ _1405_ _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3609_ _0163_ _1184_ _1185_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2988_ _1742_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2181__A2 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3433__A2 _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3960_ g.g_y\[2\].g_x\[4\].t.w_si net123 g.g_y\[2\].g_x\[4\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2911_ _0551_ _0553_ _0554_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3891_ net66 _3891_/E g.g_y\[4\].g_x\[2\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_2773_ _0422_ _0424_ _0425_ g.g_y\[4\].g_x\[6\].t.r_h _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2842_ net67 _0380_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3256_ _0701_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3325_ _0941_ _0942_ g.g_y\[1\].g_x\[0\].t.r_h _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2069_ _1520_ _1522_ _1555_ _1518_ _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2138_ _1611_ _1613_ _1614_ _1618_ _1626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2207_ _1688_ _1690_ _1691_ _1692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3187_ _0798_ _0799_ _0801_ _0807_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3718__B _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3406__A2 _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3110_ _0597_ _0598_ _0741_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3041_ net58 _0629_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3874_ g.g_y\[4\].g_x\[6\].t.w_na _3874_/E _3874_/RN g.bi_l\[38\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2825_ _0422_ _0424_ _0474_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1959__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3943_ g.g_y\[3\].g_x\[0\].t.out_sc _3943_/E g.g_y\[3\].g_x\[0\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2756_ g.g_y\[3\].g_x\[6\].t.r_h _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2687_ g.bi_l\[34\]\[0\] g.g_y\[4\].g_x\[2\].t.r_h _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_5_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3308_ _1451_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3239_ _0839_ _0859_ _0862_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_52_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout87 g.g_y\[6\].g_x\[2\].t.out_sc net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout98 g.g_y\[7\].g_x\[2\].t.out_sc net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout32 g.g_y\[0\].g_x\[4\].t.out_sc net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout76 g.g_y\[5\].g_x\[2\].t.out_sc net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout43 g.g_y\[1\].g_x\[7\].t.out_sc net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout65 g.g_y\[4\].g_x\[0\].t.out_sc net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout54 g.g_y\[3\].g_x\[1\].t.out_sc net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_9_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3590_ _1752_ _1761_ _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2541_ g.g_y\[5\].g_x\[7\].t.r_h _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2610_ _0263_ _0265_ _0270_ _0261_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_50_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3563__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2472_ g.g_y\[4\].g_x\[0\].t.r_d _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout123_I net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3077__C _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3024_ _0653_ _0652_ _0660_ _0661_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3788_ g.g_y\[6\].g_x\[7\].t.out_sc _3788_/E g.g_y\[6\].g_x\[7\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_3857_ net75 _3857_/E g.g_y\[5\].g_x\[1\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_2808_ _0401_ _0402_ _0457_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_18_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3926_ g.g_y\[3\].g_x\[3\].t.w_si net114 g.g_y\[3\].g_x\[3\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2739_ g.g_y\[2\].g_x\[6\].t.r_v _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_6_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2596__A2 _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1972_ g.bi_l\[13\]\[0\] g.g_y\[1\].g_x\[5\].t.r_v _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3642_ g.g_y\[4\].g_x\[1\].t.r_h _0526_ _0527_ _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3711_ _1020_ _1268_ _1575_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2339__A2 _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3573_ _1302_ _1153_ _1155_ _1156_ g.g_y\[7\].g_x\[7\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2455_ _0125_ _1712_ _1723_ _1727_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3536__A1 _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2524_ _0189_ _0190_ _0191_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_11_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2386_ _1625_ _1628_ g.g_y\[6\].g_x\[3\].t.r_h _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4056_ g.g_y\[0\].g_x\[1\].t.w_si net129 g.g_y\[0\].g_x\[1\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3007_ _0234_ _0236_ _0644_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3909_ g.g_y\[3\].g_x\[7\].t.w_dh _3909_/E _3909_/RN g.bi_l\[31\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_6_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1961__S _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3802__D net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2171_ _1657_ _1641_ _1658_ _1654_ _1659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2240_ _1724_ _1725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_38_Left_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2715__B _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1955_ _1447_ net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1886_ _1377_ _1379_ _1380_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3625_ _1623_ _1195_ _1197_ _1198_ g.g_y\[5\].g_x\[3\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2438_ _1645_ _0110_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_47_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3487_ _1085_ _1474_ _1483_ _1455_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2507_ g.g_y\[4\].g_x\[7\].t.r_d _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3556_ _1143_ _1144_ _1146_ g.g_y\[0\].g_x\[0\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input16_I in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2369_ net79 _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4039_ net32 _4039_/E g.g_y\[0\].g_x\[4\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_62_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2723__A2 _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4036__CLK net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2962__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3272_ _1638_ _1639_ _0892_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3341_ _0955_ _0958_ _0938_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3410_ g.g_y\[1\].g_x\[3\].t.r_d _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input8_I in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2154_ g.g_y\[6\].g_x\[2\].t.r_v _1642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2223_ g.bi_l\[41\]\[1\] net74 g.g_y\[5\].g_x\[1\].t.r_d _1708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_36_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2085_ g.g_y\[1\].g_x\[3\].t.r_v _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_16_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2987_ _0615_ _0620_ _0625_ _0613_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_8_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1869_ _1337_ _1346_ _1363_ _1339_ _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1938_ _1421_ _1422_ _1423_ _1432_ _1433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3608_ _0163_ net16 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3539_ _1441_ _1130_ _1131_ g.g_y\[0\].g_x\[1\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2841_ _0487_ _0488_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2910_ g.bi_l\[16\]\[0\] g.g_y\[2\].g_x\[0\].t.r_v _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3890_ g.g_y\[4\].g_x\[2\].t.w_si net111 g.g_y\[4\].g_x\[2\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2772_ _0255_ _0258_ g.g_y\[4\].g_x\[5\].t.r_h _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2206_ g.g_y\[0\].g_x\[1\].t.r_h _1691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3255_ _0724_ _0875_ _0876_ _0877_ g.g_y\[2\].g_x\[4\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3324_ net11 _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2068_ _1487_ _1517_ _1457_ _1558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2137_ _1601_ _1609_ _1624_ _1603_ _1625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3186_ _0796_ _0795_ _0812_ _0791_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_48_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2926__A2 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3040_ _0667_ _0669_ _0674_ _0665_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_58_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3873_ g.g_y\[4\].g_x\[6\].t.w_dh _3873_/E _3873_/RN g.bi_l\[38\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2824_ _0422_ _0255_ _0258_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3942_ g.g_y\[3\].g_x\[0\].t.w_si net111 g.g_y\[3\].g_x\[0\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2755_ _0405_ _0406_ _0407_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2686_ _0189_ _0190_ _0343_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3169_ g.g_y\[1\].g_x\[6\].t.r_v _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3307_ _0889_ _0887_ _0926_ g.g_y\[2\].g_x\[2\].t.r_d _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3238_ _0853_ _0852_ _0860_ _0861_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_55_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout33 net34 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_1_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout55 g.g_y\[3\].g_x\[2\].t.out_sc net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout44 net45 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout88 g.g_y\[6\].g_x\[2\].t.out_sc net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout99 g.g_y\[7\].g_x\[2\].t.out_sc net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout77 g.g_y\[5\].g_x\[3\].t.out_sc net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout66 g.g_y\[4\].g_x\[2\].t.out_sc net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2540_ _0172_ _0206_ _0207_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout116_I net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3563__A2 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2471_ g.g_y\[4\].g_x\[0\].t.r_v _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__3315__A2 _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3023_ g.g_y\[2\].g_x\[5\].t.r_d _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3925_ net57 _3925_/E g.g_y\[3\].g_x\[3\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3787_ g.g_y\[6\].g_x\[7\].t.out_sc _3787_/E g.g_y\[6\].g_x\[7\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3856_ g.g_y\[5\].g_x\[1\].t.w_si net110 g.g_y\[5\].g_x\[1\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2807_ g.bi_l\[29\]\[0\] g.g_y\[3\].g_x\[5\].t.r_h _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2738_ g.g_y\[3\].g_x\[6\].t.r_d _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2669_ _0099_ _0098_ _0106_ _0082_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_6_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2538__B _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3572_ _1299_ _1329_ _1335_ _1302_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3536__A2 _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1971_ g.bi_l\[13\]\[1\] net40 g.g_y\[1\].g_x\[5\].t.r_d _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3641_ _0028_ _1208_ _1210_ _1211_ g.g_y\[4\].g_x\[4\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_3_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3710_ _1567_ _1592_ _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2385_ _1627_ _1610_ _1619_ _0060_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_2454_ _1704_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2523_ g.bi_l\[32\]\[0\] g.g_y\[4\].g_x\[0\].t.r_h _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput1 in[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4055_ g.g_y\[0\].g_x\[1\].t.out_sc _4055_/E g.g_y\[0\].g_x\[1\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_3006_ g.bi_l\[29\]\[0\] g.g_y\[3\].g_x\[5\].t.r_v _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3908_ net62 _3908_/E g.g_y\[3\].g_x\[7\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3839_ g.g_y\[5\].g_x\[5\].t.w_dh _3839_/E _3839_/RN g.bi_l\[45\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XTAP_TAPCELL_ROW_60_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2170_ _1643_ _1644_ _1646_ _1657_ _1658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1954_ g.bi_l\[63\]\[0\] _1418_ _1373_ _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3509__A2 _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1885_ g.bi_l\[57\]\[0\] g.g_y\[7\].g_x\[1\].t.r_h _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3624_ g.g_y\[6\].g_x\[3\].t.r_v _1622_ _0282_ _1623_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3555_ _1145_ net2 net3 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_31_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2437_ _0081_ _0103_ _0109_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2368_ _0040_ _0042_ _0043_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3486_ _1475_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2506_ _0173_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2299_ _1410_ _1412_ _1778_ _1779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4038_ g.g_y\[0\].g_x\[5\].t.out_sc _4038_/E g.g_y\[0\].g_x\[5\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_34_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2184__A1 _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3684__A1 _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2239__A2 _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2222_ _1706_ _1707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3271_ g.bi_l\[2\]\[0\] g.g_y\[0\].g_x\[2\].t.r_v _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3340_ _0937_ _0945_ _0956_ _0957_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_2084_ _1569_ _1570_ _1571_ _1572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2153_ _1638_ _1639_ _1640_ _1641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_36_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1937_ g.g_y\[7\].g_x\[6\].t.r_h _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_56_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2986_ _0581_ _0612_ _0177_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1868_ _1362_ _1342_ _1343_ _1337_ _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__1913__A1 g.bi_l\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3607_ _1183_ _0113_ _0123_ _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3538_ net28 _1445_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3469_ _0790_ _0813_ _0816_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_47_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3409__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2396__A1 _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2771_ _0257_ _0241_ _0249_ _0423_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_33_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2840_ _0285_ _0292_ _0307_ _0310_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xrotfpga2a_135 out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2205_ _1580_ _1582_ _1689_ _1690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3185_ _1406_ _1407_ _0792_ _0796_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3254_ net48 _0629_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3323_ _0898_ _0900_ _0940_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2136_ _1623_ _1605_ _1606_ _1601_ _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2067_ _1440_ _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2387__A1 g.g_y\[6\].g_x\[3\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2969_ _0583_ _0607_ _0610_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_8_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4026__CLK net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3941_ g.g_y\[3\].g_x\[0\].t.out_sc _3941_/E g.g_y\[3\].g_x\[0\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3872_ net73 _3872_/E g.g_y\[4\].g_x\[6\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_30_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2754_ g.bi_l\[31\]\[0\] g.g_y\[3\].g_x\[7\].t.r_h _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2823_ g.g_y\[4\].g_x\[4\].t.r_h _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2685_ g.bi_l\[32\]\[0\] g.g_y\[4\].g_x\[0\].t.r_h _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3306_ _0890_ _0910_ _0916_ _0889_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2119_ _1604_ _1605_ _1606_ _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3168_ _0392_ _0394_ _0794_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_1_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3237_ g.g_y\[1\].g_x\[4\].t.r_d _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xfanout89 g.g_y\[6\].g_x\[3\].t.out_sc net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout34 g.g_y\[0\].g_x\[6\].t.out_sc net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout78 g.g_y\[5\].g_x\[3\].t.out_sc net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout45 g.g_y\[2\].g_x\[0\].t.out_sc net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3099_ _0485_ _0730_ _0731_ g.g_y\[3\].g_x\[2\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout56 g.g_y\[3\].g_x\[3\].t.out_sc net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout67 g.g_y\[4\].g_x\[2\].t.out_sc net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3021__A2 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3635__I1 _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2835__A2 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3571__I0 _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2470_ _0138_ _0139_ g.g_y\[5\].g_x\[0\].t.r_h _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3022_ _0647_ _0648_ _0649_ _0653_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__3079__A2 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3924_ g.g_y\[3\].g_x\[4\].t.out_sc _3924_/E g.g_y\[3\].g_x\[4\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_3786_ g.g_y\[6\].g_x\[7\].t.w_si net118 g.g_y\[6\].g_x\[7\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2668_ _0167_ _0325_ _0326_ _0327_ g.g_y\[5\].g_x\[3\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3855_ net74 _3855_/E g.g_y\[5\].g_x\[1\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2737_ g.g_y\[3\].g_x\[6\].t.r_v _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2806_ _0452_ _0454_ _0455_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2599_ g.g_y\[5\].g_x\[5\].t.r_h _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3490__A2 _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ g.g_y\[1\].g_x\[5\].t.r_v _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3571_ _1403_ _1154_ _1373_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3640_ g.g_y\[5\].g_x\[4\].t.r_v _0047_ _0438_ _0028_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_43_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2522_ net65 g.bi_l\[32\]\[1\] g.g_y\[4\].g_x\[0\].t.r_d _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2384_ _1627_ _1620_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2453_ _0123_ _1717_ _1726_ _1705_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4054_ g.g_y\[0\].g_x\[2\].t.w_na _4054_/E _4054_/RN g.bi_l\[2\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3005_ _1461_ _1462_ _0642_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput2 in[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3838_ net81 _3838_/E g.g_y\[5\].g_x\[5\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3907_ net63 _3907_/E g.g_y\[3\].g_x\[7\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_6_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3769_ g.g_y\[7\].g_x\[3\].t.w_dh _3769_/E _3769_/RN g.bi_l\[59\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_14_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2577__I1 _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ _1441_ _1442_ _1443_ _1446_ g.g_y\[7\].g_x\[7\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1884_ net96 g.bi_l\[57\]\[1\] _1378_ _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3485_ _1477_ _0988_ _1083_ _1084_ g.g_y\[0\].g_x\[6\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3623_ _0318_ _1196_ _0316_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3554_ net9 _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_31_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2505_ g.g_y\[4\].g_x\[7\].t.r_v _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2298_ g.bi_l\[54\]\[0\] g.g_y\[6\].g_x\[6\].t.r_v _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2367_ g.g_y\[5\].g_x\[4\].t.r_h _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2436_ _0105_ _0108_ g.g_y\[5\].g_x\[2\].t.r_v _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4037_ g.g_y\[0\].g_x\[5\].t.out_sc _4037_/E g.g_y\[0\].g_x\[5\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_22_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2221_ g.g_y\[5\].g_x\[1\].t.r_v _1706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2152_ g.bi_l\[2\]\[0\] g.g_y\[0\].g_x\[2\].t.r_v _1640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3270_ g.g_y\[1\].g_x\[2\].t.r_d _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2083_ g.bi_l\[59\]\[0\] g.g_y\[7\].g_x\[3\].t.r_v _1571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_36_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1867_ _1340_ _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1936_ _1429_ _1409_ _1430_ _1426_ _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_44_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2985_ _0614_ _0626_ g.g_y\[3\].g_x\[7\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1913__A2 g.g_y\[0\].g_x\[6\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3468_ g.g_y\[0\].g_x\[6\].t.r_v _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3606_ _1725_ _1729_ _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3537_ _1128_ _1129_ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2419_ _0088_ _0090_ _0091_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3399_ _0800_ _1005_ _1010_ _0998_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3942__CLK net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3657__A2 _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrotfpga2a_136 out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2396__A2 _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2770_ _0257_ _0250_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3322_ g.bi_l\[9\]\[0\] g.g_y\[1\].g_x\[1\].t.r_h _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2135_ _1604_ _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2204_ g.bi_l\[2\]\[0\] _1583_ _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3184_ _0791_ _0797_ _0808_ _0810_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_0_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3253_ _0867_ _0869_ _0873_ _0865_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2066_ _1519_ _1556_ g.g_y\[7\].g_x\[5\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_14_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1919_ g.bi_l\[54\]\[0\] _1413_ _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_60_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2387__A2 _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2899_ g.g_y\[5\].g_x\[0\].t.r_v _0152_ _0542_ g.g_y\[4\].g_x\[0\].t.r_v _0543_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2968_ _0601_ _0600_ _0608_ _0609_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_4_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1822__A1 g.bi_l\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2378__A2 _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3871_ net72 _3871_/E g.g_y\[4\].g_x\[6\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XTAP_TAPCELL_ROW_18_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3940_ g.g_y\[3\].g_x\[1\].t.w_na _3940_/E _3940_/RN g.bi_l\[25\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2753_ net62 g.bi_l\[31\]\[1\] g.g_y\[3\].g_x\[7\].t.r_d _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2822_ _0439_ _0470_ _0471_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3318__A1 g.g_y\[3\].g_x\[0\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2684_ _0338_ _0340_ _0341_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3305_ _0885_ _0888_ _0918_ _0925_ g.g_y\[2\].g_x\[2\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_68_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2118_ g.bi_l\[43\]\[0\] g.g_y\[5\].g_x\[3\].t.r_v _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2049_ g.g_y\[7\].g_x\[3\].t.r_d _1540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3167_ g.bi_l\[22\]\[0\] _0789_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3098_ net54 _0682_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3236_ _0846_ _0847_ _0849_ _0853_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_52_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout79 g.g_y\[5\].g_x\[4\].t.out_sc net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout68 g.g_y\[4\].g_x\[3\].t.out_sc net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout46 g.g_y\[2\].g_x\[2\].t.out_sc net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout57 g.g_y\[3\].g_x\[3\].t.out_sc net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout35 g.g_y\[1\].g_x\[0\].t.out_sc net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2532__A2 _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__B _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3021_ _0638_ _0645_ _0658_ _0640_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_61_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3854_ net76 _3854_/E g.g_y\[5\].g_x\[2\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA__3539__A1 _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3923_ net58 _3923_/E g.g_y\[3\].g_x\[4\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2805_ g.bi_l\[27\]\[0\] g.g_y\[3\].g_x\[3\].t.r_h _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4016__CLK net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3785_ g.g_y\[6\].g_x\[7\].t.out_sc _3785_/E g.g_y\[6\].g_x\[7\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_2667_ g.g_y\[5\].g_x\[2\].t.out_sc _0274_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2736_ _1773_ _0388_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2598_ _0230_ _0260_ _0261_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_6_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3711__A1 _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3219_ g.bi_l\[20\]\[0\] g.g_y\[2\].g_x\[4\].t.r_v _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_17_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2886__I _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3570_ _1404_ _1428_ _1435_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout121_I net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2521_ _0188_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_11_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2383_ _0002_ _0004_ _0058_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2452_ _1718_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4053_ g.g_y\[0\].g_x\[2\].t.w_dh _4053_/E _4053_/RN g.bi_l\[2\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 in[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3004_ g.bi_l\[13\]\[0\] _0641_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3837_ net81 _3837_/E g.g_y\[5\].g_x\[5\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3768_ net100 _3768_/E g.g_y\[7\].g_x\[3\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3906_ g.g_y\[3\].g_x\[7\].t.w_si net112 g.g_y\[3\].g_x\[7\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3699_ _0971_ _1258_ _0585_ _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2719_ _1747_ _0373_ _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_69_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2726__A2 _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_2_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3151__A2 _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1952_ net107 _1445_ _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1883_ g.g_y\[7\].g_x\[1\].t.r_d _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3622_ _0319_ _0321_ _0322_ _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2965__A2 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2504_ g.g_y\[6\].g_x\[7\].t.r_v _1361_ _0171_ g.g_y\[5\].g_x\[7\].t.r_v _0172_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3484_ _1074_ _1079_ _1081_ _1452_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2435_ _0099_ _0098_ _0106_ _0107_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3553_ _1137_ _1140_ _1141_ _0013_ _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_24_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2297_ _1773_ _1774_ _1776_ _1777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2366_ _1782_ _1783_ _0041_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4036_ g.g_y\[0\].g_x\[5\].t.w_si net131 g.g_y\[0\].g_x\[5\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2220_ g.g_y\[6\].g_x\[1\].t.r_d _1705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2082_ g.bi_l\[59\]\[1\] net100 g.g_y\[7\].g_x\[3\].t.r_d _1570_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2151_ g.bi_l\[2\]\[1\] net29 g.g_y\[0\].g_x\[2\].t.r_d _1639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2984_ _0615_ _0620_ _0625_ _0177_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_16_9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1866_ _1339_ _1347_ _1358_ _1360_ _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_1935_ _1411_ _1412_ _1414_ _1429_ _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3605_ _0129_ _0131_ _0132_ _0146_ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_31_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2418_ g.g_y\[5\].g_x\[2\].t.r_v _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3467_ _1068_ net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3536_ _1044_ _1683_ _1696_ _1699_ _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3398_ _1006_ _1008_ _1009_ _0800_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_3_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3145__I _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2349_ _0024_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input14_I in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4019_ g.g_y\[1\].g_x\[1\].t.w_dh _4019_/E _4019_/RN g.bi_l\[9\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3290__A1 _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrotfpga2a_137 out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_53_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3042__A1 _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3252_ _0837_ _0864_ _0445_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3321_ g.g_y\[1\].g_x\[0\].t.r_d _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2065_ _1520_ _1522_ _1555_ _1457_ _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2134_ _1603_ _1610_ _1619_ _1621_ _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3183_ _0791_ _0809_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2203_ _1686_ _1321_ _1687_ _1688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input6_I in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3656__I0 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2967_ g.g_y\[2\].g_x\[7\].t.r_d _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1849_ _1340_ _1342_ _1343_ _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1918_ g.g_y\[6\].g_x\[6\].t.r_v _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3584__A2 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2898_ _0155_ _0158_ g.g_y\[5\].g_x\[0\].t.r_v _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_4_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3519_ _1659_ _1662_ g.g_y\[7\].g_x\[2\].t.r_v _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2847__A1 _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3272__A1 _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3870_ g.g_y\[4\].g_x\[6\].t.w_si net119 g.g_y\[4\].g_x\[6\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2821_ _0029_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3263__A1 _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3566__A2 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2752_ g.g_y\[3\].g_x\[7\].t.r_h _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2683_ g.g_y\[4\].g_x\[1\].t.r_v _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__3318__A2 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3235_ _0838_ _0844_ _0858_ _0840_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3304_ _0922_ _0924_ _0885_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3579__B _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2048_ g.g_y\[7\].g_x\[3\].t.r_h _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_2117_ g.bi_l\[43\]\[1\] net77 g.g_y\[5\].g_x\[3\].t.r_d _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3166_ _1406_ _1407_ _0792_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3097_ _0728_ _0729_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout69 g.g_y\[4\].g_x\[4\].t.out_sc net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3999_ g.g_y\[1\].g_x\[5\].t.w_dh _3999_/E _3999_/RN g.bi_l\[13\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
Xfanout58 g.g_y\[3\].g_x\[4\].t.out_sc net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout47 g.g_y\[2\].g_x\[2\].t.out_sc net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3932__CLK net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout36 g.g_y\[1\].g_x\[1\].t.out_sc net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2393__B _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3020_ _1461_ _1462_ _0642_ _0638_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3853_ net76 _3853_/E g.g_y\[5\].g_x\[2\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3784_ net94 _3784_/E g.g_y\[7\].g_x\[0\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_41_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3922_ g.g_y\[3\].g_x\[4\].t.w_si net112 g.g_y\[3\].g_x\[4\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2804_ net56 g.bi_l\[27\]\[1\] _0453_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_14_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2735_ _1770_ _1794_ _0387_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2597_ _1492_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2666_ _0316_ _0318_ _0323_ _0314_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3149_ _0777_ _0589_ _0606_ _0609_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3218_ _1525_ _1526_ _0841_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2450__A2 _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1952__A1 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2451_ _1564_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2520_ g.g_y\[4\].g_x\[0\].t.r_h _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout114_I net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2382_ _0002_ _1512_ _1515_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4052_ net29 _4052_/E g.g_y\[0\].g_x\[2\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3003_ g.g_y\[1\].g_x\[5\].t.r_v _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput4 in[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_62_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3905_ net63 _3905_/E g.g_y\[3\].g_x\[7\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3836_ g.g_y\[5\].g_x\[5\].t.w_si net118 g.g_y\[5\].g_x\[5\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3767_ net100 _3767_/E g.g_y\[7\].g_x\[3\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2718_ _0210_ _0138_ _0154_ _0157_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2761__B _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3698_ _1299_ _1329_ _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2649_ g.g_y\[4\].g_x\[3\].t.r_d _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_69_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3439__A1 _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4006__CLK net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3611__A1 _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1882_ g.g_y\[7\].g_x\[1\].t.r_h _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_3621_ _0285_ _0305_ _0312_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3552_ _1132_ _1134_ _1136_ _1320_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1951_ _1444_ _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2503_ g.g_y\[6\].g_x\[7\].t.r_v _1364_ _1368_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2365_ g.bi_l\[45\]\[0\] g.g_y\[5\].g_x\[5\].t.r_h _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3483_ _1069_ _1071_ _1073_ _1314_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2434_ g.g_y\[5\].g_x\[2\].t.r_d _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_63_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4035_ g.g_y\[0\].g_x\[5\].t.out_sc _4035_/E g.g_y\[0\].g_x\[5\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_2296_ g.bi_l\[38\]\[0\] _1775_ _1776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_39_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3587__B _1730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3819_ net86 _3819_/E g.g_y\[6\].g_x\[0\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_30_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2341__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2081_ g.g_y\[7\].g_x\[3\].t.r_v _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2150_ g.g_y\[0\].g_x\[2\].t.r_v _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_17_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1934_ g.g_y\[7\].g_x\[6\].t.r_v _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_44_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2983_ _0621_ _0623_ _0624_ g.g_y\[3\].g_x\[7\].t.r_h _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_71_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1865_ _1339_ _1359_ _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3604_ _0135_ _0152_ _0159_ _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3535_ _1127_ _1690_ _1698_ _1673_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_3_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3466_ _1065_ _1067_ g.g_y\[0\].g_x\[7\].t.r_h _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2417_ _1642_ _1644_ _0089_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2348_ g.g_y\[5\].g_x\[4\].t.r_v _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3397_ _0859_ _0862_ g.g_y\[1\].g_x\[4\].t.r_h _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2279_ _1367_ _1359_ _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1921__I1 _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4018_ net36 _4018_/E g.g_y\[1\].g_x\[1\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_47_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2617__A2 _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3290__A2 _1639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Left_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2202_ g.bi_l\[0\]\[0\] _1322_ _1687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3182_ g.g_y\[1\].g_x\[6\].t.out_sc _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3251_ _0866_ _0874_ g.g_y\[2\].g_x\[4\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3320_ _0937_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2133_ _1603_ _1620_ _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2064_ _1523_ _1547_ _1554_ _1520_ _1555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_53_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2856__A2 _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1917_ g.bi_l\[54\]\[1\] net92 g.g_y\[6\].g_x\[6\].t.r_d _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2966_ _0591_ _0593_ _0594_ _0601_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2897_ _0540_ _0541_ g.g_y\[4\].g_x\[1\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1848_ g.bi_l\[47\]\[0\] g.g_y\[5\].g_x\[7\].t.r_v _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3518_ _0890_ _0910_ _1112_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_71_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2847__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3449_ _1041_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3272__A2 _1639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2854__B _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2751_ _0401_ _0402_ _0403_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2820_ _0441_ _0463_ _0469_ _0028_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_53_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2682_ _1707_ _1708_ _0339_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3165_ g.bi_l\[6\]\[0\] g.g_y\[0\].g_x\[6\].t.r_v _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3234_ _1525_ _1526_ _0841_ _0838_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3303_ _0878_ _0871_ _0923_ _0695_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2047_ _1421_ _1422_ _1537_ _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2116_ g.g_y\[5\].g_x\[3\].t.r_v _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_52_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3254__A2 _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3096_ _0504_ _0503_ _0517_ _0520_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_9_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout37 g.g_y\[1\].g_x\[1\].t.out_sc net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3595__B _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout59 g.g_y\[3\].g_x\[5\].t.out_sc net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3998_ net41 _3998_/E g.g_y\[1\].g_x\[5\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2949_ g.g_y\[2\].g_x\[6\].t.r_h _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_4_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout48 g.g_y\[2\].g_x\[3\].t.out_sc net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_9_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2359__I1 _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3921_ net58 _3921_/E g.g_y\[3\].g_x\[4\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_2734_ _1770_ _1796_ _1799_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3783_ net95 _3783_/E g.g_y\[7\].g_x\[0\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3852_ g.g_y\[5\].g_x\[2\].t.w_si net117 g.g_y\[5\].g_x\[2\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2803_ g.g_y\[3\].g_x\[3\].t.r_d _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_14_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2596_ _0232_ _0252_ _0259_ _1510_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2665_ _0283_ _0313_ _0037_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3635__S _1773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3217_ g.bi_l\[4\]\[0\] g.g_y\[0\].g_x\[4\].t.r_v _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3148_ _0583_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3079_ _0685_ _0712_ _0713_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1952__A2 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2381_ g.g_y\[6\].g_x\[4\].t.r_h _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2450_ _1720_ _0010_ _0120_ _0121_ g.g_y\[6\].g_x\[2\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4051_ net29 _4051_/E g.g_y\[0\].g_x\[2\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3002_ g.g_y\[2\].g_x\[5\].t.r_d _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput5 in[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_62_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3904_ g.g_y\[4\].g_x\[0\].t.w_na _3904_/E _3904_/RN g.bi_l\[32\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3835_ net80 _3835_/E g.g_y\[5\].g_x\[5\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3766_ g.g_y\[7\].g_x\[3\].t.w_si net128 g.g_y\[7\].g_x\[3\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2717_ _0135_ _0145_ _0156_ _0136_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3697_ _0777_ _0605_ _0973_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2579_ net69 g.bi_l\[36\]\[1\] g.g_y\[4\].g_x\[4\].t.r_d _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2648_ _0294_ _0296_ _0297_ _0301_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_65_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3611__A2 _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1950_ _1439_ _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2502_ _0167_ _0168_ _0169_ _0170_ g.g_y\[6\].g_x\[0\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3620_ _1510_ _1191_ _1193_ _1194_ g.g_y\[5\].g_x\[5\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1881_ g.g_y\[7\].g_x\[0\].t.r_d _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3551_ _1138_ _1142_ g.g_y\[0\].g_x\[0\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3482_ _1075_ _1082_ g.g_y\[0\].g_x\[6\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2364_ _0036_ _0038_ _0039_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2433_ _0093_ _0094_ _0095_ _0099_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_63_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4034_ g.g_y\[0\].g_x\[6\].t.w_na _4034_/E _4034_/RN g.bi_l\[6\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XTAP_TAPCELL_ROW_39_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2295_ g.g_y\[4\].g_x\[6\].t.r_v _1775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3818_ g.g_y\[6\].g_x\[1\].t.out_sc _3818_/E g.g_y\[6\].g_x\[1\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3749_ g.g_y\[7\].g_x\[7\].t.w_dh _3749_/E _3749_/RN g.bi_l\[63\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XTAP_TAPCELL_ROW_30_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2341__A2 _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output20_I net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2080_ g.g_y\[0\].g_x\[3\].t.r_d _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_36_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1933_ _1405_ _1416_ _1425_ _1427_ _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__2399__A2 _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2982_ _0415_ _0418_ g.g_y\[3\].g_x\[6\].t.r_h _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1864_ g.g_y\[6\].g_x\[7\].t.out_sc _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3603_ _1612_ _1177_ _1179_ _1180_ g.g_y\[6\].g_x\[2\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3465_ _1333_ _1312_ _1326_ _1066_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_3534_ _1691_ _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2278_ _1364_ _1368_ _1759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2347_ _0019_ _0021_ _0022_ g.g_y\[6\].g_x\[4\].t.r_v _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2416_ g.bi_l\[50\]\[0\] g.g_y\[6\].g_x\[2\].t.r_v _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3396_ _0861_ _0845_ _0854_ _1007_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4017_ net36 _4017_/E g.g_y\[1\].g_x\[1\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_62_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3587__A1 _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2132_ net89 _1620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_49_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2201_ _1319_ _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3181_ _0802_ _0806_ _0807_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3250_ _0867_ _0869_ _0873_ _0445_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2063_ _1550_ _1553_ g.g_y\[7\].g_x\[4\].t.r_h _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_71_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3569__A1 _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1847_ g.bi_l\[47\]\[1\] net83 _1341_ _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1916_ _1410_ _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2965_ _0582_ _0589_ _0606_ _0584_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2896_ net64 _1757_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3592__I1 _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3517_ _0890_ _0912_ _0915_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3448_ _1043_ _1046_ _1041_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3379_ _0992_ net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_55_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2681_ g.bi_l\[41\]\[0\] g.g_y\[5\].g_x\[1\].t.r_v _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2750_ g.bi_l\[29\]\[0\] g.g_y\[3\].g_x\[5\].t.r_h _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2870__B _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3302_ _0707_ _0710_ _0878_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2115_ g.g_y\[6\].g_x\[3\].t.r_d _1603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3164_ g.g_y\[1\].g_x\[6\].t.r_d _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3233_ _0840_ _0845_ _0854_ _0856_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_3095_ _0512_ _0511_ _0519_ _0496_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2046_ g.bi_l\[61\]\[0\] g.g_y\[7\].g_x\[5\].t.r_h _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_52_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout27 g.g_y\[0\].g_x\[0\].t.out_sc net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3997_ net40 _3997_/E g.g_y\[1\].g_x\[5\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
Xfanout49 net50 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout38 g.g_y\[1\].g_x\[3\].t.out_sc net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_17_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2948_ _0587_ _0589_ _0582_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2879_ _0356_ _0342_ _0348_ _0525_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_13_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3851_ net76 _3851_/E g.g_y\[5\].g_x\[2\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3920_ g.g_y\[3\].g_x\[5\].t.w_na _3920_/E _3920_/RN g.bi_l\[29\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2664_ _0315_ _0324_ g.g_y\[5\].g_x\[3\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3782_ g.g_y\[7\].g_x\[0\].t.w_si net119 g.g_y\[7\].g_x\[0\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2733_ g.g_y\[4\].g_x\[6\].t.r_d _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2802_ g.g_y\[3\].g_x\[3\].t.r_h _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_14_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2595_ _0232_ _0255_ _0258_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_1_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3147_ _0775_ _0600_ _0608_ _0584_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3078_ _0453_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3216_ g.g_y\[1\].g_x\[4\].t.r_d _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2029_ g.g_y\[7\].g_x\[5\].t.r_h _1520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2986__A2 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2380_ _0023_ _0054_ _0055_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3154__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ g.g_y\[0\].g_x\[2\].t.w_si net129 g.g_y\[0\].g_x\[2\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3001_ _0638_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput6 in[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3701__I1 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3834_ g.g_y\[5\].g_x\[6\].t.out_sc _3834_/E g.g_y\[5\].g_x\[6\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_62_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3903_ g.g_y\[4\].g_x\[0\].t.w_dh _3903_/E _3903_/RN g.bi_l\[32\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__2968__A2 _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3765_ net101 _3765_/E g.g_y\[7\].g_x\[3\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2716_ _0150_ _0010_ _0371_ _0372_ g.g_y\[5\].g_x\[1\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2647_ _0284_ _0292_ _0307_ _0286_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3696_ _0946_ _1251_ _1252_ _1256_ g.g_y\[2\].g_x\[0\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2578_ g.g_y\[4\].g_x\[4\].t.r_h _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3384__A2 _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2895__A1 _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1880_ _1374_ _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2501_ net83 _1743_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3481_ _1314_ _1079_ _1081_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_51_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3550_ _1320_ _1140_ _1141_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_3_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3375__A2 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ g.g_y\[0\].g_x\[6\].t.w_dh _4033_/E _4033_/RN g.bi_l\[6\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2363_ g.bi_l\[43\]\[0\] g.g_y\[5\].g_x\[3\].t.r_h _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2432_ _0091_ _0090_ _0104_ _0082_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2294_ g.bi_l\[38\]\[1\] net71 g.g_y\[4\].g_x\[6\].t.r_d _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3748_ net109 _3748_/E g.g_y\[7\].g_x\[7\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_62_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3817_ g.g_y\[6\].g_x\[1\].t.out_sc _3817_/E g.g_y\[6\].g_x\[1\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_30_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3679_ _0592_ _1239_ _1241_ _1242_ g.g_y\[2\].g_x\[6\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_6_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1863_ _1351_ _1356_ _1357_ _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1932_ _1426_ net106 _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_68_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3602_ _0110_ _0079_ _1643_ _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_44_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2981_ _0417_ _0400_ _0410_ _0622_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_16_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3464_ _1327_ _1333_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3533_ _1693_ _0122_ _1125_ _1126_ g.g_y\[0\].g_x\[2\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2415_ _0084_ _0085_ _0087_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2277_ _1751_ _1755_ _1758_ g.g_y\[6\].g_x\[7\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2346_ _1535_ _1550_ _1553_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_35_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3395_ _0861_ _0855_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4016_ g.g_y\[1\].g_x\[1\].t.w_si net122 g.g_y\[1\].g_x\[1\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3587__A2 _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2131_ _1615_ _1617_ _1618_ _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2062_ _1551_ _1538_ _1552_ _1524_ _1553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_49_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2200_ _1678_ _1683_ _1684_ _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3180_ g.g_y\[1\].g_x\[6\].t.r_h _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__3569__A2 _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2964_ _1307_ _1308_ _0586_ _0582_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1846_ g.g_y\[5\].g_x\[7\].t.r_d _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1915_ g.g_y\[6\].g_x\[6\].t.r_v _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2895_ _0122_ _0537_ _0539_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_4_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3516_ g.g_y\[0\].g_x\[2\].t.r_v _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3378_ g.bi_l\[15\]\[0\] _0804_ _0976_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3447_ _1041_ _1047_ _1052_ g.g_y\[1\].g_x\[1\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2329_ _1752_ _1761_ _0007_ _1365_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_input12_I in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3496__A1 _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1982__A1 g.bi_l\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2680_ _0335_ _0336_ _0337_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3232_ _0840_ _0855_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3301_ g.g_y\[2\].g_x\[1\].t.r_h _0920_ _0921_ g.g_y\[2\].g_x\[2\].t.r_h _0922_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2045_ _1528_ _1534_ _1535_ _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2114_ _1601_ _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3163_ g.g_y\[1\].g_x\[6\].t.r_v _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input4_I in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3094_ _0724_ _0725_ _0726_ _0727_ g.g_y\[3\].g_x\[3\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_72_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout28 g.g_y\[0\].g_x\[0\].t.out_sc net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2947_ _0176_ _0178_ _0588_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3996_ g.g_y\[1\].g_x\[5\].t.w_si net126 g.g_y\[1\].g_x\[5\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_17_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout39 g.g_y\[1\].g_x\[3\].t.out_sc net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1829_ _1319_ _1321_ _1323_ _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_32_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2878_ _0356_ _0349_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3026__C _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2141__A1 _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2444__A2 _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3781_ net95 _3781_/E g.g_y\[7\].g_x\[0\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3850_ g.g_y\[5\].g_x\[3\].t.w_na _3850_/E _3850_/RN g.bi_l\[43\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__3641__A1 _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2801_ _0448_ _0450_ _0440_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2663_ _0316_ _0318_ _0323_ _0037_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2732_ _0385_ net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2594_ _0248_ _0247_ _0256_ _0257_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_1_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2900__I g.g_y\[3\].g_x\[0\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3215_ _0838_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_65_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2028_ _1487_ _1517_ _1518_ _1519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_59_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3146_ _0601_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3077_ _0687_ _0705_ _0711_ _0306_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_72_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3979_ net45 _3979_/E g.g_y\[2\].g_x\[0\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_68_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3000_ g.g_y\[2\].g_x\[5\].t.r_v _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_19_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 in[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3833_ net82 _3833_/E g.g_y\[5\].g_x\[6\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3764_ net102 _3764_/E g.g_y\[7\].g_x\[4\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3902_ net64 _3902_/E g.g_y\[4\].g_x\[0\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_2715_ _0332_ _0360_ _0362_ _0013_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2577_ _0238_ _0240_ _0231_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3695_ _0963_ _1254_ _1255_ _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2646_ _0306_ _0288_ _0289_ _0284_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_69_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3605__A1 _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3129_ _0758_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2026__B _1516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2647__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3072__A2 _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3480_ _1060_ _1067_ _1080_ _1313_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2500_ _0133_ _0160_ _1385_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2431_ _0084_ _0085_ _0087_ _0091_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4032_ net33 _4032_/E g.g_y\[0\].g_x\[6\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_2362_ net77 g.bi_l\[43\]\[1\] _0037_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2293_ _1772_ _1773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_22_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3747_ net108 _3747_/E g.g_y\[7\].g_x\[7\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_62_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3816_ g.g_y\[6\].g_x\[1\].t.w_si net117 g.g_y\[6\].g_x\[1\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_30_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3678_ _0818_ _0787_ _0393_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2629_ _0287_ _0288_ _0289_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2980_ _0417_ _0411_ _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1862_ g.g_y\[6\].g_x\[7\].t.r_h _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_1931_ g.g_y\[7\].g_x\[6\].t.r_d _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3601_ _0116_ _1178_ _1612_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_44_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput10 in[2] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3463_ _1331_ _1334_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3532_ _1116_ _1121_ _1123_ _1452_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2414_ g.bi_l\[34\]\[0\] _0086_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3394_ g.g_y\[1\].g_x\[4\].t.r_h _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2276_ net92 _1757_ _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2345_ _1545_ _1536_ _1544_ _0020_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_4015_ net37 _4015_/E g.g_y\[1\].g_x\[1\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_62_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2538__A1 _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2130_ g.g_y\[6\].g_x\[3\].t.r_h _1618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2061_ _1539_ _1541_ _1542_ _1551_ _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_49_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1914_ _1406_ _1407_ _1408_ _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2963_ _0584_ _0590_ _0602_ _0604_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_1845_ g.g_y\[5\].g_x\[7\].t.r_v _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3515_ _1441_ _1109_ _1110_ g.g_y\[0\].g_x\[3\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_31_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2894_ _0538_ _0340_ _0352_ _0356_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_69_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2328_ _1364_ _1368_ _1752_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3377_ _0809_ _0988_ _0990_ _0991_ g.g_y\[1\].g_x\[7\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3446_ _0901_ _1049_ _1051_ _1041_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2259_ _1742_ _1743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_40_Left_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3496__A2 _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3162_ g.g_y\[2\].g_x\[6\].t.r_v _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3554__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3231_ g.g_y\[1\].g_x\[4\].t.out_sc _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3300_ _0752_ _0756_ g.g_y\[2\].g_x\[1\].t.r_h _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2044_ g.g_y\[7\].g_x\[4\].t.r_v _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2113_ g.g_y\[6\].g_x\[3\].t.r_v _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3093_ g.g_y\[3\].g_x\[2\].t.out_sc _0629_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout29 g.g_y\[0\].g_x\[2\].t.out_sc net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2946_ g.bi_l\[31\]\[0\] g.g_y\[3\].g_x\[7\].t.r_v _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3995_ net41 _3995_/E g.g_y\[1\].g_x\[5\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2877_ _0086_ _0523_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ g.bi_l\[0\]\[0\] _1322_ _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_13_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3429_ _0906_ _0905_ _0913_ _0891_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_51_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3166__A1 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3780_ g.g_y\[7\].g_x\[1\].t.w_na _3780_/E _3780_/RN g.bi_l\[57\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2800_ _0027_ _0030_ _0449_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2731_ _0382_ _0384_ g.g_y\[4\].g_x\[7\].t.r_h _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_14_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2662_ _0319_ _0321_ _0322_ _0316_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_41_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2593_ g.g_y\[4\].g_x\[5\].t.r_d _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_1_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3145_ _0276_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3214_ g.g_y\[1\].g_x\[4\].t.r_v _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_65_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2027_ _1457_ _1518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3076_ _0687_ _0707_ _0710_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_72_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2929_ _0189_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3978_ g.g_y\[2\].g_x\[1\].t.out_sc _3978_/E g.g_y\[2\].g_x\[1\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_9_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3318__B _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 in[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3614__A2 _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3901_ net64 _3901_/E g.g_y\[4\].g_x\[0\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_19_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3763_ net102 _3763_/E g.g_y\[7\].g_x\[4\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3832_ g.g_y\[5\].g_x\[6\].t.w_si net118 g.g_y\[5\].g_x\[6\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2714_ _0364_ _0366_ _0368_ _0370_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3694_ _0963_ net12 _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2576_ _1491_ _1493_ _0239_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_10_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2645_ _0287_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3128_ _0538_ _0351_ _0759_ _0335_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_65_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3605__A2 _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3059_ g.g_y\[2\].g_x\[2\].t.r_h _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2361_ g.g_y\[5\].g_x\[3\].t.r_d _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2430_ _0082_ _0092_ _0100_ _0102_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_4031_ net34 _4031_/E g.g_y\[0\].g_x\[6\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2292_ g.g_y\[4\].g_x\[6\].t.r_v _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_63_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3746_ g.g_y\[7\].g_x\[7\].t.w_si net127 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3815_ g.g_y\[6\].g_x\[1\].t.out_sc _3815_/E g.g_y\[6\].g_x\[1\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XTAP_TAPCELL_ROW_30_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3677_ _0825_ _1240_ _0592_ _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2559_ _0224_ net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2628_ g.bi_l\[27\]\[0\] g.g_y\[3\].g_x\[3\].t.r_v _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_38_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ _1420_ _1424_ g.g_y\[7\].g_x\[6\].t.r_h _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_44_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2556__A2 _1743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3600_ _0068_ _0061_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1861_ _1353_ _1354_ _1355_ _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3531_ _1111_ _1113_ _1115_ _1581_ _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3557__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 in[3] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2344_ _1524_ net103 _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_58_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3462_ _0993_ _1063_ _1064_ g.g_y\[0\].g_x\[7\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3393_ _0982_ _0984_ _1004_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3108__I1 _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2413_ g.g_y\[4\].g_x\[2\].t.r_v _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2275_ _1756_ _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4014_ g.g_y\[1\].g_x\[2\].t.out_sc _4014_/E g.g_y\[1\].g_x\[2\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_15_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3729_ g.g_y\[0\].g_x\[3\].t.r_h _1098_ _1099_ _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2538__A2 _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2786__A2 _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2060_ g.g_y\[7\].g_x\[4\].t.r_h _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_49_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1913_ g.bi_l\[6\]\[0\] g.g_y\[0\].g_x\[6\].t.r_v _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2962_ _0584_ _0603_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2893_ _0341_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1844_ g.g_y\[6\].g_x\[7\].t.r_d _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3726__A1 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3514_ net30 _1039_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3445_ _0977_ _0979_ _1050_ _0901_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2327_ _0002_ _0004_ _0005_ g.g_y\[6\].g_x\[6\].t.r_h _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3376_ _0970_ _0972_ _0974_ _0928_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2258_ _1438_ _1742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2189_ g.g_y\[7\].g_x\[1\].t.r_v _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_47_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3717__A1 _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2456__A1 _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2112_ _1567_ _1592_ _1599_ g.g_y\[7\].g_x\[3\].t.r_v _1600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3161_ _0393_ _0787_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3230_ _0850_ _0852_ _0853_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2043_ _1530_ _1532_ _1533_ _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3092_ _0715_ _0717_ _0722_ _0713_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_72_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1827_ g.g_y\[0\].g_x\[0\].t.r_h _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2945_ _1307_ _1308_ _0586_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3994_ g.g_y\[1\].g_x\[6\].t.out_sc _3994_/E g.g_y\[1\].g_x\[6\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2876_ _0495_ _0516_ _0522_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_17_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3428_ _0908_ _0988_ _1034_ _1035_ g.g_y\[1\].g_x\[3\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_68_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3359_ _0972_ _0974_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_51_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2989__A2 _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2661_ _0105_ _0108_ g.g_y\[5\].g_x\[2\].t.r_h _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2730_ _0203_ _0183_ _0194_ _0383_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_14_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2592_ _0242_ _0243_ _0244_ _0248_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3565__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2668__A1 _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3213_ g.g_y\[3\].g_x\[4\].t.r_v _0463_ _0836_ g.g_y\[2\].g_x\[4\].t.r_v _0837_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3075_ _0701_ _0700_ _0708_ _0709_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3144_ _0603_ _1746_ _0773_ g.g_y\[3\].g_x\[0\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_65_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2026_ _1489_ _1509_ _1516_ _1480_ _1517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3977_ g.g_y\[2\].g_x\[1\].t.out_sc _3977_/E g.g_y\[2\].g_x\[1\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA__2840__A1 _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2928_ _0543_ _0570_ _0571_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2859_ g.g_y\[3\].g_x\[1\].t.r_h _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_5_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput9 in[1] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1873__A2 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3831_ net82 _3831_/E g.g_y\[5\].g_x\[6\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XTAP_TAPCELL_ROW_62_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3900_ g.g_y\[4\].g_x\[0\].t.w_si net110 g.g_y\[4\].g_x\[0\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2822__A1 _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3762_ g.g_y\[7\].g_x\[4\].t.w_si net128 g.g_y\[7\].g_x\[4\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2713_ _0332_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2644_ _0286_ _0293_ _0302_ _0304_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_2_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3693_ _1253_ _0920_ _0930_ _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2575_ g.bi_l\[45\]\[0\] g.g_y\[5\].g_x\[5\].t.r_v _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3127_ _0354_ _0358_ _0538_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3058_ _0690_ _0692_ _0686_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3613__I0 _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2009_ net90 g.bi_l\[52\]\[1\] g.g_y\[6\].g_x\[4\].t.r_d _1500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2291_ g.g_y\[5\].g_x\[6\].t.r_d _1771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2360_ g.g_y\[5\].g_x\[3\].t.r_h _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_63_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4030_ g.g_y\[0\].g_x\[6\].t.w_si net130 g.g_y\[0\].g_x\[6\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2271__A2 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3814_ g.g_y\[6\].g_x\[2\].t.w_na _3814_/E _3814_/RN g.bi_l\[50\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XTAP_TAPCELL_ROW_22_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3745_ net108 _3745_/E g.g_y\[7\].g_x\[7\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_42_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3676_ _0775_ _0783_ _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2627_ g.bi_l\[27\]\[1\] net56 g.g_y\[3\].g_x\[3\].t.r_d _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2558_ g.bi_l\[47\]\[0\] _1787_ _0209_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2489_ _0155_ _0158_ _0135_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2832__I _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3211__A1 _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3514__A2 _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1911__I g.g_y\[0\].g_x\[6\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1860_ g.bi_l\[48\]\[0\] g.g_y\[6\].g_x\[0\].t.r_h _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_44_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3461_ net34 _1039_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3530_ _1117_ _1124_ g.g_y\[0\].g_x\[2\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 in[4] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2343_ _1535_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2274_ _1438_ _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3392_ _0982_ _0813_ _0816_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2412_ g.bi_l\[34\]\[1\] net66 g.g_y\[4\].g_x\[2\].t.r_d _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4013_ g.g_y\[1\].g_x\[2\].t.out_sc _4013_/E g.g_y\[1\].g_x\[2\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_47_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1989_ _1456_ _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3744__A2 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3728_ _1085_ _1077_ _1101_ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3659_ _0832_ _0657_ _0663_ _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2171__A1 _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3671__A1 _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1843_ _1337_ _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1912_ g.bi_l\[6\]\[1\] net33 g.g_y\[0\].g_x\[6\].t.r_d _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2961_ g.g_y\[2\].g_x\[7\].t.out_sc _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2892_ _0536_ _0346_ _0355_ _0333_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3513_ _1107_ _1108_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3444_ _0953_ _0955_ _0958_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2326_ _1512_ _1515_ g.g_y\[6\].g_x\[5\].t.r_h _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2257_ _1702_ _1731_ _1378_ _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3375_ _0976_ _0981_ _0986_ _0989_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2217__A2 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2188_ g.g_y\[0\].g_x\[1\].t.r_d _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3717__A2 _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3427__B _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2153__A1 _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3008__I1 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2042_ g.bi_l\[52\]\[0\] g.g_y\[6\].g_x\[4\].t.r_v _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2111_ g.g_y\[0\].g_x\[3\].t.r_v _1595_ _1598_ _1599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3160_ _0390_ _0413_ _0786_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3091_ _0685_ _0712_ _0453_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2695__A2 _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3993_ g.g_y\[1\].g_x\[6\].t.out_sc _3993_/E g.g_y\[1\].g_x\[6\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1826_ net27 g.bi_l\[0\]\[1\] _1320_ _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2944_ g.bi_l\[15\]\[0\] _0585_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2875_ _0518_ _0521_ g.g_y\[3\].g_x\[2\].t.r_v _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3358_ _0777_ _0605_ _0973_ _1307_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3427_ _1019_ _1021_ _1023_ _0928_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_68_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2309_ _1786_ _1787_ _1788_ _1789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_0_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3289_ _0891_ _0897_ _0907_ _0909_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA_input10_I in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2749__I0 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout128_I net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2660_ _0107_ _0092_ _0100_ _0320_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_26_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2591_ _0231_ _0240_ _0254_ _0233_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3212_ g.g_y\[3\].g_x\[4\].t.r_v _0465_ _0468_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_1_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2025_ _1489_ _1512_ _1515_ _1516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3074_ g.g_y\[2\].g_x\[3\].t.r_d _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input2_I in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3143_ _1745_ _0771_ _0772_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2927_ _0142_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_28_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3976_ g.g_y\[2\].g_x\[1\].t.w_si net122 g.g_y\[2\].g_x\[1\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2840__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3093__A2 _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1809_ g.bi_l\[63\]\[1\] net108 _1303_ _1304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2356__A1 _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2789_ g.g_y\[5\].g_x\[4\].t.r_v _0047_ _0438_ g.g_y\[4\].g_x\[4\].t.r_v _0439_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_25_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2858_ _0501_ _0503_ _0504_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_37_Left_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2131__I1 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3440__B _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2347__A1 _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4022__CLK net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3830_ g.g_y\[5\].g_x\[7\].t.w_na _3830_/E _3830_/RN g.bi_l\[47\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3761_ net103 _3761_/E g.g_y\[7\].g_x\[4\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XANTENNA__2122__I1 _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2822__A2 _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2712_ _0332_ _0363_ _0369_ g.g_y\[5\].g_x\[1\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2574_ _0234_ _0236_ _0237_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2643_ _0286_ _0303_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3692_ _0752_ _0756_ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2008_ g.g_y\[6\].g_x\[4\].t.r_h _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_3126_ _0733_ _0749_ _0757_ g.g_y\[3\].g_x\[1\].t.r_v _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3057_ _0287_ _0288_ _0691_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_45_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3959_ net50 _3959_/E g.g_y\[2\].g_x\[4\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_9_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2290_ g.g_y\[5\].g_x\[6\].t.r_v _1770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3813_ g.g_y\[6\].g_x\[2\].t.w_dh _3813_/E _3813_/RN g.bi_l\[50\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3744_ _1132_ _1134_ _1294_ _1296_ g.g_y\[0\].g_x\[0\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2557_ _0167_ _0221_ _0222_ _0223_ g.g_y\[5\].g_x\[7\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3675_ _0820_ _0822_ _0823_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2626_ g.g_y\[3\].g_x\[3\].t.r_v _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2488_ _0134_ _0145_ _0156_ _0157_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_38_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3109_ g.bi_l\[16\]\[0\] g.g_y\[2\].g_x\[0\].t.r_h _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2798__A1 _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3039__A2 _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput13 in[5] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3460_ _1061_ _1062_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3391_ _1000_ _1002_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout110_I net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2411_ _0083_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2273_ _1753_ _1754_ _1755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2342_ _1751_ _0017_ _0018_ g.g_y\[6\].g_x\[5\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4012_ g.g_y\[1\].g_x\[2\].t.w_si net122 g.g_y\[1\].g_x\[2\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1988_ _1455_ _1466_ _1476_ _1478_ _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3727_ _0019_ _0021_ _1093_ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3589_ _0002_ _0004_ _0005_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2704__A1 _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2609_ _0230_ _0260_ _1492_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3658_ _0198_ _1222_ _1224_ _1225_ g.g_y\[3\].g_x\[7\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2960_ _0595_ _0600_ _0601_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3671__A2 _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1842_ g.g_y\[6\].g_x\[7\].t.r_v _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_1911_ g.g_y\[0\].g_x\[6\].t.r_v _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2891_ _0347_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3512_ _1578_ _1577_ _1594_ _1597_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3374_ _0970_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3443_ _1027_ _1029_ _1048_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2325_ _1514_ _1498_ _1506_ _0003_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2187_ _1672_ g.g_y\[7\].g_x\[2\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2256_ _1734_ _1736_ _1738_ _1732_ _1740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3662__A2 _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2153__A2 _1639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2392__A2 _1743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2041_ g.bi_l\[52\]\[1\] net90 _1531_ _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2110_ _1588_ _1587_ _1596_ _1597_ _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3090_ _1756_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2943_ g.g_y\[1\].g_x\[7\].t.r_v _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3992_ g.g_y\[1\].g_x\[6\].t.w_si net124 g.g_y\[1\].g_x\[6\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1825_ g.g_y\[0\].g_x\[0\].t.r_d _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2874_ _0512_ _0511_ _0519_ _0520_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_13_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2308_ g.bi_l\[47\]\[0\] g.g_y\[5\].g_x\[7\].t.r_h _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_fanout90_I net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3357_ _0607_ _0610_ _0583_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_13_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3426_ _0848_ _1026_ _1031_ _1033_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_68_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3796__CLK net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2239_ _1703_ _1712_ _1723_ _1705_ _1724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_0_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3288_ _0891_ _0908_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2071__A1 _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1949__A2 _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2590_ _0253_ _0236_ _0237_ _0231_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_22_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3562__A1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3211_ _0774_ _0834_ _0835_ g.g_y\[2\].g_x\[5\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3142_ _0616_ _0548_ _0564_ _0567_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_65_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2024_ _1505_ _1504_ _1513_ _1514_ _1515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3073_ _0694_ _0696_ _0697_ _0701_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2857_ g.g_y\[3\].g_x\[2\].t.r_v _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3975_ g.g_y\[2\].g_x\[1\].t.out_sc _3975_/E g.g_y\[2\].g_x\[1\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_9_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2926_ _0545_ _0562_ _0569_ _0556_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1808_ g.g_y\[7\].g_x\[7\].t.r_d _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2356__A2 _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2788_ g.g_y\[5\].g_x\[4\].t.r_v _0049_ _0052_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3409_ _0993_ _1017_ _1018_ g.g_y\[1\].g_x\[4\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2347__A2 _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3544__A1 _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3760_ g.g_y\[7\].g_x\[5\].t.w_na _3760_/E _3760_/RN g.bi_l\[61\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2711_ _0364_ _0366_ _0368_ _0332_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2573_ g.bi_l\[29\]\[0\] g.g_y\[3\].g_x\[5\].t.r_v _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3691_ g.g_y\[3\].g_x\[0\].t.r_v _0562_ _0935_ _0946_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2642_ net68 _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3125_ _0752_ _0756_ g.g_y\[2\].g_x\[1\].t.r_v _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2007_ _1495_ _1497_ _1488_ _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3056_ g.bi_l\[27\]\[0\] g.g_y\[3\].g_x\[3\].t.r_v _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2026__A1 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3958_ g.g_y\[2\].g_x\[5\].t.out_sc _3958_/E g.g_y\[2\].g_x\[5\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3889_ net66 _3889_/E g.g_y\[4\].g_x\[2\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_18_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2909_ g.bi_l\[16\]\[1\] net44 _0552_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__A2 _1743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1863__I1 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_56_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3812_ net87 _3812_/E g.g_y\[6\].g_x\[2\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_42_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3743_ _1389_ _1295_ _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3674_ _1235_ _1238_ g.g_y\[3\].g_x\[1\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2556_ net82 _1743_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2487_ g.g_y\[5\].g_x\[0\].t.r_d _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ g.g_y\[4\].g_x\[3\].t.r_d _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_10_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3108_ _0736_ _0738_ _0739_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3039_ _0637_ _0664_ _0235_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4012__CLK net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2722__A2 _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2789__A2 _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3738__A1 _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 in[6] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2341_ net91 _1757_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3390_ _0832_ _0657_ _1001_ _1461_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2410_ g.g_y\[4\].g_x\[2\].t.r_v _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2272_ _1338_ _1346_ _1363_ _1367_ _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4011_ g.g_y\[1\].g_x\[2\].t.out_sc _4011_/E g.g_y\[1\].g_x\[2\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3726_ _1406_ _1277_ _1280_ _1281_ g.g_y\[0\].g_x\[6\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1987_ _1477_ _1455_ _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3657_ g.g_y\[4\].g_x\[7\].t.r_v _0197_ _0580_ _0198_ _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_7_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2539_ _1341_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2608_ _0262_ _0271_ g.g_y\[5\].g_x\[5\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2704__A2 _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3588_ _1676_ _1165_ _1167_ _1168_ g.g_y\[7\].g_x\[1\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_2_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1910_ g.g_y\[7\].g_x\[6\].t.r_d _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_60_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2890_ _0349_ _0532_ _0534_ _0535_ g.g_y\[4\].g_x\[2\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_71_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1841_ _1299_ _1329_ _1335_ g.g_y\[7\].g_x\[7\].t.r_v _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_52_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3511_ _1106_ _1587_ _1596_ _1568_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2324_ _1514_ _1507_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3373_ _1564_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3442_ _1027_ _0912_ _0915_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2186_ net97 _1671_ _1565_ _1672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2255_ _1733_ _1739_ g.g_y\[7\].g_x\[1\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2870__A1 _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3709_ _0880_ _0705_ _1022_ _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2613__A1 _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2040_ g.g_y\[6\].g_x\[4\].t.r_d _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3991_ g.g_y\[1\].g_x\[6\].t.out_sc _3991_/E g.g_y\[1\].g_x\[6\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_2942_ g.g_y\[2\].g_x\[7\].t.r_d _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2873_ g.g_y\[3\].g_x\[2\].t.r_d _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_17_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1824_ g.g_y\[0\].g_x\[0\].t.r_h _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_13_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2307_ net83 g.bi_l\[47\]\[1\] g.g_y\[5\].g_x\[7\].t.r_d _1787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3356_ _1299_ _1329_ _0971_ _0585_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_2238_ _1706_ _1708_ _1709_ _1703_ _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3287_ g.g_y\[1\].g_x\[2\].t.out_sc _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3425_ _1019_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_68_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2169_ g.g_y\[7\].g_x\[2\].t.r_v _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_48_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3890__CLK net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3562__A2 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3210_ net49 _0682_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3141_ _0545_ _0555_ _0566_ _0546_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_65_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2023_ g.g_y\[6\].g_x\[5\].t.r_d _1514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3072_ _0686_ _0692_ _0706_ _0688_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_15_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1807_ _1301_ _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ g.g_y\[2\].g_x\[2\].t.w_na _3974_/E _3974_/RN g.bi_l\[18\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2925_ _0565_ _0568_ _0545_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2856_ _0083_ _0085_ _0502_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2787_ _0277_ _0436_ _0437_ g.g_y\[4\].g_x\[5\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3408_ net39 _0883_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3339_ g.g_y\[1\].g_x\[0\].t.r_d _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3544__A2 _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout133_I net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2710_ _0210_ _0212_ _0367_ _0364_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3690_ _0938_ _0952_ _0959_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3786__CLK net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2572_ g.bi_l\[29\]\[1\] net59 _0235_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2641_ _0298_ _0300_ _0301_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3124_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3055_ _1573_ _1574_ _0689_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2026__A2 _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2006_ _1456_ _1458_ _1496_ _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_26_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3957_ g.g_y\[2\].g_x\[5\].t.out_sc _3957_/E g.g_y\[2\].g_x\[5\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_60_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2839_ _0486_ _0300_ _0309_ _0286_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2908_ g.g_y\[2\].g_x\[0\].t.r_d _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3888_ net68 _3888_/E g.g_y\[4\].g_x\[3\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XANTENNA__3462__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2265__A2 _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3811_ net87 _3811_/E g.g_y\[6\].g_x\[2\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_59_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3742_ _0129_ _0131_ _1135_ _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2624_ _0284_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3673_ _1236_ _1237_ _0335_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2555_ _0209_ _0214_ _0219_ _0207_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2486_ _1384_ _1386_ _0147_ _0134_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_38_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3038_ _0666_ _0675_ g.g_y\[3\].g_x\[5\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3107_ g.g_y\[2\].g_x\[1\].t.r_v _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_65_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput15 in[7] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2271_ _1752_ _1356_ _1366_ _1339_ _1753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2340_ _0015_ _0016_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4010_ g.g_y\[1\].g_x\[3\].t.w_na _4010_/E _4010_/RN g.bi_l\[11\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_55_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1986_ g.g_y\[0\].g_x\[5\].t.out_sc _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_43_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2170__C _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3725_ _1069_ _1071_ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2607_ _0263_ _0265_ _0270_ _1492_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3587_ _0125_ _1722_ _1730_ _1676_ _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3656_ _0620_ _1223_ _0615_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2538_ _0174_ _0197_ _0205_ _1362_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2469_ net15 _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1903__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1840_ g.g_y\[0\].g_x\[7\].t.r_v _1331_ _1334_ _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_25_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3510_ _1588_ _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3441_ _1043_ _1046_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2323_ g.g_y\[6\].g_x\[5\].t.r_h _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2254_ _1734_ _1736_ _1738_ _1378_ _1739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3372_ _0970_ _0975_ _0987_ g.g_y\[1\].g_x\[7\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4002__CLK net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2185_ _1669_ _1670_ _1671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2870__A2 _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2622__A2 _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1969_ _1456_ _1458_ _1459_ _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3639_ _0475_ _1209_ _0473_ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3708_ _0641_ _1262_ _1264_ _1266_ g.g_y\[1\].g_x\[5\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_54_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3629__A1 _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3990_ g.g_y\[1\].g_x\[7\].t.w_na _3990_/E _3990_/RN g.bi_l\[15\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_72_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1823_ _1313_ _1315_ _1317_ _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2941_ _0582_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2872_ _0506_ _0507_ _0508_ _0512_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_40_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2915__I0 _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3424_ _1019_ _1024_ _1032_ g.g_y\[1\].g_x\[3\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2306_ g.g_y\[5\].g_x\[7\].t.r_h _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3355_ _1331_ _1334_ g.g_y\[0\].g_x\[7\].t.r_v _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2237_ _1705_ _1713_ _1719_ _1721_ _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3286_ _0903_ _0905_ _0906_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2168_ _1637_ _1648_ _1653_ _1655_ _1656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_45_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2099_ _1467_ _1469_ _1586_ _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_0_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_59_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2531__A1 _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3331__I0 _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3140_ _0560_ _0532_ _0769_ _0770_ g.g_y\[3\].g_x\[1\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3071_ _1573_ _1574_ _0689_ _0686_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2022_ _1499_ _1500_ _1501_ _1505_ _1513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3973_ g.g_y\[2\].g_x\[2\].t.w_dh _3973_/E _3973_/RN g.bi_l\[18\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_1806_ g.g_y\[7\].g_x\[7\].t.r_v _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_2786_ net70 _0380_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2855_ g.bi_l\[34\]\[0\] g.g_y\[4\].g_x\[2\].t.r_v _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_13_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2924_ _0544_ _0555_ _0566_ _0567_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2761__A1 _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3338_ _0551_ _0553_ _0947_ _0937_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_3407_ _1015_ _1016_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3269_ g.g_y\[1\].g_x\[2\].t.r_v _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_62_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2640_ g.g_y\[4\].g_x\[3\].t.r_h _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA_fanout126_I net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2571_ g.g_y\[3\].g_x\[5\].t.r_d _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2743__A1 _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2005_ g.bi_l\[61\]\[0\] g.g_y\[7\].g_x\[5\].t.r_v _1496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3123_ _0745_ _0744_ _0753_ _0754_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3054_ g.bi_l\[11\]\[0\] g.g_y\[1\].g_x\[3\].t.r_v _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3956_ g.g_y\[2\].g_x\[5\].t.w_si net124 g.g_y\[2\].g_x\[5\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2907_ g.g_y\[2\].g_x\[0\].t.r_v _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2769_ g.g_y\[4\].g_x\[5\].t.r_h _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2838_ _0301_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3887_ net68 _3887_/E g.g_y\[4\].g_x\[3\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_13_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3880__CLK net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3810_ g.g_y\[6\].g_x\[2\].t.w_si net116 g.g_y\[6\].g_x\[2\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3741_ _1322_ _1139_ _1292_ _1293_ _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3453__A2 _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3205__A2 _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2554_ _0172_ _0206_ _1341_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_30_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2623_ g.g_y\[4\].g_x\[3\].t.r_v _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_6_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3672_ _0538_ _0351_ _0759_ _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2449__B _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2485_ _0153_ _0138_ _0154_ _0136_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__2184__B _1658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3037_ _0667_ _0669_ _0674_ _0235_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3106_ _0335_ _0336_ _0737_ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_21_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3939_ g.g_y\[3\].g_x\[1\].t.w_dh _3939_/E _3939_/RN g.bi_l\[25\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_14_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3776__CLK net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 in[8] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2270_ _1357_ _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3724_ _1278_ _1279_ _1316_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1985_ _1472_ _1474_ _1475_ _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_43_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2937__A1 _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2606_ _0266_ _0268_ _0269_ _0263_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3586_ _1736_ _1166_ _1734_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2537_ _0174_ _0200_ _0204_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3655_ _0621_ _0623_ _0624_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2399_ net88 _0072_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2468_ _0093_ _0094_ _0137_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2960__I1 _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3353__A1 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3408__A2 _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1947__I _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2395__A2 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3371_ _0976_ _0981_ _0986_ _0970_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3440_ _1044_ _1695_ _1045_ _1680_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_4_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2322_ _1413_ _0000_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2184_ _1657_ _1641_ _1658_ _1637_ _1670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2253_ _1375_ _1397_ _1737_ _1734_ _1738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_20_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3647__A2 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1968_ g.bi_l\[61\]\[0\] g.g_y\[7\].g_x\[5\].t.r_v _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1899_ _1388_ _1392_ _1393_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3707_ _1265_ _1005_ _0798_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3569_ _1338_ _1361_ _1369_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3638_ g.g_y\[4\].g_x\[3\].t.r_h _0477_ _0478_ _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3574__A1 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__A2 _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2940_ g.g_y\[2\].g_x\[7\].t.r_v _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_29_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1822_ g.bi_l\[6\]\[0\] _1316_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2871_ _0504_ _0503_ _0517_ _0496_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_13_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3354_ g.g_y\[1\].g_x\[7\].t.r_d _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3423_ _0848_ _1026_ _1031_ _1019_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_68_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2305_ _1782_ _1783_ _1784_ _1785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2236_ _1705_ _1720_ _1721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2167_ _1654_ net98 _1655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_29_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3285_ g.g_y\[1\].g_x\[2\].t.r_h _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2098_ g.bi_l\[4\]\[0\] _1470_ _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_0_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2021_ _1488_ _1497_ _1511_ _1490_ _1512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3070_ _0688_ _0693_ _0702_ _0704_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3972_ net46 _3972_/E g.g_y\[2\].g_x\[2\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2923_ g.g_y\[3\].g_x\[0\].t.r_d _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1805_ g.g_y\[0\].g_x\[7\].t.r_d _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2785_ _0434_ _0435_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2854_ _0498_ _0499_ _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2761__A2 _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3406_ _0839_ _0844_ _0858_ _0861_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3710__A1 _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3337_ _0953_ _0941_ _0954_ _0939_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_68_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2219_ _1703_ _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3199_ _0775_ _0783_ _0825_ _0592_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3268_ g.g_y\[2\].g_x\[2\].t.r_v _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2504__A2 _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2268__A1 _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout119_I net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2570_ g.g_y\[3\].g_x\[5\].t.r_v _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__2743__A2 _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3122_ g.g_y\[2\].g_x\[1\].t.r_d _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_10_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ _1491_ _1493_ _1494_ _1495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3053_ g.g_y\[2\].g_x\[3\].t.r_d _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2431__A1 _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3955_ g.g_y\[2\].g_x\[5\].t.out_sc _3955_/E g.g_y\[2\].g_x\[5\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3886_ g.g_y\[4\].g_x\[3\].t.w_si net112 g.g_y\[4\].g_x\[3\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2906_ _0548_ _0549_ g.g_y\[3\].g_x\[0\].t.r_h _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2768_ _1775_ _0420_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2837_ _0276_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2699_ _0347_ _0346_ _0355_ _0356_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_67_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3740_ _1322_ net10 _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2553_ _0208_ _0220_ g.g_y\[5\].g_x\[7\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2622_ g.g_y\[6\].g_x\[3\].t.r_v _1622_ _0282_ g.g_y\[5\].g_x\[3\].t.r_v _0283_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_50_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_34_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_30_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ _0733_ _0749_ _0757_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2716__A2 _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2484_ net15 g.g_y\[5\].g_x\[0\].t.r_h _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3105_ g.bi_l\[25\]\[0\] g.g_y\[3\].g_x\[1\].t.r_v _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3141__A2 _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2652__A1 _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Left_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3036_ _0670_ _0672_ _0673_ _0667_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2007__I1 _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3869_ net71 _3869_/E g.g_y\[4\].g_x\[6\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XTAP_TAPCELL_ROW_21_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3938_ net53 _3938_/E g.g_y\[3\].g_x\[1\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XPHY_EDGE_ROW_52_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_72_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 in[9] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_70_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3371__A2 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3723_ g.g_y\[0\].g_x\[5\].t.r_h _1077_ _1078_ _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1984_ g.g_y\[0\].g_x\[5\].t.r_h _1475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_43_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3654_ _0777_ _0605_ _0611_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3870__CLK net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3585_ _1375_ _1397_ _1737_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2605_ _0049_ _0052_ g.g_y\[5\].g_x\[4\].t.r_h _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2467_ g.bi_l\[41\]\[0\] g.g_y\[5\].g_x\[1\].t.r_h _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2536_ _0193_ _0192_ _0202_ _0203_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_2_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2398_ _1756_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2228__I1 _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3019_ _0640_ _0646_ _0654_ _0656_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_61_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2321_ _1770_ _1794_ _1800_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3370_ _0982_ _0984_ _0985_ _0976_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2183_ _1660_ _1650_ _1661_ _1654_ _1669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2252_ _1374_ _1399_ _1401_ _1737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2743__B _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3574__B _1516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ g.bi_l\[61\]\[1\] net104 _1457_ _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1898_ g.g_y\[7\].g_x\[0\].t.r_v _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3706_ _1006_ _1008_ _1009_ _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3637_ _0441_ _0463_ _0469_ _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3499_ _1590_ _1597_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2519_ _0184_ _0185_ _0186_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3568_ _1145_ _1152_ _3568_/ZN vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3574__A2 _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3484__B _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3915__D net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2870_ _0498_ _0499_ _0500_ _0504_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1821_ g.g_y\[0\].g_x\[6\].t.r_h _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2304_ g.bi_l\[45\]\[0\] g.g_y\[5\].g_x\[5\].t.r_h _1784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3353_ _0724_ _0967_ _0968_ _0969_ g.g_y\[2\].g_x\[0\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3284_ _0846_ _0847_ _0904_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3422_ _1027_ _1029_ _1030_ _0848_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2166_ g.g_y\[7\].g_x\[2\].t.r_d _1654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2235_ g.g_y\[6\].g_x\[1\].t.out_sc _1720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2097_ _1580_ _1582_ _1584_ _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2999_ g.g_y\[4\].g_x\[5\].t.r_v _0252_ _0636_ g.g_y\[3\].g_x\[5\].t.r_v _0637_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2020_ _1510_ _1493_ _1494_ _1488_ _1511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_72_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ net47 _3971_/E g.g_y\[2\].g_x\[2\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_2853_ g.bi_l\[18\]\[0\] g.g_y\[2\].g_x\[2\].t.r_v _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_15_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2922_ _0141_ _0143_ _0557_ _0544_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_17_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1804_ g.g_y\[0\].g_x\[7\].t.r_v _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3538__A2 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2784_ _0232_ _0240_ _0254_ _0257_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_31_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3267_ _0498_ _0887_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3710__A2 _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3336_ net11 g.g_y\[1\].g_x\[0\].t.r_h _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3405_ _0853_ _0852_ _0860_ _0840_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_72_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2149_ g.g_y\[7\].g_x\[2\].t.r_d _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2218_ g.g_y\[6\].g_x\[1\].t.r_v _1703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3198_ _0607_ _0610_ _0775_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2268__A2 _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3121_ _0596_ _0598_ _0741_ _0745_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2003_ g.bi_l\[45\]\[0\] g.g_y\[5\].g_x\[5\].t.r_v _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3456__A1 _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3052_ _0686_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2431__A2 _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ g.g_y\[2\].g_x\[6\].t.w_na _3954_/E _3954_/RN g.bi_l\[22\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2836_ _0481_ _0482_ _0483_ _0484_ g.g_y\[4\].g_x\[4\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3885_ g.g_y\[4\].g_x\[3\].t.out_sc _3885_/E g.g_y\[4\].g_x\[3\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_2905_ net13 _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2767_ _0390_ _0413_ _0419_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2698_ g.g_y\[4\].g_x\[1\].t.r_d _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3319_ g.g_y\[1\].g_x\[0\].t.r_v _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_64_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout131_I net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3670_ _0764_ _1234_ _0762_ _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2552_ _0209_ _0214_ _0219_ _1341_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2621_ g.g_y\[6\].g_x\[3\].t.r_v _1625_ _1628_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2483_ g.g_y\[5\].g_x\[0\].t.r_h _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3035_ _0465_ _0468_ g.g_y\[3\].g_x\[4\].t.r_h _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3104_ _1680_ _1681_ _0735_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2652__A2 _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3937_ net53 _3937_/E g.g_y\[3\].g_x\[1\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3799_ net90 _3799_/E g.g_y\[6\].g_x\[4\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_61_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3868_ g.g_y\[4\].g_x\[7\].t.out_sc _3868_/E g.g_y\[4\].g_x\[7\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_2819_ _0441_ _0465_ _0468_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_21_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3668__A1 _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1983_ _1313_ _1315_ _1473_ _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2604_ _0051_ _0035_ _0044_ _0267_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_3722_ _1060_ _1067_ _1080_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3653_ _0556_ _1216_ _1217_ _1221_ g.g_y\[4\].g_x\[0\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_21_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3584_ g.g_y\[0\].g_x\[1\].t.r_v _1695_ _1701_ _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2535_ g.g_y\[4\].g_x\[7\].t.r_d _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2466_ g.g_y\[5\].g_x\[0\].t.r_d _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2397_ _0069_ _0070_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3018_ _0640_ _0655_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3050__A2 _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2386__B g.g_y\[6\].g_x\[3\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3041__A2 _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2320_ _1796_ _1799_ g.g_y\[5\].g_x\[6\].t.r_v _1800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2251_ _1636_ _1656_ _1735_ _1736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2182_ _1557_ _1666_ _1667_ _1668_ g.g_y\[7\].g_x\[3\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_48_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1966_ g.g_y\[7\].g_x\[5\].t.r_d _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1897_ _1389_ _1390_ _1391_ _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3636_ _0201_ _1204_ _1206_ _1207_ g.g_y\[4\].g_x\[6\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3567_ _1151_ net4 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3705_ _0999_ _1263_ _0641_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2449_ _0074_ _0115_ _0117_ _0013_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3498_ _1090_ _1092_ _1094_ _1095_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2518_ g.bi_l\[38\]\[0\] g.g_y\[4\].g_x\[6\].t.r_h _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_3_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1820_ net33 g.bi_l\[6\]\[1\] _1314_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3262__A2 _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3421_ _0912_ _0915_ g.g_y\[1\].g_x\[2\].t.r_h _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2303_ net80 g.bi_l\[45\]\[1\] g.g_y\[5\].g_x\[5\].t.r_d _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2234_ _1715_ _1717_ _1718_ _1719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3352_ net43 _1747_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3283_ g.bi_l\[11\]\[0\] g.g_y\[1\].g_x\[3\].t.r_h _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2165_ _1650_ _1652_ g.g_y\[7\].g_x\[2\].t.r_h _1653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2096_ g.bi_l\[2\]\[0\] _1583_ _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_0_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1949_ _1373_ _1403_ _1436_ _1371_ _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_61_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2998_ g.g_y\[4\].g_x\[5\].t.r_v _0255_ _0258_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_16_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3619_ g.g_y\[6\].g_x\[5\].t.r_v _1509_ _0229_ _1510_ _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_31_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3483__A2 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3970_ g.g_y\[2\].g_x\[2\].t.w_si net122 g.g_y\[2\].g_x\[2\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3235__A2 _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3756__CLK net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1803_ _1298_ _1803_/Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2783_ _0248_ _0247_ _0256_ _0233_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_31_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2852_ g.bi_l\[18\]\[1\] net46 g.g_y\[2\].g_x\[2\].t.r_d _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2921_ _0563_ _0548_ _0564_ _0546_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_53_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3404_ _0855_ _0988_ _1013_ _1014_ g.g_y\[1\].g_x\[5\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_0_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3474__A2 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2217_ g.g_y\[0\].g_x\[1\].t.r_v _1695_ _1701_ _1676_ _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3197_ _0820_ _0822_ _0823_ g.g_y\[2\].g_x\[6\].t.r_h _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3266_ _0495_ _0516_ _0886_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3335_ g.g_y\[1\].g_x\[0\].t.r_h _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_64_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2148_ g.g_y\[7\].g_x\[2\].t.r_h _1636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2079_ g.g_y\[0\].g_x\[3\].t.r_v _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3456__A2 _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3120_ _0751_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3051_ g.g_y\[2\].g_x\[3\].t.r_v _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2002_ g.bi_l\[45\]\[1\] net80 _1492_ _1493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3953_ g.g_y\[2\].g_x\[6\].t.w_dh _3953_/E _3953_/RN g.bi_l\[22\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__3208__A2 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2766_ _0415_ _0418_ g.g_y\[3\].g_x\[6\].t.r_v _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3884_ g.g_y\[4\].g_x\[4\].t.w_na _3884_/E _3884_/RN g.bi_l\[36\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2835_ net68 _0274_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2719__A1 _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2904_ _0506_ _0507_ _0547_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__1942__A2 _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2697_ _0188_ _0190_ _0343_ _0347_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__3144__A1 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3318_ g.g_y\[3\].g_x\[0\].t.r_v _0562_ _0935_ g.g_y\[2\].g_x\[0\].t.r_v _0936_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_68_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3249_ g.g_y\[2\].g_x\[3\].t.r_h _0871_ _0872_ _0867_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_24_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2620_ _0277_ _0280_ _0281_ g.g_y\[5\].g_x\[4\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3667__C _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout124_I net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2551_ _0215_ _0217_ _0218_ g.g_y\[5\].g_x\[7\].t.r_h _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2482_ _0136_ _0140_ _0149_ _0151_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__3126__A1 _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3103_ g.bi_l\[9\]\[0\] g.g_y\[1\].g_x\[1\].t.r_v _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3034_ _0467_ _0451_ _0460_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_58_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3936_ g.g_y\[3\].g_x\[1\].t.w_si net111 g.g_y\[3\].g_x\[1\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3798_ g.g_y\[6\].g_x\[5\].t.out_sc _3798_/E g.g_y\[6\].g_x\[5\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_3867_ g.g_y\[4\].g_x\[7\].t.out_sc _3867_/E g.g_y\[4\].g_x\[7\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2749_ net59 g.bi_l\[29\]\[1\] g.g_y\[3\].g_x\[5\].t.r_d _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2818_ _0459_ _0458_ _0466_ _0467_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__3668__A2 _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1906__A2 _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3595__A1 g.g_y\[6\].g_x\[3\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1982_ g.bi_l\[6\]\[0\] _1316_ _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_35_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3721_ _1764_ _1766_ _1072_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2603_ _0051_ _0045_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3583_ _1593_ _1161_ _1163_ _1164_ g.g_y\[7\].g_x\[3\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2534_ _0201_ _0185_ _0186_ _0193_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3652_ _0573_ _1219_ _1220_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2396_ _1602_ _1609_ _1624_ _1627_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2465_ _0134_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1833__A1 _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1887__I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3017_ g.g_y\[2\].g_x\[5\].t.out_sc _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3919_ g.g_y\[3\].g_x\[5\].t.w_dh _3919_/E _3919_/RN g.bi_l\[29\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_6_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3754__D net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2313__A2 _1792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout130 net131 net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3577__A1 _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2552__A2 _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2250_ _1636_ _1659_ _1662_ _1735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2181_ net99 _1445_ _1668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2091__I1 _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1965_ g.g_y\[7\].g_x\[5\].t.r_v _1456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3704_ _1454_ _1479_ _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_59_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1896_ g.bi_l\[0\]\[0\] g.g_y\[0\].g_x\[0\].t.r_v _1391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3635_ _0420_ _0388_ _1773_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2517_ net71 g.bi_l\[38\]\[1\] g.g_y\[4\].g_x\[6\].t.r_d _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3497_ _1468_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3566_ _1151_ net4 _1145_ _3566_/ZN vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2379_ _1531_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2448_ _1645_ _0079_ _0119_ g.g_y\[6\].g_x\[2\].t.r_d _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input17_I in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4049_ net30 _4049_/E g.g_y\[0\].g_x\[2\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_3_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_49_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2782__A2 _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_67_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3691__B _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3351_ _0936_ _0960_ _0552_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3420_ _0914_ _0897_ _0907_ _1028_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2302_ g.g_y\[5\].g_x\[5\].t.r_h _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_2233_ g.g_y\[6\].g_x\[1\].t.r_h _1718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2164_ _1377_ _1379_ _1651_ _1652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input9_I in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3282_ _0899_ _0900_ _0902_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2095_ g.g_y\[0\].g_x\[2\].t.r_h _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1948_ _1336_ _1370_ _1303_ _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1879_ g.g_y\[7\].g_x\[0\].t.r_h _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2997_ _0485_ _0634_ _0635_ g.g_y\[3\].g_x\[6\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3618_ _0265_ _1192_ _0263_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3549_ _1686_ net10 _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_8_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3704__A1 _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2920_ net13 g.g_y\[3\].g_x\[0\].t.r_h _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_15_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2782_ _0250_ _0010_ _0431_ _0433_ g.g_y\[4\].g_x\[6\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1802_ net8 net7 _1297_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2851_ _0497_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_13_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3403_ _0998_ _1000_ _1002_ _0928_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3334_ _0939_ _0943_ _0949_ _0951_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2147_ _1523_ _1547_ _1634_ _1635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2216_ g.g_y\[0\].g_x\[1\].t.r_v _1697_ _1700_ _1701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3196_ _0659_ _0662_ g.g_y\[2\].g_x\[5\].t.r_h _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3265_ _0495_ _0518_ _0521_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2078_ _1566_ g.g_y\[7\].g_x\[4\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2673__A1 _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2200__I1 _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2077__S _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2001_ g.g_y\[5\].g_x\[5\].t.r_d _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3050_ g.g_y\[4\].g_x\[3\].t.r_v _0305_ _0684_ g.g_y\[3\].g_x\[3\].t.r_v _0685_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_61_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3952_ net51 _3952_/E g.g_y\[2\].g_x\[6\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3883_ g.g_y\[4\].g_x\[4\].t.w_dh _3883_/E _3883_/RN g.bi_l\[36\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2903_ g.bi_l\[25\]\[0\] g.g_y\[3\].g_x\[1\].t.r_h _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2834_ _0473_ _0475_ _0479_ _0471_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2696_ _0353_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2765_ _0409_ _0408_ _0416_ _0417_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_5_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3144__A2 _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3317_ _0565_ _0568_ g.g_y\[3\].g_x\[0\].t.r_v _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3179_ _0803_ _0804_ _0805_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3248_ _0707_ _0710_ g.g_y\[2\].g_x\[3\].t.r_h _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2646__A1 _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2550_ _1796_ _1799_ g.g_y\[5\].g_x\[6\].t.r_h _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_fanout117_I net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3683__C _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2481_ _0136_ _0150_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3126__A2 _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3102_ g.g_y\[2\].g_x\[1\].t.r_d _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3033_ _0467_ _0461_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3204__B _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3866_ g.g_y\[4\].g_x\[7\].t.w_si net117 g.g_y\[4\].g_x\[7\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3935_ net54 _3935_/E g.g_y\[3\].g_x\[1\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3797_ g.g_y\[6\].g_x\[5\].t.out_sc _3797_/E g.g_y\[6\].g_x\[5\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_26_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2748_ g.g_y\[3\].g_x\[5\].t.r_h _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_2817_ g.g_y\[3\].g_x\[4\].t.r_d _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2679_ g.bi_l\[25\]\[0\] g.g_y\[3\].g_x\[1\].t.r_v _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_14_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3595__A2 _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1981_ _1467_ _1469_ _1471_ _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3720_ _1272_ _1273_ _1276_ g.g_y\[1\].g_x\[1\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2602_ g.g_y\[5\].g_x\[4\].t.r_h _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3582_ _1567_ _1592_ _1599_ _1593_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2533_ _0184_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3651_ _0573_ net14 _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2395_ _0068_ _1617_ _1626_ _1603_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_47_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2464_ g.g_y\[5\].g_x\[0\].t.r_v _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_64_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3016_ _0650_ _0652_ _0653_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3849_ g.g_y\[5\].g_x\[3\].t.w_dh _3849_/E _3849_/RN g.bi_l\[43\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3918_ net60 _3918_/E g.g_y\[3\].g_x\[5\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_6_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout131 net132 net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout120 net121 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3577__A2 _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2180_ _1633_ _1635_ _1664_ _1631_ _1667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_18_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ g.g_y\[0\].g_x\[5\].t.r_d _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3634_ _0427_ _1205_ _0201_ _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1895_ g.bi_l\[0\]\[1\] net27 g.g_y\[0\].g_x\[0\].t.r_d _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3703_ _0832_ _0657_ _1001_ _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2447_ _0081_ _0103_ _0109_ _1645_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3740__A2 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3496_ _0019_ _0021_ _1093_ _1090_ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2516_ g.g_y\[4\].g_x\[6\].t.r_h _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3565_ net5 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2059__A2 _1528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2378_ _0025_ _0047_ _0053_ _1530_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4048_ g.g_y\[0\].g_x\[3\].t.out_sc _4048_/E g.g_y\[0\].g_x\[3\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XTAP_TAPCELL_ROW_54_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3559__A2 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2301_ _1777_ _1779_ _1780_ _1781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3350_ _0963_ net12 _0965_ _0961_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2289__A2 _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2232_ _1611_ _1613_ _1716_ _1717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2163_ g.bi_l\[57\]\[0\] g.g_y\[7\].g_x\[1\].t.r_h _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3281_ g.bi_l\[9\]\[0\] _0901_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_51_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2094_ net29 g.bi_l\[2\]\[1\] _1581_ _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1878_ g.g_y\[7\].g_x\[7\].t.r_h _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3617_ _0266_ _0268_ _0269_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1947_ _1440_ _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2996_ net59 _0380_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3479_ _1331_ _1334_ _1060_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3548_ _1127_ _1119_ _1139_ _1686_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_8_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3704__A2 _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2850_ g.g_y\[2\].g_x\[2\].t.r_v _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_15_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2781_ _0386_ _0426_ _0428_ _0432_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1801_ net9 _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_13_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3402_ _0800_ _1005_ _1010_ _1012_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3333_ _0939_ _0950_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3264_ g.g_y\[2\].g_x\[2\].t.r_d _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2146_ _1523_ _1550_ _1553_ _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2077_ net101 _1563_ _1565_ _1566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2215_ _1691_ _1690_ _1698_ _1699_ _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3195_ _0661_ _0646_ _0654_ _0821_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_15_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2781__B _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2979_ g.g_y\[3\].g_x\[6\].t.r_h _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1936__A1 _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2000_ g.g_y\[5\].g_x\[5\].t.r_v _1491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_26_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3882_ net70 _3882_/E g.g_y\[4\].g_x\[4\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3951_ net52 _3951_/E g.g_y\[2\].g_x\[6\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_2833_ _0439_ _0470_ _0029_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2902_ g.g_y\[3\].g_x\[0\].t.r_d _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2764_ g.g_y\[3\].g_x\[6\].t.r_d _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2695_ _0341_ _0340_ _0352_ _0333_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_5_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3316_ _0774_ _0933_ _0934_ g.g_y\[2\].g_x\[1\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3247_ _0709_ _0693_ _0702_ _0870_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__2407__A2 _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2129_ _1499_ _1500_ _1616_ _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__2067__I _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3178_ g.bi_l\[15\]\[0\] g.g_y\[1\].g_x\[7\].t.r_h _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2894__A2 _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2480_ g.g_y\[5\].g_x\[0\].t.out_sc _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3101_ g.g_y\[2\].g_x\[1\].t.r_v _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_38_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3032_ g.g_y\[3\].g_x\[4\].t.r_h _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3796_ g.g_y\[6\].g_x\[5\].t.w_si net120 g.g_y\[6\].g_x\[5\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3865_ g.g_y\[4\].g_x\[7\].t.out_sc _3865_/E g.g_y\[4\].g_x\[7\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XFILLER_0_33_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2615__I _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3934_ net55 _3934_/E g.g_y\[3\].g_x\[2\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2816_ _0452_ _0454_ _0455_ _0459_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2747_ _0396_ _0398_ _0399_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2678_ g.bi_l\[25\]\[1\] net53 g.g_y\[3\].g_x\[1\].t.r_d _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_72_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2800__A2 _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2619__A2 _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1980_ g.bi_l\[4\]\[0\] _1470_ _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3650_ _1218_ _0526_ _0536_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3044__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2601_ _0215_ _0217_ _0264_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3581_ _1635_ _1162_ _1633_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2463_ _0129_ _0131_ _0132_ g.g_y\[6\].g_x\[0\].t.r_v _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2532_ _0173_ _0182_ _0199_ _0175_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_2_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2394_ _1618_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4064_ g.g_y\[0\].g_x\[0\].t.w_na _4064_/E _4064_/RN g.bi_l\[0\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3015_ g.g_y\[2\].g_x\[5\].t.r_h _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_3_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout42_I net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3848_ net78 _3848_/E g.g_y\[5\].g_x\[3\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3779_ g.g_y\[7\].g_x\[1\].t.w_dh _3779_/E _3779_/RN g.bi_l\[57\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3917_ net60 _3917_/E g.g_y\[3\].g_x\[5\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfanout132 net133 net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout121 net134 net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout110 net111 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3274__A2 _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2537__A1 _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1899__I0 _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1963_ g.g_y\[0\].g_x\[5\].t.r_v _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3633_ _0376_ _0384_ _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1894_ g.g_y\[0\].g_x\[0\].t.r_v _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_3702_ _0585_ _1257_ _1259_ _1261_ g.g_y\[1\].g_x\[7\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_16_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3495_ _1550_ _1553_ _1535_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2446_ _0074_ _0080_ _0111_ _0118_ g.g_y\[6\].g_x\[2\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2515_ _0180_ _0182_ _0173_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3564_ _1145_ _1150_ _3564_/ZN vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2377_ _0025_ _0049_ _0052_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4047_ g.g_y\[0\].g_x\[3\].t.out_sc _4047_/E g.g_y\[0\].g_x\[3\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_66_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2186__S _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2300_ g.g_y\[5\].g_x\[6\].t.r_v _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2231_ g.bi_l\[50\]\[0\] g.g_y\[6\].g_x\[2\].t.r_h _1716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_0_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3280_ g.g_y\[1\].g_x\[1\].t.r_h _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2162_ _1539_ _1541_ _1649_ _1650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2093_ g.g_y\[0\].g_x\[2\].t.r_d _1581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2995_ _0632_ _0633_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1877_ _1336_ _1370_ _1371_ _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3616_ _0232_ _0252_ _0259_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3547_ _1697_ _1700_ _1127_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1946_ _1439_ _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3478_ g.g_y\[0\].g_x\[5\].t.r_h _1077_ _1078_ _1316_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2429_ _0082_ _0101_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_67_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3403__B _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3165__A1 g.bi_l\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2140__A2 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2515__I1 _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3640__A2 _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2780_ _1451_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3401_ _0998_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_13_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3459__A2 _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2214_ g.g_y\[0\].g_x\[1\].t.r_d _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3194_ _0661_ _0655_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3263_ _0774_ _0882_ _0884_ g.g_y\[2\].g_x\[3\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3332_ net35 _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2145_ g.g_y\[7\].g_x\[3\].t.r_h _1633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2076_ _1564_ _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1929_ _1421_ _1422_ _1423_ _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2978_ _0616_ _0618_ _0619_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_16_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_70_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2263__I _1745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3950_ g.g_y\[2\].g_x\[6\].t.w_si net124 g.g_y\[2\].g_x\[6\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ net69 _3881_/E g.g_y\[4\].g_x\[4\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2832_ _1440_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2763_ _0401_ _0402_ _0403_ _0409_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_9_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2901_ _0544_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2694_ _0334_ _0336_ _0337_ _0341_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3177_ net42 g.bi_l\[15\]\[1\] g.g_y\[1\].g_x\[7\].t.r_d _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3315_ net45 _0883_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3246_ _0709_ _0703_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2128_ g.bi_l\[52\]\[0\] g.g_y\[6\].g_x\[4\].t.r_h _1616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2059_ _1548_ _1528_ _1549_ _1545_ _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_24_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2591__A2 _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2334__A2 _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3031_ _0621_ _0623_ _0668_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3100_ g.g_y\[3\].g_x\[1\].t.r_d _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3933_ net55 _3933_/E g.g_y\[3\].g_x\[2\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3795_ g.g_y\[6\].g_x\[5\].t.out_sc _3795_/E g.g_y\[6\].g_x\[5\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_61_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2948__I1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3864_ g.g_y\[5\].g_x\[0\].t.out_sc _3864_/E g.g_y\[5\].g_x\[0\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_2746_ g.g_y\[3\].g_x\[6\].t.r_v _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2815_ _0440_ _0450_ _0464_ _0442_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_1_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2677_ _0334_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3229_ g.g_y\[1\].g_x\[4\].t.r_h _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__2261__A1 _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2600_ _0215_ _1796_ _1799_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3580_ _1636_ _1656_ _1663_ _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_43_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout122_I net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2555__A2 _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2393_ _1557_ _0065_ _0066_ _0067_ g.g_y\[6\].g_x\[4\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2462_ _1399_ _1401_ g.g_y\[7\].g_x\[0\].t.r_v _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2531_ _0198_ _0178_ _0179_ _0173_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_2_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4063_ g.g_y\[0\].g_x\[0\].t.w_dh _4063_/E _4063_/RN g.bi_l\[0\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3014_ _0591_ _0593_ _0651_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_46_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3916_ g.g_y\[3\].g_x\[5\].t.w_si net123 g.g_y\[3\].g_x\[5\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3847_ net78 _3847_/E g.g_y\[5\].g_x\[3\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3778_ net96 _3778_/E g.g_y\[7\].g_x\[1\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_46_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2729_ _0203_ _0195_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout133 net134 net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout100 g.g_y\[7\].g_x\[3\].t.out_sc net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout111 net115 net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout122 net126 net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_40_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_0_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3980__CLK net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1962_ _1453_ g.g_y\[7\].g_x\[6\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ _1384_ _1386_ _1387_ _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3632_ _0422_ _0424_ _0425_ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3563_ net5 net4 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3701_ _1260_ _0981_ _0803_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2514_ _1340_ _1342_ _0181_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2445_ _0115_ _0117_ _0074_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2376_ _0043_ _0042_ _0050_ _0051_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3494_ g.g_y\[1\].g_x\[4\].t.r_v _0857_ _1091_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_3_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4046_ g.g_y\[0\].g_x\[3\].t.w_si net130 g.g_y\[0\].g_x\[3\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_27_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2455__A1 _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2230_ _1353_ _1354_ _1714_ _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2161_ g.bi_l\[59\]\[0\] g.g_y\[7\].g_x\[3\].t.r_h _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2092_ g.g_y\[0\].g_x\[2\].t.r_h _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_61_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1945_ _1438_ _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2994_ _0399_ _0398_ _0414_ _0417_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_16_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3615_ _1362_ _1187_ _1189_ _1190_ g.g_y\[5\].g_x\[7\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1876_ _1303_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3546_ _1132_ _1134_ _1136_ _1137_ _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_31_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2428_ net76 _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3477_ _1482_ _1485_ g.g_y\[0\].g_x\[5\].t.r_h _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2359_ _0032_ _0034_ _0024_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4029_ net33 _4029_/E g.g_y\[0\].g_x\[6\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_input15_I in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3165__A2 g.g_y\[0\].g_x\[6\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3380__I _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3400_ _0998_ _1003_ _1011_ g.g_y\[1\].g_x\[5\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3331_ _0945_ _0948_ _0937_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2144_ _1600_ _1630_ _1631_ _1632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2213_ _1686_ _1321_ _1687_ _1691_ _1698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3193_ g.g_y\[2\].g_x\[5\].t.r_h _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3262_ net47 _0883_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input7_I in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2075_ _1451_ _1564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1928_ g.bi_l\[61\]\[0\] g.g_y\[7\].g_x\[5\].t.r_h _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1859_ net85 g.bi_l\[48\]\[1\] g.g_y\[6\].g_x\[0\].t.r_d _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2977_ _0565_ _0568_ _0563_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3529_ _1581_ _1121_ _1123_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_12_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3147__A2 _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3310__A2 _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2454__I _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2900_ g.g_y\[3\].g_x\[0\].t.r_v _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2762_ _0399_ _0398_ _0414_ _0391_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2831_ _0472_ _0480_ g.g_y\[4\].g_x\[4\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3880_ g.g_y\[4\].g_x\[4\].t.w_si net115 g.g_y\[4\].g_x\[4\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3377__A2 _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2693_ _0333_ _0342_ _0348_ _0350_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3314_ _0931_ _0932_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2127_ _1612_ _1613_ _1614_ _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3176_ g.g_y\[1\].g_x\[7\].t.r_h _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3245_ _0820_ _0822_ _0868_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2058_ _1529_ _1532_ _1533_ _1548_ _1549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_24_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3531__A2 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3030_ _0621_ _0415_ _0418_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3863_ g.g_y\[5\].g_x\[0\].t.out_sc _3863_/E g.g_y\[5\].g_x\[0\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3932_ g.g_y\[3\].g_x\[2\].t.w_si net114 g.g_y\[3\].g_x\[2\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3794_ g.g_y\[6\].g_x\[6\].t.w_na _3794_/E _3794_/RN g.bi_l\[54\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2745_ _1772_ _1774_ _0397_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2814_ _0443_ _0446_ _0447_ _0440_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2676_ g.g_y\[3\].g_x\[1\].t.r_v _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3522__A2 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1836__A2 _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3159_ _0390_ _0415_ _0418_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3228_ _0798_ _0799_ _0851_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_64_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3139__B _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2269__I _1745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2530_ _0176_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_fanout115_I net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2392_ net89 _1743_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2461_ _1395_ _1383_ _1394_ _0130_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_23_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4062_ net27 _4062_/E g.g_y\[0\].g_x\[0\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3013_ g.bi_l\[22\]\[0\] g.g_y\[2\].g_x\[6\].t.r_h _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3846_ g.g_y\[5\].g_x\[3\].t.w_si net120 g.g_y\[5\].g_x\[3\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3915_ net59 _3915_/E g.g_y\[3\].g_x\[5\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_19_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3440__A1 _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3777_ net96 _3777_/E g.g_y\[7\].g_x\[1\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2659_ _0107_ _0101_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2728_ _0200_ _0204_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout134 net1 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout101 g.g_y\[7\].g_x\[3\].t.out_sc net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3782__CLK net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout112 net113 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout123 net126 net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1961_ net104 _1450_ _1452_ _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_56_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1892_ g.bi_l\[48\]\[0\] g.g_y\[6\].g_x\[0\].t.r_v _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3700_ _0982_ _0984_ _0985_ _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2513_ g.bi_l\[47\]\[0\] g.g_y\[5\].g_x\[7\].t.r_v _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3725__A2 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3631_ _1200_ _1203_ g.g_y\[5\].g_x\[1\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3562_ net8 net7 _1148_ _3562_/ZN vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3493_ g.g_y\[1\].g_x\[4\].t.r_v _0859_ _0862_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_3_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2444_ _0068_ _0061_ _0116_ _1612_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2375_ g.g_y\[5\].g_x\[4\].t.r_d _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4045_ g.g_y\[0\].g_x\[3\].t.out_sc _4045_/E g.g_y\[0\].g_x\[3\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_3829_ g.g_y\[5\].g_x\[7\].t.w_dh _3829_/E _3829_/RN g.bi_l\[47\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__3468__I g.g_y\[0\].g_x\[6\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2455__A2 _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2160_ _1641_ _1647_ g.g_y\[7\].g_x\[2\].t.r_v _1648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2091_ _1572_ _1577_ _1578_ _1579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1957__A1 _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3614_ g.g_y\[6\].g_x\[7\].t.r_v _1361_ _0171_ _1362_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1875_ _1338_ _1361_ _1369_ _1302_ _1370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_61_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1944_ _1297_ net2 _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2993_ _0409_ _0408_ _0416_ _0391_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3476_ _1484_ _1466_ _1476_ _1076_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_2427_ _0096_ _0098_ _0099_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3545_ _1320_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2289_ _1411_ _1768_ _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3820__CLK net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2358_ _1529_ _1532_ _0033_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4028_ g.g_y\[0\].g_x\[7\].t.out_sc _4028_/E g.g_y\[0\].g_x\[7\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3970__CLK net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3330_ _0946_ _0553_ _0947_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2667__A2 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2143_ _1540_ _1631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2212_ _1684_ _1683_ _1696_ _1673_ _1697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3192_ _0789_ _0818_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3261_ _1444_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_64_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2074_ _1561_ _1562_ _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_46_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ net104 g.bi_l\[61\]\[1\] g.g_y\[7\].g_x\[5\].t.r_d _1422_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1858_ _1352_ _1353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2976_ _0567_ _0550_ _0559_ _0617_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_3459_ _1311_ _1310_ _1330_ _1333_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_55_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3528_ _1106_ _1098_ _1122_ _1580_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_64_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3866__CLK net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3605__B _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2830_ _0473_ _0475_ _0479_ _0029_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2761_ _0393_ _0394_ _0395_ _0399_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2692_ _0333_ _0349_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3244_ _0820_ _0659_ _0662_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2888__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3313_ _0739_ _0738_ _0750_ _0754_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2057_ g.g_y\[7\].g_x\[4\].t.r_v _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_2126_ g.bi_l\[50\]\[0\] g.g_y\[6\].g_x\[2\].t.r_h _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3175_ _0798_ _0799_ _0801_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3688__I1 _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2959_ g.g_y\[2\].g_x\[7\].t.r_h _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_16_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ g.g_y\[5\].g_x\[0\].t.w_si net110 g.g_y\[5\].g_x\[0\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2813_ _0442_ _0451_ _0460_ _0462_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3931_ net55 _3931_/E g.g_y\[3\].g_x\[2\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XANTENNA__3047__A2 _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3793_ g.g_y\[6\].g_x\[6\].t.w_dh _3793_/E _3793_/RN g.bi_l\[54\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_41_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2744_ g.bi_l\[38\]\[0\] g.g_y\[4\].g_x\[6\].t.r_v _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2675_ g.g_y\[4\].g_x\[1\].t.r_d _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3227_ g.bi_l\[13\]\[0\] g.g_y\[1\].g_x\[5\].t.r_h _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2109_ g.g_y\[0\].g_x\[3\].t.r_d _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_37_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3158_ g.g_y\[2\].g_x\[6\].t.r_d _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3089_ _0714_ _0723_ g.g_y\[3\].g_x\[3\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3210__A2 _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2572__I1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2460_ net94 _1376_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_2_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2391_ _0057_ _0059_ _0063_ _0055_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4061_ net27 _4061_/E g.g_y\[0\].g_x\[0\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_34_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3012_ _0647_ _0648_ _0649_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3776_ g.g_y\[7\].g_x\[1\].t.w_si net118 g.g_y\[7\].g_x\[1\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3845_ net77 _3845_/E g.g_y\[5\].g_x\[3\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3914_ g.g_y\[3\].g_x\[6\].t.out_sc _3914_/E g.g_y\[3\].g_x\[6\].t.r_v vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA__3440__A2 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout102 g.g_y\[7\].g_x\[4\].t.out_sc net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2658_ g.g_y\[5\].g_x\[2\].t.r_h _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2727_ _0277_ _0379_ _0381_ g.g_y\[4\].g_x\[7\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout113 net115 net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2589_ _0234_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_69_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout124 net125 net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3259__A2 _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1891_ g.bi_l\[48\]\[1\] net85 _1385_ _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3630_ _1201_ _1202_ _1707_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1960_ _1451_ _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2443_ _1625_ _1628_ _0068_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3492_ g.g_y\[0\].g_x\[4\].t.r_v _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3561_ _1148_ _1149_ _3561_/ZN vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2512_ _0176_ _0178_ _0179_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2374_ _0036_ _0038_ _0039_ _0043_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4044_ g.g_y\[0\].g_x\[4\].t.w_na _4044_/E _4044_/RN g.bi_l\[4\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3828_ net84 _3828_/E g.g_y\[5\].g_x\[7\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_3759_ g.g_y\[7\].g_x\[5\].t.w_dh _3759_/E _3759_/RN g.bi_l\[61\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output21_I net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3404__A2 _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ g.g_y\[0\].g_x\[3\].t.r_v _1578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2992_ _0631_ net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1874_ _1338_ _1364_ _1368_ _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1943_ _1372_ _1437_ g.g_y\[7\].g_x\[7\].t.w_dh vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3613_ _0214_ _1188_ _0209_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3475_ _1477_ _1484_ _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2426_ g.g_y\[5\].g_x\[2\].t.r_h _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_43_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3544_ _0129_ _0131_ _1135_ _1132_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2288_ _1764_ _1766_ _1767_ _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2357_ g.bi_l\[52\]\[0\] g.g_y\[6\].g_x\[4\].t.r_v _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4027_ g.g_y\[0\].g_x\[7\].t.out_sc _4027_/E g.g_y\[0\].g_x\[7\].t.r_d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_50_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2373__A2 _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3260_ _0879_ _0881_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1875__A1 _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3616__A2 _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2073_ _1548_ _1528_ _1549_ _1524_ _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2142_ _1602_ _1622_ _1629_ _1593_ _1630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2211_ _1674_ _1675_ _1677_ _1684_ _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3191_ _0790_ _0811_ _0817_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2975_ _0567_ _0560_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1926_ g.g_y\[7\].g_x\[5\].t.r_h _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_1857_ g.g_y\[6\].g_x\[0\].t.r_h _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3527_ _1595_ _1598_ _1106_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2107__A2 _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3458_ _1060_ _1324_ _1332_ _1300_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2409_ g.g_y\[5\].g_x\[2\].t.r_d _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3389_ _0659_ _0662_ _0639_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2337__A2 _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3810__CLK net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2760_ _0391_ _0400_ _0410_ _0412_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2691_ g.g_y\[4\].g_x\[1\].t.out_sc _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3243_ g.g_y\[2\].g_x\[4\].t.r_h _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3312_ _0930_ _0744_ _0753_ _0734_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2125_ net87 g.bi_l\[50\]\[1\] g.g_y\[6\].g_x\[2\].t.r_d _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2056_ _1524_ _1536_ _1544_ _1546_ _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_3174_ g.bi_l\[13\]\[0\] _0800_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_16_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1909_ g.g_y\[7\].g_x\[6\].t.r_h _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2025__A1 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2958_ _0597_ _0598_ _0599_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_8_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2889_ _0491_ _0528_ _0530_ _0432_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_67_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3930_ g.g_y\[3\].g_x\[3\].t.w_na _3930_/E _3930_/RN g.bi_l\[27\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_3792_ net93 _3792_/E g.g_y\[6\].g_x\[6\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_46_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3861_ g.g_y\[5\].g_x\[0\].t.out_sc _3861_/E g.g_y\[5\].g_x\[0\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
X_2743_ _0393_ _0394_ _0395_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2812_ _0442_ _0461_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2674_ g.g_y\[5\].g_x\[1\].t.r_d _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3157_ _0784_ net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3226_ _0846_ _0847_ _0849_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2039_ _1529_ _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2246__A1 _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2108_ _1580_ _1582_ _1584_ _1588_ _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_37_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3688__S _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3088_ _0715_ _0717_ _0722_ _0453_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_60_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2390_ _0023_ _0054_ _1531_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4060_ g.g_y\[0\].g_x\[0\].t.w_si net129 g.g_y\[0\].g_x\[0\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3011_ g.bi_l\[20\]\[0\] g.g_y\[2\].g_x\[4\].t.r_h _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_64_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2779__A2 _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3913_ net61 _3913_/E g.g_y\[3\].g_x\[6\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_19_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3775_ net97 _3775_/E g.g_y\[7\].g_x\[1\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3844_ net79 _3844_/E g.g_y\[5\].g_x\[4\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_42_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2726_ net71 _0380_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout103 g.g_y\[7\].g_x\[4\].t.out_sc net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2657_ _0266_ _0268_ _0317_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2588_ _0233_ _0241_ _0249_ _0251_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
Xfanout125 net126 net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout114 net115 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3209_ _0831_ _0833_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1817__I1 _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout120_I net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1890_ g.g_y\[6\].g_x\[0\].t.r_d _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3560_ _1147_ net7 _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2442_ g.g_y\[6\].g_x\[1\].t.r_h _0113_ _0114_ g.g_y\[6\].g_x\[2\].t.r_h _0115_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2373_ _0024_ _0034_ _0048_ _0026_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3491_ _1441_ _1088_ _1089_ g.g_y\[0\].g_x\[5\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2511_ g.bi_l\[31\]\[0\] g.g_y\[3\].g_x\[7\].t.r_v _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4043_ g.g_y\[0\].g_x\[4\].t.w_dh _4043_/E _4043_/RN g.bi_l\[4\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3827_ net84 _3827_/E g.g_y\[5\].g_x\[7\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3758_ net105 _3758_/E g.g_y\[7\].g_x\[5\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2709_ _0153_ _0155_ _0158_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_30_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2924__A2 _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3689_ _0695_ _1247_ _1249_ _1250_ g.g_y\[2\].g_x\[2\].t.w_na vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_15_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3168__A2 _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3340__A2 _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1942_ _1373_ _1403_ _1436_ _1303_ _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_61_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2991_ g.bi_l\[31\]\[0\] _0406_ _0615_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_16_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1873_ _1357_ _1356_ _1366_ _1367_ _1368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3612_ _0215_ _0217_ _0218_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2703__B _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3543_ g.g_y\[7\].g_x\[0\].t.r_v _1399_ _1401_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_43_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3474_ _1069_ _1071_ _1073_ _1074_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2425_ _0036_ _0038_ _0097_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2356_ _0028_ _0030_ _0031_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2287_ _1764_ _1431_ _1434_ _1767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4026_ g.g_y\[0\].g_x\[7\].t.w_si net130 g.g_y\[0\].g_x\[7\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2070__A2 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2684__I1 _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2833__A1 _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _1673_ _1685_ _1692_ _1694_ _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3190_ _0813_ _0816_ g.g_y\[1\].g_x\[6\].t.r_v _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3313__A2 _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1875__A2 _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2072_ _1551_ _1538_ _1552_ _1545_ _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2141_ _1602_ _1625_ _1628_ _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1925_ _1417_ _1418_ _1419_ _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2974_ _0563_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1856_ _1348_ _1349_ _1350_ _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3526_ g.g_y\[0\].g_x\[1\].t.r_h _1119_ _1120_ _1583_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__3552__A2 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2339_ _1489_ _1497_ _1511_ _1514_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3457_ _1325_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2408_ g.g_y\[5\].g_x\[2\].t.r_v _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3388_ _1454_ _1479_ _0999_ _0641_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4009_ g.g_y\[1\].g_x\[3\].t.w_dh _4009_/E _4009_/RN g.bi_l\[11\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_15_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2690_ _0344_ _0346_ _0347_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3311_ _0745_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_7_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2124_ _1611_ _1612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3173_ g.g_y\[1\].g_x\[5\].t.r_h _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3242_ _0837_ _0864_ _0865_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input5_I in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2055_ _1545_ net102 _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1839_ _1325_ _1324_ _1332_ _1333_ _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1908_ _1375_ _1397_ _1402_ _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_32_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2957_ g.bi_l\[16\]\[0\] g.g_y\[2\].g_x\[0\].t.r_h _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2888_ _0086_ _0493_ _0533_ g.g_y\[4\].g_x\[2\].t.r_d _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3509_ _1590_ _0122_ _1104_ _1105_ g.g_y\[0\].g_x\[4\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1839__A2 _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3452__A1 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3791_ net93 _3791_/E g.g_y\[6\].g_x\[6\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
XFILLER_0_58_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ g.g_y\[5\].g_x\[1\].t.w_na _3860_/E _3860_/RN g.bi_l\[41\]\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2742_ g.bi_l\[22\]\[0\] g.g_y\[2\].g_x\[6\].t.r_v _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_26_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2811_ net58 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2673_ _0277_ _0330_ _0331_ g.g_y\[5\].g_x\[2\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2107_ _1578_ _1577_ _1594_ _1568_ _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_37_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3156_ _0781_ _0783_ g.g_y\[2\].g_x\[7\].t.r_h _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3691__A1 g.g_y\[3\].g_x\[0\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3087_ _0718_ _0720_ _0721_ _0715_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3225_ g.bi_l\[11\]\[0\] _0848_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_64_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2038_ g.g_y\[6\].g_x\[4\].t.r_v _1529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__2246__A2 _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3989_ g.g_y\[1\].g_x\[7\].t.w_dh _3989_/E _3989_/RN g.bi_l\[15\]\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_0_13_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2182__A1 _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3434__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1996__A1 _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3737__A2 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3950__CLK net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3010_ net49 g.bi_l\[20\]\[1\] g.g_y\[2\].g_x\[4\].t.r_d _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3843_ net79 _3843_/E g.g_y\[5\].g_x\[4\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_34_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3912_ g.g_y\[3\].g_x\[6\].t.w_si net112 g.g_y\[3\].g_x\[6\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3774_ net98 _3774_/E g.g_y\[7\].g_x\[2\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_4
X_2656_ _0266_ _0049_ _0052_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2725_ _1756_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout104 g.g_y\[7\].g_x\[5\].t.out_sc net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2587_ _0233_ _0250_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout115 net121 net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout126 net133 net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3208_ _0832_ _0645_ _0658_ _0661_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3139_ _0732_ _0758_ _0760_ _0432_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_64_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3490_ net31 _1039_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2510_ g.bi_l\[31\]\[1\] net62 _0177_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout113_I net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3846__CLK net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2441_ _1725_ _1729_ g.g_y\[6\].g_x\[1\].t.r_h _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2372_ _0027_ _0030_ _0031_ _0024_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4042_ net31 _4042_/E g.g_y\[0\].g_x\[4\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XPHY_EDGE_ROW_20_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3996__CLK net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3826_ g.g_y\[5\].g_x\[7\].t.w_si net116 g.g_y\[5\].g_x\[7\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3757_ net105 _3757_/E g.g_y\[7\].g_x\[5\].t.r_d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA__2171__B _1658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2708_ _0319_ _0321_ _0365_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2639_ _0242_ _0243_ _0299_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3688_ _0917_ _0887_ _0498_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2160__I1 _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2612__A2 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1872_ g.g_y\[6\].g_x\[7\].t.r_d _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1941_ _1404_ _1428_ _1435_ g.g_y\[7\].g_x\[7\].t.r_h _1436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_61_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2990_ _0481_ _0627_ _0628_ _0630_ g.g_y\[3\].g_x\[7\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_9_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3611_ _0174_ _0197_ _0205_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3473_ _1314_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3542_ g.g_y\[1\].g_x\[0\].t.r_v _0952_ _1133_ _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2286_ _1426_ _1416_ _1425_ _1765_ _1766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_2424_ g.bi_l\[43\]\[0\] g.g_y\[5\].g_x\[3\].t.r_h _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2355_ g.bi_l\[36\]\[0\] g.g_y\[4\].g_x\[4\].t.r_v _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_67_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4025_ g.g_y\[0\].g_x\[7\].t.out_sc _4025_/E g.g_y\[0\].g_x\[7\].t.r_h vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XANTENNA__2842__A2 _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3809_ net87 _3809_/E g.g_y\[6\].g_x\[2\].t.r_h vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_2
XTAP_TAPCELL_ROW_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2833__A2 _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _1618_ _1617_ _1626_ _1627_ _1628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2071_ _1557_ _1558_ _1559_ _1560_ g.g_y\[7\].g_x\[5\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1855_ g.bi_l\[54\]\[0\] g.g_y\[6\].g_x\[6\].t.r_h _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1924_ g.bi_l\[63\]\[0\] g.g_y\[7\].g_x\[7\].t.r_h _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2973_ g.g_y\[3\].g_x\[7\].t.r_h _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3525_ _1697_ _1700_ g.g_y\[0\].g_x\[1\].t.r_h _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3456_ _1327_ _1746_ _1059_ g.g_y\[1\].g_x\[0\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2269_ _1745_ _1751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2338_ _1505_ _1504_ _1513_ _1490_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2407_ _1643_ _0079_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3387_ _1482_ _1485_ g.g_y\[0\].g_x\[5\].t.r_v _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4008_ net38 _4008_/E g.g_y\[1\].g_x\[3\].t.r_v vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_33_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2815__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Left_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_60_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2990__A1 _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3310_ _0747_ _0532_ _0927_ _0929_ g.g_y\[2\].g_x\[2\].t.w_si vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2123_ g.g_y\[6\].g_x\[2\].t.r_h _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3172_ net40 g.bi_l\[13\]\[1\] g.g_y\[1\].g_x\[5\].t.r_d _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3241_ _0445_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2054_ g.g_y\[7\].g_x\[4\].t.r_d _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1838_ g.g_y\[0\].g_x\[7\].t.r_d _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1907_ _1399_ _1401_ _1374_ _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2956_ net44 g.bi_l\[16\]\[1\] g.g_y\[2\].g_x\[0\].t.r_d _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2887_ _0495_ _0516_ _0522_ _0086_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3508_ _1095_ _1100_ _1102_ _1452_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3439_ _1044_ _1697_ _1700_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__3461__A2 _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3790_ g.g_y\[6\].g_x\[6\].t.w_si net127 g.g_y\[6\].g_x\[6\].t.out_sc vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2672_ net75 _0072_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2741_ g.bi_l\[22\]\[1\] net51 g.g_y\[2\].g_x\[6\].t.r_d _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2810_ _0456_ _0458_ _0459_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3224_ g.g_y\[1\].g_x\[3\].t.r_h _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
.ends

